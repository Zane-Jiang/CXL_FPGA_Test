// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
sNTofcDXWFbY41shhy/pwf0pMiv6u8kwNvaxPmq2FLoUB3rCd2fExVVKRnCndoRD
gDoqkcWoHs2TNtCfKyK622sg0vciptr45/9gW0cHrxys9pVrAVZKXW/N7BtSvRV/
lWYDuW1iUZ6g172YOSz+W1hwgeiOU2NvWuGerTL6cvEjUClRQjs8Ig==
//pragma protect end_key_block
//pragma protect digest_block
yMNQqEyjgQlytfHHtnOZlVGqV0o=
//pragma protect end_digest_block
//pragma protect data_block
JmiuLn5I2ir2HxEXm/3EffPc1wo6tTkvq07vz3jAQbi4rd29cFRIEMAxXEr98QgJ
V1cCPdOc5hOaRbwgz9bw+a76JxV4JKN3Wzc8biWUCfvZGredLzH0GE3PifbrpRYm
XgJb5s3uaOvRP8JtJhvxHcbTXXLKbbSdw2E7RS6k0nwkXrh85J9VnDyu19wkXZ2a
ERp50hT38PLy5DTzqN9H+DUZdf18w0jRBLt4md9Xk5Gh+cF15wmZZqhVzOVVlj/G
OfZf80NTnrhYEpGtCpnNcjotXQsTrtZZozkQa9BtxKcxIknLutjCeHaYg0KTOAv7
q9W60zkbXcm+qVVT2PNJV+o+QnoPkidXxhJQseetVeevysSCi/XeDM07gu6kRseU
dC/bm5gGNjzapbX5buYKwXT+jJ/GI+5V7U0vp4S8LHsvgoQ+K9r4DN/T+iELl/BR
QG4aHddxTez/WbsvP1VeZblLPYvOUXG0ZZp8FyG3KkJZTL3e/9+6W0ZpNeEP7BMV
sMTAJfRVNxu29u8KZULHcJ4zTkYs1Ti63x+vViEd61cTCGATf7sdDVoVP4Y0ANxZ
10Vs392QFNJye8i41s0k3Iielbg79GRy8vrtu8HWsHJzhK1Kj81rYq43QcxsEkqX
iaENNg/XUbCM1EvbMOPuIu4k7wZ5j7GII7KqU1tP26DPHl2VeFTOFGxhTOTAEKgF
rrN9lhgKH5QGjsB1ceDXDfC1UbpXUgJpPMA72IxdJLoculJ8jznxuXabDHYJqw3h
/mvE5JCOblY7BUYhzpzI+Xh8oqULVPiAJYLPZpgZ/67n1cQSSxPK8epTn9oMxH1N
daFz89UqmwNZSmgpvFAmEdUoMiBOwO1Qo6eA5Elc13aFHLkGsviDyEJBdKDUP2Bu
i+u5aXIjNgNumQKZyNgq9Y/xQD0bSk7H0r5Vs5r4oKAgJyI7/hhobbNOUMnb0yA0
HZLaXd3uznBQwXiwSzzZrRJprlvahoCwmd5VVT7UmqixpP8Cy+FqALPL9d+L8BPl
/5tPE0jrmTaa4Yc14eWUqxAJMlI6AnUF59pdnoaQoF2MYlwk78W1fu7oG+GfPez0
HNuzc3MiPe0TvicW9YVaQe5FZQmecB66AxevKHwRBX9N6IjBt+4TNEn+Ki6oxsm7
BH3a7/1JSiEWTo/Q20xp3Dxs+ENzhDYJfFM9m/0yb5wzUsukRDtv3Ps0VGlyTrGm
/0zw6wXVQ5qaDLcAst8O/6Mm5tT8tw2QSvZGY7voR+K+FlB0oi2eu9oMtypbK/TX
ggwpdFvRvQkBfhQG6YedTt6d6dA2fL5OUcRsL7+/S13fBXzxppxJ/635OsS0sRSz
30kNnPq6c0SOmtAGf/ZoAgn6fn1yFp2pKi8SWskoJ7dEXii2v5LanJ6bVtzXkyiB
wjhTtKwBVYSF17FcrWN4S4H8R26Sv3ajx9ZFhUiOncTZdN49H9+Ix8hSMb9jL8lu
5dfkhaBqGFMM587Xj/eA84CsIueEdr/3CnVmxEB4cFN3orj/XI3chGyqeGUu/Bf2
ayz27jTbGuUfxWpDgrf0+elnDPtyQITWX0HA+2i1Uds6dSQcI6RM8fnK6gKJalW1
k9m4X9OJsA7KrVNNb6gDbLa/fxzOZez17i6QpG9JnOer2VeC4yvJadjCb8CLg3Le
Z4jZPEdJcQ8vXBwqY0Ppy7dwN6xXGqwXs+caZ3E1yXbwj/YvaLWZUucklEqdyyVd
jGFao04Q2D0PyHnZKo95hnx6AvhTNhcmLQbYj1yIfXj7ahqh+yO9q47PJCnfPkaV
wVyefqNBkCu6sfviCj6eww0NTV36klj2YZNAb2hRtHSoaok+Ivy76FgiMzHsX2YR
nZb+k/QM6amUknPVnIuPWqTyPkfn2SMQ81L7Bdot6dsPD2oQzKFgLu6hnRtcSflh
BKPgL+JYUnlmqhVOzpUwyh/q2JIJRtGE255jYYZsFMWX/uwcDQSYxC/jd7HDo0AQ
WZ85/t2EMpt9YXFxDHyp30Pgp5GB/c0f2oa7KHav2dkZwqR2JMxd620ce5P/ZHoQ
q49+QLfFYTHEM1kI06IzlN/jl/Km5mnR7XBdegTnBGO1xHBKqnLzDjtualFf+3g6
DpG2SwBkF0DEOghxLyn+hlXS+xQWlaXT1Ef8O7QrUKWG9k/IMvQoqhwNOsenpBZG
poVprL8eABvl7ca3nOT8AYHj1LpTWe8iNUvD/aQd/4HA+tgLLmegQ5qysx6Y01+m
hUvNB4o58LHf1HH4X8FAbhayXfU6DZRKv8ZLcy4oSlyTXutqq75/Ybt0Csdyv3u7
UjtyTDIPI9hgi8/gXhQbn8U7aab6j+CqcPtDERzbySQtGIhLCbcF7r2CRxZPN8Xz
ebUyKncfAmolxsrUFBCvrydg8kQRV+741QtCWIL9wJhEzZ5Q0cSFeO+HsJ8PvYmt
5iTgCV240vVI33UX3bGf4t9dFCKXp5nWZE0kSdQrnI/rO2pankNUbQt8ZZcf6I1D
kguaI+SDIZSBA9+6uXyWsZNKcPVV8Bd02Tn+u9Do5Qcl2aPJrI3zzF7rDPy5gkaL
4L5QrBf+ditSp/4lpmTvoHqIC+OtFiSWhq0/aRY4OoDUCb0tAvctYk6O2f9aza2c
Ezs9S/D4wbecafZwnzMis9dKX8nfyuTxaArA2iQBdsz/KrNIkG9u23hJg1XZYpUi
39n7C7wkNT1vPIYVg9S4yQlAiSYdFYBZRjVJUljMDu/H0EL8lMFm+lDvBv89LWUb
5LUnsvPdQ9ZD2PjRgEuIs6fRP27jBUd14fYj+7HykgxYNLTJt5qjx1zH3rxRQkEi
1W0eq8gP5NPLSnUYVfshIMi7UhsH7i9+8bqm09n33rV+5c+mFwx9qoiZJVTIZ1y7
FIEG1NXiLwAm0nj6cqS16hjsiCkHvuox1ZgIulip44nrjA1ivaF3TdrLeMdTb7kR
v3rOhIH0eFE7zn0WrzpA8YRU0ZqQLBY1TeRFVmWFxHSLUXnuJlycXqgc4PfR6V+O
u9UCDb0PGOpmm5LvggVFBzxnJ1vXvzG2g5k7StXUK/kEboQqIscDsxGJPx2XxU3s
Qqkc7TPUBBa1jLSUxn6TnrzprENNjNorDKJqM1Sib3w7CrGYWnjbrINbojORN8Rz
+deaJY6CwsEJffdMf7cU8qWGkwBoPPqbe/7nXjH+iU6GKNYV5AgEm3/YMHKFHndl
2dG5nzgM8UQ3vbtDORdLk/OkNZZZFjfTgRYw9zhUsjEMa0Wec5ta6PkeTmqLOcw7
GDODiMghwSBcWy1uAbbrA1e5bdAd19pdYrwUDOFb2EGBKrk27JT77hRwxqCWhd5+
mwylwkivy1EK/kX6Hlkq1HfOiS1fuaSezM4X5c7XZtqbzDK36LAiOg5R1p9CK1Ox
UYlb09mDlp4Fe2XznRC+lL1kankEFrqZxUsEBB3o5Y1nnVMuUtMkoLjfJVB1lbqf
wlW5gHbhyWdDsV1Dl6HyYKnRfA3pqmZ9z7Z8TQC8mZRfCc1jkMge3XhNYRHhMiyF
HLg6P4aW7DsSk/q7nn4o0vOv6jmb/b179kSKmCLlNY/84BKTR825amYdRs942NDe
90wqpA28txOsgOPsXkFu4P0XRYajVjqmH1cQUxgktdS46eAMqL3e+EB55WPTrMDL
jWrnAHm/ivI60y+nO2Ym0c8mEsWoNzTuefCRMYFEOFaqNz+yJXWKTBLXQLlWa33w
PK0e9ZFoVW5m6q+YE1xwLDRkIvSGM5EPbl9oj7XX/VyvZYdNXXtKhOVTG9+YmuOg
CziD1wkJRfS/PL8bwQhjDEMQqkS5AqlazgEWGFkc+HPJhmM3YVQ2iV9WlAfo6D7S
C9bcITqKGTiJmS4dywmA/uAElNeen7dp50h0J2nbZzpyiGsBqOB7rJEXiIetyiIz
uMbp54TcfHGTCN6IIcYyJiqwY+TwG5fc8X4El8duuLEOJkIfsKg0GJGrt3Cjtg28
Y5fX4xs1SVcbiGQp5spgey5eM/cVbKhnrUv4oTPIP4Uo9w7wKFalijEmtVmqReYj
DlmN17HmepaiMXPXZAeiNjmghaS5KzSUJyguXPRnUz6Fi4bQQGboR7FdnFJz25yY
7wul/+qpIkAodRwo7CVFN+7Bid/YpjaQ1J8Mce0nBIzqXRVxbmX7XnoicMprpxG8
uXnz9zIPmwaH6G3uWdZv/fNtQmWGi1Jdl3jVDq5DDdI/z5L7rAUL+NkiPoXRsLOg
VmA3rwcjANQuYGdqpz4v1Wj2l0TwApcx2+bNxKOm12AiGKAuBLfHy3sDt3R4Yg3X
70lnBM2oenuNxQbGCwldv+WBHADpcJOVVGEhnvrF8TVf70AdtAFwWWcdzCYnNQTV
f9tz3mJVEHuNoMZObUSBcpxs16w/RtjnTSrWcCoSXf2G8J1cnh2QlixE+RlTT74F
szTK291ktap1zCyPNNgK4zY1MqMmBAucF+7KpzA2S8eJdQyfQsO82Ft8OSvEeYJi
s6c3HY4JXkbbqmgVhFk0vRbTemuRTrxWPZnwsGvOlM+6MMQIGmtwMfRvuk4rTAfy
MPSnhZpVtGJfkIQoY614GUa1HIV3M0goXmRnAZDQXHSGHi2eFP9pDbfOytPkh9SA
sb2TRi67zNuerucrWIW0BbFm6YMx7cpLFRMj64q1KstzGr0tUUvCzzvo86OH1dou
fNKbC1g2bwiIVMZCn2ABiSOpb3M9LpVO4qtRNSZKu1VX1tBFgT0yVITBayE+XR2q
gJ8KMYdmiF/8y1RRWWMk6b+bDVenlPgWlTNaD7WnZwUMFxzGhc2nIhPyENr/XeKM
6Xq2+NtwBgOpGWgSsJ9Z1cSRTZ+6P3HvOnvGAGRBZ90Yoo4Se76dOFOMrRhUa3aV
GpuywUOP12I4uuCn4ClY4qiReZz8c4YcmD54RF6lfUdtfQl0EdDtdT1XoufWFNIa
3BQSpBvJrEBFRsrkkMH6Xmq/XbkW0HhYol9FhgozuTqBOg+QORh2zavmJFuvcZk1
ksVEDzp2kek2Ft7CgOYW/PZtUgioMcaHP0IqPc6VfyTdHUH9/fCeVIC6RRKFHFBC
0t0N3B9vmgkNX/1LoAp8oiZA8Oo4koCZB2gz6zNaPVwOq4c7nKYeLLJqGASctEBD
OOqw9sxndokw8rrYAar/CrzvwQbiaN7d5uZc6f6wedwp0h/VElAAY8NV68rBA15r
nmBWDcemSCsBWGZ3q1uopYtb7kT0D7EmjCBlDSjGOng03xazZpCEKd5vTS5rDQdv
9A0pz9WyXQhgPT5geo1CaQUBM39Tj+H6f04pozLyyH1hcYFhOImsLsk1dsI48Xgp
Tq8c+v15IQgCpjoJQtNO4Ob1NIPlop2np0fTiz3xagbP0tHfQbMbNskidRLPI3mM
i96H3GOnTiIt6t3hhu+nZ4mnDzahj2eJtLJWP7p3oJ9ZrBPbRC5KdROfv44QwI0g
bc5J46ZBrJ3CFtP3n8vrzSG4mqBgCFYTyIcXyQfTkdtQ7FlTjsfSOHMLZuXuM2m2
VJ/qislH2x9oJFqWWXaHfreFGN9yXnb7d7IxqIDXT54fNaS3HAK7jcmjgd1N28j5
NDW1fDi4GDQRCEIKreyYT4wbhYolATINbOIeY/V3xcclBB+jQClSg+kvJ6ZAORre
0FpMbiEYNvyU0T321cjwGAu01Ui/eWPq3UFB5tdxi1Agl44zWPPkl9pK9U6jEEkO
q3nQZUHJTKab8DDjhcBv+t7oq3d004k8D+BMAej52unDMkZwXkHwL5f30UQx+9Ul
0j0P/FmEhh50ykzEEdYDGQlPrpKwsWdfdQdL/pxiHgbZbkMcpIB04NIxYifQUIoe
gvEFYvMSHu0dDRBOaTLJuNG5wZgW+Y6qse1dgyeBiNaRmxhOErvNpADP6QaQi1tZ
UWraDteRS3cLFcZTEAsCbwn9qA0NfFmNGQDeugg85XRkU/nN8xng5m69HuXahLgA
TmMJ8ycZSqbtQKY/swZMujZCsPuPN2KCKYtpVbQ8FvMeWbgM8oQwN7V0k/2fOIP2
92lA3fvRbd/gVGWswZGd4VH/gOUj7/tTQYz+1kMmsty3OQJ3p2/CRLcjnz29yKVN
cC7XrDi1XjpqzUVBTGjnCbhAxs1o5+KQsGjKxx11WVE72Fiz7ixzLCMvLQrMXl0p
Yu92F3Pk3h2WvxmE2+7L1ZXEOQoNu7CXS6NIzay66Qb64DEEBU7sg5oVOdGdyOhO
XLMIJxtKwzjQ9OpuiHO/4DI7umTocn5eREJUNxMc0TaWSOgTLCqQyWPeXmawPw//
GUQrMu52Gk+Iztm3J7ibTvPeR5CdxnKrBZOMzq5LrLzB43KWV/+jlaOwem5CJn5n
IpX0qoVk+vb8BYzljT7S0nNGS8n7Ya4G55BUdOP7WKvnT7ZtfPSD4uAbcLVN+Xow
P4DJ+Rrj0lWgF1sXwY/oQ+u5E8c6K94uF+BOby2nJYWSLs6IPyec0aD1UWaFzXv1
UvgqUBvT4KKTFWh/UlJEl/NYYHguFVhpoajg6cmW5BceOE955j9gdHpXI4yMd6Gi
cNOU6EdSOmFCgbXClxUqlmbEHGZezHG6UZQz/QD7p65F5g+Sqx1fZyItFPUvGNMS
wbpd58RoECvKmppoiNeY6rMymOPQdwBlNCeJ8mqO5o/U/9bUdqdqj7Y9ZGoT4X9T
voGrEfw6Zmy/maBBjfFsEXI/3lipvrNGNPSg7pr/XC+/EXgGo24uJD8aUeL6uinG
NpW+MolaGj1bmw9PaffenmDlD8AH1OMgsR8WXftJw1EnJ6uWeZq9CddGykSJu4Vl
1yGOg6hRVJ5x2BLCgqfjn+186WngrRSTvzDBgss0BNdpYe50c6+eIWOMAHkgoLTA
16eDFqRAJZMgjTSQXKdus8VINkNrJ6BIJ434kj/PJ20zMxJITwNpBU8ncRqPEmKL
xhTK+/6rTEoOwlR8H1IDpBs2Mjo05H24YVXJKUTbPktTZaAOLxzf7szMuPQm562i
OTB8ih0ogh2IBCew4tgUY09XKYWFyG3qXVfmZoiE9PJQ19nsrUl+fu1W5k4/uoXL
ba7B2nER4u9AfoA2fTi37mYYYbRrPFeDSaFnoiu+InUY8137vYhO9h8Q/ntGyTkC
YrF+zwyIs6k448jbXtmbwHSutwA3i55jzbMR1NVSzyNy64nVsLgktZDT53mxO7Fj
hF415JJDuEq4AH7euZ7YhJmec/4e8fltr8NPYMMDbipRZeoQwFEXBZoiVB9T7b6m
U9ZcL9kyt9jdHa/eRBXdJxmsJ5CCoMxxNuO/zsB9y/L+HqB+8Z7iOuxRRF2hvwkW
6WWlOd1e65IzcEb7mAB28tWdqD1qxCeGEGqt2ZN6HGtRSUdS6oOQxYTHyE60wdPN
cPXGCxq3wt1dbMFfpOH/PYi3hxQb7dr+qXkeu/WhGJgFfb8A+kPhAkAOt26q0Fo7
Uvyv8gqmwhX4egabNDhYdyuaeVSKJmRmmGZdfbO7iY9n+yfS6BG4cOaRs7nrvO3v
ZmB7o3fhJKb7pephNeRQ1L0sleMiEL29oQRU/iT2qQyAycCSCI0fhszJ55qESVes
630RuzCMgskPZHII7amd1JpAN/1eItLiwzcAm6x1Kq5w0GQB+CBzKEXl1rHNXygT
stTTaPzLjpxP12pEu9WQPLirNBZ89Gqjw0VC9+r9H/A/WJKGUFtZIwYIEfsDxbAa
c+bUPAmK9o0hKrxlXsJC3rRJjw2nzVhhz1hfh3I/Zd5jgqYC7bgghIdVeWjuuZtG
nXR8OXR7uwRFmjzIdTOLRLlEBC3O0VuFb8QcQRvlWv6TNQaraCh82f2ECot6L956
K6MUHa48nF4jscRkGdEX3UXoliMubWxAgplS1b7nw2jo830jYKST0epgThVOY70A
dReC1HpYgFUksRtiVPxRTIrAoTB0DC7HNGAldB4WzpqV7OxkIYOz1lo10HhCJjcg
8cJS20OHIGK55/Kvdo3oQp9wF7KtjiM6KEw00RG7tEJnbd5iWnwkYdWzenf4K2t5
cYX9gfE6swnMrPyzovp3jPyxZJASQr7N4qaSzj5/MGf20i1AXKuwcswbKioQGtul
dGsw2Fm/klrqa1YuY6bZqBV2K2zxfv0pD0RXcOLvpmchoM1eKP1flDiheG9bH+Cg
yJSKOhDbghpe6CDdPo+CkZbuV8GsgCkIny625NO3GdscVSOveOcwljtfXnaCFtqt
Nwhu3uG1+SV0XHTeF+vfnnLjoi2CaCciCblYQ+gMew5rizp72sjRZZCWJjId7nV0
2YYZqreRCDiqRBIio+EgdfV12S8q7qFVpTbfQ3FWtfz/1iynZTw9ePgITaUUmnFH
ImsZ6ggcrbalST7t5aiBszk9fyCQDL9S38bHGOKfr10ICfjHbKn7PP871fm0VUFq
tDTda0+QRH26h5PzDkaY17RcguKbiRU4DV1PYeB7OcKpwM5TZPA6mbcjMPlRoxQi
kKd8KZPZijCKfu2Rzuw5/5vWJWZ+hqkh2DE+HjJvDK9Y+BeEMGFhZ3fCwBIGGbf5
2TFRJSv8Ry6vjP78qnOscinLBQXMiWn5b0XCKkbO/Kqcvdbl2M84PZJJKdRUW0Zv
6SmSPLzx6WkBVq9fA8B4rXKHHKgnaZgf/qmjY289O4lzKRiW3q8FjTDEQJLC+8CH
/GDRrQeR/I6rDd0khtoyE6h5vcB0AQdJaNQV/qXCFfTcIWLk5Je3ujYnQ+V2QJyT
twSDRXTC3+/+rLxGea86lAUvBktJu5I5Qm/NyHewy8oApc+FwgSLgmS3lyQiOfS4
A1xJSrfjmWa0sx9AzjDlbENhvaW2gLRModayUUaMNyEHaBgojo+QHR5oVC5cbbpH
eraADxbqEVhBA6L2r8lC17Y0t+b4Og1ZKockSittin5J5eVmKapMddHCg4Bhv3Yn
1B8huk7tMbx4s0rQZasdjUoWG4lSqjCv0+V4apj8MFecaAheG8propyjXyRPYdRj
KAStaPVIXKgKEKktpjm1Fl9I1FxG2DRpLefp/AdpqX+FuyMxnifK70LCYA8m2OR6
cnModQRPpeinGg8vjoEb5TSN1fu+xh81Hqx4vLMPWcvZ5XrzBgNi97m/qtKL6KvF
NNxT8EXwFjHOO9xDIQLN+tjFyl0jIlMdyy/wIWDi1F/GsXFF+WDqYl4OhQHL48rD
sLr0vGjd5gsDSYu+Ff5OGsZWlbuIfu29tKR+bzXWQ9noUSrlaM9cYYm4DzhShOnn
/4/lX+KbxOjkwPoNVhI5pwrMpupVjaOSQAPe9zLRwC3LZdB+R3vqYveyNREhuxam
N+1DxKCMHWQF/y6vfYScp+YMQMGrY3EyAtAtQoChAxWhn5F3jrv6vhdRbrag/+Ub
VM75wgEdyu0iBZMRhmn/pcwGyc2I2cjK0ctdZhaHHiHGJLkyMCTiDBYvkTHhiaeT
CtWD4hOohsjnAdi9FSwXUH4aCkHpZivXpkWNf6ffqS/XSFDe8vpJUY/57TkdVsLE
ewvV2Ej++S8CqjLFbFwyK1Jiv5GVe6EuAY2TtYLhruf9DauS9W3ZDxmVHoWdZzxa
oXKECFSGAy/64VTcRK/P0UwNC8sYT36hu9uEK+SHRGVbDLJmHkAr7+EvOHD1qB6+
bpsSRKn+MmYOopzq5EVNPcx0aPvzEyWZ/mNxEKmqed0MDWmhahVJ8JFamUNou8vx
x7VxM1EHpgKnDjhb7tOmwicjraNa91UlbdNdtSksTMY2vzErPESfZTenbbFLZpqN
08aDE+Jy5A/ezj0RIqoiUClIPjCrvKXl06xuzkhLnKuzbwE5OxkBlOxxXBZTzhQZ
S/HBf0S9zIYgMrGvH9WCtza9BjibCYOtHK5moGy0KbRF7uexGu5w5YZHuL1MKKj1
rAbrxnQbVhQg4s+G1tEWajpW7LeoCx0BOA5yazp3jSVvGK+9qaulb2ckGYhHG/GG
okmV1bwuvie0vjIm1dkNxF3z90c4pZKU5Jm7eUy77fg04IY+hKIVjpfTr5nTQ8Dd
kykcWKnoYNjYbWNcWeieh1MIOb1GZHAz8lHd1cFYMEvgzlIwzrFt1JSbgRYkQ1gu
OF83eNL1WRQfafgt/U8jF8bEBVwg91F6+liT9Ho6rI1Ov6wozc3UbtJ35pCKzE+h
rH42QhzKDBFd1dXRZbTELb6EljS1PZMJbsCO5jenprx3RKbkEGgGn7+K1h8G4zev
+p/hzESYQ5+TYFcsG1UGxIPwEDMRUT7HgZTn9i8TVOjTFOQlfL3E8Z/fPzhMVmUY
LZa9lxJa2tLvrK8vfxpRZ+gvGhkX3oKN6XfBCYby7Qsf7sE3FfMkjIv3X/RP2D6W
Dr55OjdWCOIszyhsI3UzWI6fsfdB1eGvNp5lX18+lNLZitFfAF69CIuJgGOCQ85u
QIQXiyT0Y4BjZ50Sg3Eq7wgbvZg97rvxFUoV76JfZXBAdkoJdFqPAbkCv6ZDVK4d
IIzuBdKzf6pAmCD5cF8dtk0aMoRhiVW3DwCfgDJX770M9KzhoKzU6x7d/KssQMpO
XyH+3jOS94sEg7UMM2mu2GaanarI3+piUVKYF06B2QKQSIVFi23QLfl0jhXJloBS
WBoAF36h6h4QPCIrkqiGC44aJf8KVaAXRpTy2ubRmgKOUyNVStQe8KRsFCYnZ0pJ
/uww5VMGfRK/Mha2sAgxrK3yjcyYx9g6vmLa66Ijq6JDPxBwTrT0UvQpjWBrx44F
j6M6U4wj6w0CH8tQb98Mgb9uR17gaI7Hh5uaqZF2xlTaNZtXRRfV3kPNXdMB/y41
qIpCFFm883Iix431eTKjXMnAXOfkn8/KIhnQUI6lfnfW62e0exR/OfuseGu8daoQ
Re8ypEzP7zOCe95ZkEsGiXmXeolQSCClGnkNi9T9BWwN2dMC6/lkJBhGlbUtZkrS
ClaVgzkRwkF7JN9K0vHySiamWH6faHQ/W5aQrKnN8TMhVzQ+tcOu5+y6W3V4Jd1K
rHaLZLD1saujuH2dDtvXGlh1GTGtGB8WjTOwPnubdJxyrP9jB184lRQO5ITKnQwk
yrZdnQpK1S3bn5U3ZRvxeNw/ahOxGCy0PZviSGdlZpHHvJDOZJv2JaeshGB4gBs6
YzjBF8Sf5m/CEbIeErc+MvFYfQ8xOndNuyP6hGQ0p202pnNfZiWhLO1cfLcTeDsi
F3NuveXFXwTxLrpz53MYOwFr/J9PZlm7loK5jksModWe8vZtMF/kdxlOVx7ynxFg
Mk2gGnPlzAyabwVKvGIHtGNm+2QfAGz9c84hvxHGlJ8NMVWcyq3g5x1RWVGSpvlY
mS9ag40TQhTjw8W7fd7azTjTUBFqqSAFWH5L0xjzBPsAKhvcQ6YbT4y4jqeRgAwZ
obKhGZsmmTAwcvwrR3kw1RLBDcjAnuOB1J+weeAqCSj7mwrdAnke3EfEeQOPsQ4a
Q8p6YRZrLzHDpEMcBEXVUkVcSeXTwZnl+GkGYJR5S93h9C6gs8oC1CfoPiIhIXdV
rCB2SjDcpIZPhp0HUPAesUERFlOpJTL42lBkR3AT8B1tQN9hEvEK14RSj/gLzwiS
QPp7YZ6PeYBNMhlsqVGXur4XPZqPpUnm90ZPRs4emuDzJM9ZZBsI/EypamQSz9Pr
vl/0mGjxjmcPTNIBDZ5E+ET6XqkbZ0uA7FzfEvWZgLKbssmNRcPAabPcqsxgns1N
i4QeoeNZi92pNAVVQ2rPegyZh3zlwa6GzoHN2zzuVphI+rnb39hbZrsS6HfSv4+D
kwjt7BNHH9z/QkaqmXTXx9Mr+tzHO3xw7XfhnfruU226Pw9em9wuaGiw5Lc3Tggw
qOoVr4Nj0oi91HwGnWu9GyXIxXFvSSVgvcln3EMjLYB2Eb9Nu5iCS2oyWCU+EjtD
GacuQiEB70ppAA/JrRo0OYxEv/Y23ZFKRSNG+yAyqUXJ95p28xoeqG2fgccnTBfj
o1CutXSVNzH6Cuo3gjTiExyrGjoduiLpQlLQk0i6V6FQbXgR0Pdv5TWoOK7L9bq5
OLCrPOeBjgkXDJ5zBqVOETs8Zi6q6UHo0hvGNSTCu5FBKz+8bi5uKuex1rjTe1jc
0afoDks40j14dFJNzwtPX8qcBaIYfywyRuFpBu3OeeKcWM2dExNPcgKba90H+RAR
EWlaB43vWJZWSzLf9gluNQwM3KIlyg3yK/DbveIKQEE0Gz0OPTwETfoMv5nj33wF
Bqr8a1NSwadRHMJBcAT2Na6dFex0nocstVgo7SUzvWUEXlIPw8fSEumaiojExuaf
plVis21Qqtt71odhkH4p7MUR/frYYQE7Tcmo/UbjaQr2TKImZGZicE8nUFBzRwDv
sSp5yquhU6IS+ySibPJxGuZhPPP6cYswEjVaUqijBtwKQnIgFZ1xYMCpmI/wMZ+F
cy22gs58AtpKqtHX1+M6NBYn6MnqweEqmJTVPbxFt3R+n5x4VTe0UhzNu+pGEt8/
QNRyPjDcYaepUM68ioFkx6N/meBuwbMcb7gscuB4Ll6m+BGFw3uhPtdle3SiYRGQ
VHVIGvrCMEvS4U9UcZZ9ym1yJ7PvJj0PS3FK6lqcyfFYTg1U61MzhhtVjilLWGcw
/+EiziUGc1+JfvBMv2oerEqNR9FG0DuKUNGSR24G7oaNG6WT++i1HjwWL5+nsUKT
6Synw1bHKww/tIyEGQe45rrPrkJP0IG2w/JAdDU0iYik+Lf8D7HJOdstIPxAoyH2
1KwuAsbifwOnLyiDOFKscYwkiQ/vT+ZQioh1SEGDc28UV8vt7fPBsbVqDTBQjwvu
2QQpfN4XW7iqn2ByH1zMbkOm2167GeCYCzvGdqtLxltfJjxZS7hUz2/xyqzelsiG
N4xC7MVMwcjaoJ4HvfTla6IqqRlEqFlaXyBE3HbOlELlS4/G+eDiGg8oMd/Abq/0
HV1KaQLfmcOB7Wj4RRnmxZMxD/NOJ5Fz6QMAewxHaG+qZ2rnKJGCuIXQzBdfVp0T
df0kBYMW0OfR1AJmOrnxdDrVEBvIiWy3EK/vPNRrw74pgbnrPF15TBT+UXa37R/Q
kqGTZd8HBxPKZVgORR/Fx3wQEhyAq3PRSab/WKQPsepqnUc+GKBCIwJulgLJEjCN
MVrUkd+VO5U0bBr540g4NT26nF8Z79wY1e2hLbRVnJkkPlrEu0Vce/t4kgraplUc
63Nt6vMBqw7pQMMyydJz9NZct4CfQ8QE1b/oHCqUSMl65j0n74CMTxXrc/dQXAYK
KA2J92cto0BtnrpGM7xABCiuTPnQ4hbgkQ78d/Xmut/Fp72LtmJ1YnSbOy3RIp7w
rFf0LeXE+2AxdpwAE723smZYz+JJkOnu7vhaclV9sySIgXA0vBosi8iEkZNf/lHC
sPhmCgv8gPwBREJKnnHwGVpBBLEZODbGcRssvicZ4ztXBzxJHMFkgvdw3n2cVfHd
N7Y4fhFGN+Re2NUBaxy2mCGquDWaG0gKKK0F5oHeh5zUhIciFVUYFZrqq5ZhiQBp
d1XRfFrsAXEFVXIfFE/30w07wnFQIZze07K8S6aUlySy1GdPPg3Gr4dIHGkYmQIk
gCZqTpe2Nl3AAHvxyzujHc/NGArDKeBvf1Dt1+wnlpTq1RCgZu/plWSM4dSOfAi8
MsJ5BYKvyRG6gy7fMGYobfRfNkw5fKH18wTkYl3+MVkIvSAfIRMrJ8qPBvv/YAx7
e4G8BiOmN5MsERlkLuGwhZV+JtIyB5T9F5ZTioTMP9ReNFFKjIqVQJqhVHlEXZs6
olCk/gRrEIvXzVV/XSJa7PVlSGTZzutm5tSkBEkukUkQKoBl+S/EW/Vn5a9jDQuC
CFdDF0qxXq8CaXxEckn2BMVc02DNm0tH9YVg3thnDeaa/sC0FZyJcy6VAgFWayc0
XBd/DzZDW/nf5NJYRwzuSZvbURBu0C7MJ9rJJ3c4XH0sNiQfxH4nhVf8nPhLZ3KV
KNO2vcgcXBOBFfrgQCWBhkAHZ0jCLQgv0z1b1L1y13SXada/Oo1sa2QSbh+qYrhL
WtzS9N7WTlcShytijPWG9KFHL/4rjtSx/pA4vJ8hLG7HZHj08rgIoLir2Bk+1P2N
rt7WYT4j1vNrA5M8PByQ2Z1gDG/vFrtoMcBHOpMsm41VpWmgJlHAFm5sfWgMdEC2
6+20jEYBzUIguVl7iHCfiMv77Clj3Ks/R7eRhzgB3vbZnyKWEIKR4sefBnxBsG73
bM9kRTQZhtGYa+3coxp48NgZ/Y/XbdSqJRHNX0edyVIEnGcQdIUkXCpBDAqEN5ft
X27bXseSDbMuW1s8bksq2/xxYjUTKk04Nj+5zw46geyZNW0CMIUv8ZHvGHTCcskX
1KY68P0cqWoQ3CSMkn5kssG/GFia4Y4N4GZ+Kcc40V4dc+IBrl4vwbBCuumw37fD
OvnP5kuo3sPJFbZH5YbnJyhqkyRrikLurGee7xofZre2vewv56dEFkjEt/3XkzsS
8XNB4jwuN5wCA7doyvfFRJ7LIkz7AP1qgbNGjTUid7hn7rtwdjmdsI84OcSfaS7Q
f1ou0uK8tbJ1RfJk6eV4qjgnnEQE8x48oDxg6xW5jj1FkLdPB5b9IEKxSOK4CahF
dbLgDTLBvcJUrB0dJ8aLY4Qjq/xxJXIouCAni3NSzJ2zHT4cUsBlw/3Y5q1J8MUE
WbGp6epWWn9k8X0KrVIerKLufv2ZPBSnZINgF2oB9SNF7pUhqJRPNODmu2FevaLE
b/zFfuZm7pyjZlPwamLgGjDBDSORvjB4o+VjeLTvHU5e3AoQrdmjpNxmXgF5pY6P
soCGVQ2N8LXr3hp8fPjEL981FmiQaWWNK3HtJjO9R1nnWyR4OpgHwxebPzwBw88I
HQkX46xeGR+PoLiGy0GG4KcYbpnMZCdBbuf1/+bdwLrgp37ag9zD66QhoqA/8aPe
j1dye9Fv0l2wfTBnwXSgE1QAr3ziWXT5xbNZOEjmnF5LlVgi3KzC4SSHldvWaUov
IlUoYJU8TnsS+miou5ULaS5oxdHQzCc1KBbp2HKqkQ1/uVtTWhetiHN38ATT2RNt
LLEyRHjRG7HkCc4q3/72M+ekZYR9IaEuAezwwwNbM5kEiaYRoaf5HTjCxcTu/v2k
UsxYc0SuaiV48yngSJG5yFlA73PTuJXPp0F/zRnt88BZpNywNPu9n4zg8FWQRazA
rJjSD9gXmc9GEd0ZPDup6uqCLI4MaJbE6oHRQAxxWPeUEc/JpRLabTdSmHIZhPiM
M0jEb5S96+TX5+bxCwKI/xQ3y9/h4DKo6KcbcLlDErLrFIjkaBnjldUu3IT1nUWp
MIc0sz7il8eAHjyjKh9ZewcCrAIE3LQApGWI5QUSI5EEb1MtVvzP/C/OUYmF4GnC
VzJTmuv6WpNnCiPczTlv4CSqquAmsqjRybRSZpwzAbdv4n2xcOLlMRK0emoUU0bc
rgQdfzCCC6mrI7CvZAc6Z6Ad2nNghoQxirCYxrjWOy4wfLuI3PkrZ2UwHjMdjCVz
29Ngyy0UhcX8RUj4sX1Pw7oYYuw3gpDfCmV0oRFQbA1w4tiuIhX/8YuTFz1JJhM6
XfwG4aYDXoXlp1yFOCBpk/6P/HpQzScJ/gZ6AlxGPnkIEFMm24blMG4102BuatDt
Jn7o8eCxKWwWbcTeLTfC/NkgQ4eHMHTO9D/kEJG4OWXjbJl0NQNso2r332iNUDsf
+eSBRuQzLHyFfumzKCHloWpM9ypu/T3H47Bgd7zMC/6f5z3d34jifpC4HHy5eSLb
ZBMpmRZToX59PY7u/44nszTHHNJJSTN1GlwrNfdjLkGisp4xmDk5o6s+f70dYI9z
JbASfymm2piY4xTjxXCbr80i++WofLEzyff0KmBfaCrm2BENP3b5KLL+BPU+31kV
UKvog8SZ0K92kac4v8yXpK4+tUgslGTyYMpYrro1HYhxPr4dlmmGqcNV9TubO71f
1K5m6GFwJF/7GRjE5E1k1o+PIFe9jDZbubOyuFmXkyF15yvM2aAsb9xU6m2JUtX9
m+FWvNw64vDcwVqGBxM+7340VYxx9zFu6VxsG/wxkwLpfLdqO0xN6qPcR8EWQ/Cj
C2qLU1S0yNhME52tIbQVmXzOXzsbET65IFX/EKYG/e68r+i3zW3mc5Oks0HesYqU
6uORwZ7Bgj6clXJd/f332MjLhQ5JMLrd52/F0rj+i4VjLytO12ISSuiGJ2/Z+jSU
5j0fl0Ib3s4wE3DD9JiNJAv3SeRhRue4CMGnFYqtwhXlSpTX4PKEb4Uveu1IzXKt
4ida+L3PPYJxT+TeQPYepmI50JrVdqY2WkMLSZX4+8EbtJsh6Wp/gHaUpy/0llj8
4lB2bNyH+OVbIe/OzUliZaC9sBsQ2KidjLBflj6Jtym+kzV3Jo2G4Bz0BpCAoIeI
DUzE6JROyQ/yyKvqp73jZj5ZNw1zOR0Gbj/5R6ceVSTzv7JeBUFhgdO5uNoGu7+A
AAlZQbcnQYPyteaIXO/vGqZWkEiqtZShYejjhTNOfFg32fDMOGvaFlO/SR9gCIqn
cqjpkROArotZ4IcRYa+Qn2Mdw8cpK+4QZmw8ow74TSqI38uMobHFUm7WH035AKKf
u5XLcI1DrX58Ay8ig4xnLBPSeq84t5Up2cyhMT2T+L6oq6+5gLywOhTf9cTv6q2r
A2XK4iI2oA8X096yfjpnQVhCeGt7xN0WfoWWhJ2+g4d9VnF6c+49yDDde+m0JK0l
GlsfKq2kgbKN6Vv9gWnXH+VJrWxBDxc4gsMfjCZ3pCuPnc5AN3vPtvQ410ggeYXL
CYrfrt5IWbelcf/0KznPuKCwPJCtGQ1YddP7BLv5Dgz7PAx9kb5ZcT8HlhXCzP57
3CM9kbYMD5e3/BecuHUhYuZDm8FDtUvK5SEf3oQF9baO1dmSh8ANHZuAGrTT+Bcj
NyV2CXin2eUk6Rz8Jd56DtBdXt/uRBo6BOYybfZphkoyhi1QVNMQGMgk81W8IoAb
ifwpRC/BJEUCLB3ZCNlIu9CpEgW1zSepvIwfaXSTPjk46LUrNwEkVqqjxrUGT5ZP
R/3Z2b66mqwnf1vX000P1jO7yMLoboX3JfLVEHzinpIFLIz3Bk56Hn9c1bKccBw6
6raeJVxEXpHvgQIgK8L4j5OJb2pppUkRbj8BEL8j+rCAKpdVXauTSWgcj/jCKXpB
H3r52V8S6ph9m5eI1yfMWvTrvzM5BmVi21CXUCFcsm63mB67UacxrM6ADnuP6iLF
JAVwMnOOv+w9mW1xGl+RGYKdh4OGWmfP6S+bbbVYZa/BuOiJlLep/mbbRipcNdTT
VO4OLYbQUUIozCYwcuVO1OvjHM5RSCOmAqfc0W5z3eDWeWRCpjJ1HbS55mK9vRtO
aFHiIJ3rqscRLYR8kHRyYeIVryjzripVjLxP5r1hMHnxXQVp0xzpAq3YoJ9WTbRT
wbpmTu/jEE24g27NlkFohtehW+qkH9XpBSzkD/bwlAXA3HIW1abGux+hZIYkGTcm
HsujEYvfD2gj7oKQiQo/NDVHUSq583nEVHi59G/Pa+dR5E6cE5M/cj+EH2YWyUGO
mQj1sWotck8/cgeengyUnfjlPMaJfVDZ5PRj0OKicaa0523mikPnIWHhhOqEG+yh
BNkZE7ey7776WUKJuYOolpcp76Sb8kUWukbSa4SkTcJLuUrlS52AkcNzHQMrLmjG
b/gsiO1DI1v7TZdU/HpgZ6mVLaQe41PPUS1osEl2VvYdM7HPy6k6J09C+xWxdzFc
kYd2GUGJyGBox0dywAvjoQJOH9YM7ir6PzDLgKjB5DDHBBQM3ivQMeiDAyAq8+jK
Osk15fsU6WQXWWegZfHi4gtgMfFLXpM4exbBJYnxfpRLPE12OX4shSqOms0N0Osw
QKKjnhBlfmzPy8XJhlm9/JACa5E8xvfGI0DKVaD6AZ8O9Q4sGdL8ZMQpp06mlTHC
4XDvQ9DULmByYEdhjNlwOgkQWSweEnRRWrwUBJTJXBfcAF8EztlwJhAW7/5jgTNg
u6OXor+Jxc+7H5aVk1H7qSOeSRL6dst2DaeF9F+bMpldwUVQeYMmNvBO9XHn1ySk
Y6cEs3abHnOwvmEkGm9m9qP+40QIyReUY5YxHJAIEzpflKee5nIo9z6EbMknyrq0
OzOoeA0WSUvwAkU7mtVdXPrXE3MZUdE6xCUIj3980WV6Uf/40UIgP5/piAneRD6Z
xEalY30Fva5An4nIkwGYOPkqN755TRbJubuGJW05J3DP+Uw6uGcwjtSzNmlaCiTk
0rhkgT8/JiiaIDChK+lb3HCH/qzSqt1Atjv7STjvwo7ENCczIoSqUHbIzahb2n7C
vfSDhWFyH1ifkpbPdNOkwMlbv77ML6y+yktFK0X7iixghJ4M+SAbnT/NW0lDCy+o
lkATmLf0+q0utAvTDVTKEJ46ekHlsIzAS4hze6ckHNvhg8nP9We6kReAcLlaBQJd
D+DOwwGWchfaCLd6o10zf1zBZJRoRmKv3l+7KQ25JpFCb6NIKduCzyUMKSncYeFp
9tEDfoGMvh96NI0yljtK9Hpy89mkCuqJVaAYJ1KIy4fTTN9QuhsPyP8wFSs7fndM
nkkj4vUVywLWEg1erzlj3d0L++PE6t5hUkBNJ1066DB1O50SsgCIH96P2DmPDc23
COeoEldkHyXfO0UWEXHOfAZQFSr5/x4dkcwVUYvB0ERNIoQniTB0Vai7XXQEhJBg
q+qoCqkW7xnRkWWJKmbgGFb1OiweSVsFvH0Vyiqy8IFAHvr/r5IeuMhSymt1agg1
rcHhAXlszUJkOwPefNSmlMtYRdZqhasXjA9LW3UhEaGppKmBta616OJePOopOhiv
mZLW0L9MKFqAn6Mh1s51X/B76MoNkzjhtOC/B6e64CY9oanBlSJNdaSIuJ1z6Fbp
tOnTcsoNcCYGGRMe6FEZloQmLKZwQFbr1gwCAN1SL61lJfL3jbXv0KdMLMO7oj1R
s3d6zg+424zIbnXbRv/IcTDcfNiO6mXMS8wC7tvo0uaLmgDNth/bMPhw3oNivC1z
K6dhC0e/qevTU8Rw5LN4Bx2qmQU1iu583Wz0cAe9a5nr7eGMWVJTyNYsKjAEgRq7
D4vbDXzfIVa+7qcPs07V0EYYGOgOFIQpwf8GmK1PtAQRhVGpMBNTpG26Sd/Gzqa3
unPRr09u3xBp0VFFZfRB+kMwrZfwVKcRURIEDM/kk8Rp/PNcwu6Run8Nr8v4u0Um
O36QPx1hpuPOG9AdeUyd8APkjASJTLYbK2OKLbiGy4R3PyzFB0NIA4s7ZwV2qOKa
MwhcdN8yqNrKXCwtx1chdxv+ww0qeI/t4BBHVnzUfjGV+khQPow9pW+hoFPDXs4n
oWHQklADGHhkxZeG5eHt1akR1Y26NnWj1D+OtTWBiiHfYo0USMqebzc2Dl9i4Q9m
vucrgSFixbFP5gwJPsHftmHt2DCeIa7WpT5f4puApGsfrcUUC3hy+CRsl2Yn+obb
R9kllDKi3ttDl4tG6Kn7zsJBSRyjbXL9V4SMIvcCuxpi9BlKoJO5+pr/+hmP5dG9
fpA2LQD4E4sCF2MBV7tRsOQ6pGEOTq5D/6UvUuOMJl9swqJVPVYtN19qrfldUbD0
RbCCPk7cAniE0x9XDMFwRO54XU4F41Pp885F7SLASjjKxs90nmH+lIjIzIK/8Dul
tCCGqHk+nspgpvdwFnTFZ3EzvQA9VcRcZjCLgixAnBlS76qVBfV4gT7HC/sgvfIe
phhXWcH21xUEo4uZvwZspS2D0iADNVi/CtAj0scQr07c4xPXYbzHQMk6OJiztIfj
hB/eiHj3unrnssZVYWoGufBQpdP+Vb0l34t7PgzRbOXbU20mwN8OIXjHfv1asNsE
IbbW88pbH+hd1yNvNVzaATfunF6lCdmYiOXhrsZekakTGhMOYM/qDroCdGNE/9Ou
tbU9D+kXWa9ftd8ULTxshZAP8ClwLiT+/wM+GxwgRtAmtV+p9owInVBLZ+hZ91Fh
kiRGMq1qK6+X069bmurnBrT+B/1SnRnO7NPZA25CC2qN+AQtWa5xtDhAnwOo9MUG
juAu7LcPFyCZJACzHdu1UVd/dgW/ag3m0+0I7HE06+NMd9UE8peOIEa4yR69Tzgi
4ZCMoEjXf7ILEcR4CgXPt5DOURecYagbuGgyB5sHdOOJ64dErLXONUbus+tMWaXW
v0sH3XsuRwlkJbAg8pI9OKSDZL3I+7dcaSkOj7lRblIZxVh5LNvExUCGI4VsJvjR
WAgviVe6BPXdx43SPSFWn94Y7p9krCuikF6PjQk3kcxW47RhNpYMlDu0cvx+gMJQ
c04OlxVTuEdLsFi6RtWWwVfAcS60MpGSnmSF7iwyrHbD1PusZ7iz+sG/+XFK8jiD
wv28FmJuqSiB8JARbEG04DnaXm/JGNWNS1/oMUo3Y9n9OgfwaVU6FUUJg/92VU1C
Aj73kbWY8XYFf0KOAZwHuPFJK3qHDjK+aCv1BeobkUPk54f36O+fYEZLoUfRGcv1
V/V9rrjoU8YxJ2GTyIfBH+Vm33m8LNUn5Rl64ukUtROWas0nCdQ2Ydp1f7p6s78K
bHdWy62PyEXPbAyu+XmbVOcQ3fjZoQdGvKtIScdl70YpAEDgVuc2VmNGo+4pcm/l
zO0XKSa6mw9akfxxUqpKODb0H6X9srFnmlzrvo3+2YKcza3811BAtHVRS9YaBpNS
0ClVOKxRe1QfWa9tUGJwPyUc2N8eGTdmJcOOZeSdsF407wl7cmmhkEqOKJpbYJtn
dSIM0qmbJTSVYu11X9mo2MDoxAabMgEf/XiFx3qrPGIxt6qpEr3UhUG/f3L8t3E/
ao0RGuB893RKwIpl/caV40oVqTUJyLuYH3UzwVbr59ACLOy6Uls+Rq+hLYeW6mdV
K5gPQbHJQJt9+nNQcrKDtnNksw7t6+edncrVVJDroNTYI106dI0/ABDh4TFu8kQ9
0t0+pqWA8X/nof1UfSZ0dQO8EpP2QWwZkbzTdxuJ7bG2ywpJSG8aht2PzYO+D2dS
6rCsQy7j+0CxxaEg2FWjnfK4/aO6AdMHFyx6rofdcbUF3jsbJB2q0E42r3jjurzH
N7koBn+WQ2wVW7Xm0TJwkycbCRdIMl5ecI6rhKr8JOQHfHP361ZYIRQpThEwfvll
XO3n9G9fwD0AdQi7E8ZPzKAvzqQcqcFu1kEFH0ISQ72l9kSwXSw6HuDXEU21AKw/
6OFhItjLaq2LWuGx4zYhZHJcDlF7fMu6PFEhYn8xe19wmJ9yigW9m+9MWQe+5W8y
WeZh4ye7WZOBSSO5/pxGNmx7cFGLZUbrJmW/z+MXi86WTnt8vnW2Ps5jMhywtK1C
Rqt85E/Y1C4EvMIADZzdog9Ln4Ecvn+IiAObrbzGRljdp+nH5ClDzwrRXSPFhneG
r+E4v3PrdwMZnejOK+LddIPZDpnsrvdhsDaZYvMKHSdvWbG942NyrY69bktjROR6
vVf9CpPCs2C2q1K5i/F1atpEiZjDCbHjGKvginEGF20TACmRDoxRVxIiabqbtxWm
d1vOOjheCiawSaIsSa6pMNlbxYXM2y9iXTzgb4hbcf8yL7Pm/BFIa1+MaZW1mKb2
nhTupwTd7WwweJo80MazI9SubObxW/22AuPIVP4jbAVO9D8cFrsTnoTnUmeVyCN6
dgbWrVwe7i2SGC7ZdWEM0n1kjjto07fK+UPONX8cI9C9sqdP4AEpU0e8R1zAR1sq
J1SUNEvaiyeH98bXSAsZHLBPRDW4pz27tCpPZ8ajJg+Nz33VpG0WCrpXg4549mii
DiN6NXOTqdehK3jPWoX9ABQVy3IZJFNRfzQJxaZlK65arDaRYhWpMTPJVCBRpQ4N
HBKELCQLM9siZQaF5wshEu32mAL5YqNR/gJvEd0xKRvtOTplH+jjaJfxjBDkrIzl
Dculonp03w1IG4xFurBHcPgOJ0rBkoGUvLjOpRkwo51ivARvZnr7tERJl3yiZOuE
RO4n0vjVZq1ZGpAM9nLBWfgwnbAXF8njoaSOnFEek4s+V0hNDAa2y3hD3BkMYl36
idduep7Adm+MxoZkF+zXgqjZf1po5qX/1WGR2eADt1/zJKe/IL9QR4St0I33pfvl
1NURZ1mKXdC3X7hK3EOkmnAXq+aTPlFiWwWRCLGwdO7NLhh92UX3zN4lGdY53bow
eArUuDW+nqDM5488C3gIMe6wo/kvmzblKEhQfs6ekFhT1LipIKcG4BNr6u2S4Nku
FP/vnnAcB6lgDgPEiRjqMzFiDo01pctRk8l2CL90C0Wk/kv9MyjYuaaIs6gPbyPl
dz/mqVdwsUZ82rxOYEFQGYa6R2iHvbj3CENEvHO+90jFqRDwNc6RArkMuCWct9T9
MjIpzYZ/KZAm6WEoTuUOwHgcgfjC2n8+7ELl/kunTMXuf/w70CC3vPYqYa2yJ5h1
y+tzuMsuc+/Jmq8UAWZMI3k1ICi7QoC9lq2WUFdJUkrc6UtCv6VEShakDIAaTdAt
2c6SmMMBcAR1d75P2/YfWtu/CIOu05joCeNv0/tH5EcmEk8hU9yuQEcJyYte8Gyg
5VNjcH8BZillPk8LasVzfHW1fysWuyCLl/bUJ7gK5u0UtWM52H7EThMvWBccSBlR
w32EPwk/QuaiqJYACLvoACB527i8UCTLdxd7CpoXbqG9CjTABA/tWfOkAfwOO5JM
dwi5c4Edk6CxcfAN1iho3ltS9kWyEL47Q7Ej8ZN7oaPSFRsGBanOENmJ8c1Suep8
6hT5MbCwvEGqMrzRDVcTpHPHq7rTvOj4CFS81kEQmvxImSOsJl6mN8VRdyPXxaUr
JsLp0Py1W1pREvJgvcAkd5XrNyl/JMT/x9R7gggPAFM2mBj8n7f40LtJkYkWGQlK
foPnwIRxap64b5P3H1mpJvKbntGpqBRUZDddns9r6Z8NjJhb/4WVk25Y/RnTXT7R
BCVX++JQl465DvRF4ffltji/oiHNgDwYj6oZkwlZgmH4vHftW4N1aZMc1Jye6alb
S3hvAxbniwF6TgBTkzg68n+DfahMYtbP+G7sdIT3xr6nnTrUVK2FDs0cJ1Z2pl97
ukhkRU5A6jX2D+K8QCXPtuopol1O8vafv5QaFWgjxAyNiJEpqtmLxekVMR1oe2MX
yGUUVnMKAAibUasvG60anrd1GFRhECYs+y0aWBYBmacqDCJUOyibztJzVK2hbS7H
TMMymgPoFmYixTyX72CQhXWOnrKfkABv4e++HsAsTjl8T7O4kTgQJBQCnnw7gb2J
Y2lwt5PdFxJx/LAvgO3lqdGCI5S8VBeXZmfl2A7HG4e7NAIuzk+lv7EaeyfCp2cc
lcqXUQepl1WocDjPz5iSjGLG58Gu9870utY6J/FdmkPEumxAITxcIz11cpNtJ1DE
ApjJqxuXyK9LQo3IzMCAtKD9MuN6k6bosfSbh43y6aaZgFmBzts63AjE2pz5jFNC
x57GFviUPlMJRpaUYL+KpsNAv3nuc8gRP6XkErO+MFIG3o1ReVX3Dm5Fo6828iPj
wlvbDE47fKdwAjl+ofpTtpK5M6hd+vNOSjZBbW9z7wTVbZ0aEcuCPoaqoHJD8nXm
B0inx6RGv4NHXfksJTrK2bFSR7qKeJ8PYnGxFuxmgLG0wZAHTW0awpYzUQsbBd2h
RmKcAzmNhkvSLEdSdVhXBXNb0B4XTs5lIYF/e/U1irW3v695UFB/dEurX/6ujX4x
gFwoRg1j6ykcotOSBuIrrS+auk2IjmttL6/mhibf1M1h2EmolbAx55Xzkq1BvcQ5
cfMhO0D/KFIoYr9hBdUhRCJAjKizlM6MJCSQ8y9Ln08W57BvqQHIZVAttnLV9GZm
kMxM3G4KmKzNPLBY5mZUl/xux6X2X0mO3jnSmLnPQj/Xn8rWaUw3Nd6qOIVewDnX
3ROb0rENMGoZ/0KAp4IB0K/aAXxDWehKMijcsBw8p3q/LbkJBwC7OdAsd/sZ4btQ
YE9Y/mPomhUZhYN4TurkvYRW2OYmxNraOAX32QekTTW7yVK15nyelrFtJ7uOsIb0
gya+/2cO+0MU0jniJ9S9V16ENSnvKhxM0oM8ucoBNQy3Vh40NXy9B7Y/bY40p9wZ
GbKJ6Hft5+TfPfb2hUFBNPY6rI+9ONANanZmzHTqRG5F41tlk4V/PgsDB2vUN3e2
J4pcpg8OMF35tJ3KfdFwxp29R4abp+Ic3Q/5p2TtJTFjq+INSDI8L2d1kjV6mvoZ
ay3mGz5iFDLhGevWLyTVsQML/lJgPEjzKwouSxmBh5nx4C0OcBsPf5BQH1vlnePG
O8ScL5D8XxQJz8+he42BbKTwt1a+t0TjhnHkxPT1yaXCMzmLrQ6KIiDaWHtYYOZD
s/vlqAbI0gK4FLaRKjQ8OEGZZjP/hXD2gQW9z6OenZtguzAEz7ue0rQnZKNAcEeQ
M/jU1xAYTY0z2LflBYWxqym6KYRDL5Ht7iDzPRMzGsCTPDzK6llYM093JEMLS1t+
FJg7y+CYCfjo1HeWRDvwjfA9DgC5OTVm3Pvns5DjlK85q0fj2eJ2Wjq7uUCxVFC+
qaC6fIQUJscMGJeLYijBrGvuD+TlewVlTOuWBTQoLqoNeSSjCKshNfF2LijlA1HI
SVYC0Swe0odvNc/CwDBc2yTktek+PfYplCUN3RWqVHYGb6DsYcP+mK5s77j2vdct
5e+lujYQalaNbooDiQ95yRsoSZ45+0OzXNTiOYbk7fAt3uwtlFe5GViOHQOfUtfI
CKkw7silvQFlWyK4hxyru1k34/IftyZ1yGs8yZye9YPuHL2EzkLA1nJwdlqZH+SK
pb54x9pOgjmTYsCnyhbGuXUFT2s4n+EMP4eKtX1GNYL+jASA/3CT7LxjXhPqNmhG
NXVGiB8HKr2nZsORL+78xLGXyVPzsL+ACjL4HNbNzd3nhLqcviutxk5YXtht9pW5
2EZzaYE9gV6VfJDfKAjcjjQ7NihdebNVIPN+axD7d32KFPWexhaAS8iwjsnS/b6x
MO2/YBn54D3ceDoZ5eIH2vYORvMuaXgJRvZRd+hxxJBMGCu8FLB4ZLVI6EhMidl8
B8rYNZwYezSoa5Ki6GFxq8bBSYpgw2oT+hP98tiqEh8VVdnA9N/9/eWBEMvysLja
XAWVWJze2WgriFJfb/Y1q8MN3Ub6NvpFRkxrhuRiclxpMNZ6dJkkMcfJWc9R9JCT
5TXw5iW4hReQuKB1xa3VOTBDSMkX3lN3mu8hu53hNtWRKU1wkvVhdf7Y8WNHPGwJ
aZ87MRcbNxT7Id0c1jK0RzAcrlVYwUGd/0Sygc20F4LhihR/QeU6YzxcYey3qCNJ
ez5Dan8GD8MvB1hGD56lQUKzOGuig63QPd38dlMhNHHJmx5eACRpTVR2x/CQJSiX
Fz9YYIxbjnJrkrR6VR0L7LZGc90erSNfftSIbpKEwRRV+nO7ysB6yjFKpnb+BqYq
ciN+nxGmNtkq4ajCquocI+cDNf7VI85JOU+rBXiWaJUOJqLEgVCzlBhSpteXZMKS
LUSEt9vnlDHQ8ET38lc+AGrNJ3CcVlx+v6gjolwv8lrmUqSm5mkgUbMzC9gTVg0+
doqU1a7PyTlzrz366QiCyzlzZiCXMqGB1TgwK/zXAjPdFQWaz/AOBkXYZvKayCSq
6l0JSy+6igiwKchkoSHZS2+scfYNFXutPQE9nGktdys3MdFSm/ZsaC5h9t4c52eW
4yn8FZ4Z1zV39e+YSGh6cYjaREhldhLhxdrd3O7iX7UDePMYkOgmhkmJ6vWUEBZc
UKPpdPJEpwNOSoy8/cYKubI1PTwoFO1vpwKpzq05ANCt1/a9yWQHwIwGtC6aENxX
rpSwaN9cVn9pvI927Vb9Jx95XB75z71TZWJgNAI+L2oK0GuntRlqT18jWEhZj6kX
QPRwscL7ZIy9QAxddR23Rgry+KE7VD8rWPddY8UgYpMIaKrMfV5TX8GlSmT7163j
dyj5ZSODj/RfPL/Oakza/YwJrPmXiQwPZ6nOe0rtUqzpMGFuMTAbluQP7E5zG5D1
DvrHjtY47ThFkCv6YUAmNAoH+x1vMvxlK9jcG7bLnycXcLL5xqY4edq31CqWeFIs
Su39twiwIxxWpmF8Cwo2NjdekZtdYVaep/4XL7AJBmbRjddCJze6+IW8rWX6icCh
r4U6RxHpyMAJi6iB4+rBNc+kC702N6ICdJ1xK0tprHP8FfW2Z//hnNUa1TyTXSm1
o/8mbHH95IFjAZqdRi0Q+32X+rM0LIbhNR6cQEo07eg51Xy7tDPGVC5YWxr3ASWb
zhlMtESJJJk/jXKXgGAZtKxwXekxAZAsmC4IVZWzCCokUrRcnD3K+PSVrG9O5l38
ZB0o3HkYp6lsIqEoPV09TCv+GLV+Q7CEXoQsIEa2VJ5PqhUfQDstYWq+gAHH4nhj
Ss3ga+Ax8Fc/Um79eKuo6uYmxEMcWGBatDJRQZ8Db+EIx0NSEUYEz9aK8dFJnVj6
ICtm9KDrGfCYgE4v5CSAV7tWs9M8CWLuAECNowJ5wjd9KgEtXcxzMKYDWXZS3Bk7
O6ypGeJjcCzATgOKYe3mVeuUGXPLbYYXAtou1qqc6bLypfpCkv+JSY4dAtCjL1Ms
2eQsQH/OXHAYiWJopcC0hVFwdRZT0MtFK6flvZ14mtKOEef63mC5GN2uq8p3g6Wt
dCp0R/+vgThJEaFYYkr9mu0PCVuFyseyXR29pV7/IyHcGR18tkXmA0gcMCTVnL28
enNnGWt+hC8oCZyZF1mDD6MrMdSkNfZrYYOd1Zo9Tg89pBcarwdWOTHL08PDyq35
LqAjLt8XNFuhEWxIenjZt/8mxmuL8QUXJOpU/aT/g3rNkMtwnIwCLK4lkH6T7zPw
XSzljAVPUXz+3fKFgWgHOlLdIVAX8ETrFgNYD6UGpmZMpzlA2aq2ZcdQRhj7vEHp
cVpaU6Z2oGiDBuKl5io6KU8blKJ0IVx5BTWXqAf9M6JuP/BgXX3kj7ZyJ4Mm3a44
7/sWl3JfdGn8TOZgnzRXjrS3oNgZEhZ8lNNlto9ViiW9yuqv7d6TlIZ1rKO7hqCF
NEVKZG7Q87KnL69KdNXajedVLFrjL+4T+QtTEQkTxtAla8PM6waDBj9d8eUTVfWP
GKZgvqq5FU7cKyBp2RGYB1UHnsZdnOhWAlZerFHfn7hkiHGv/Ylsl9//fdhZooxp
ATvgjaQJxLB8smJT9CgfWLODns6n+lwrCMHF8a+rbkEMkydOtFk69Rk6pt7K/Pum
gVmwgTUTtIX/bzN6yWmJ5zbagEL9r46m+L6FHJMszTSH6XkxEri+uWNuYzR/cPM6
Qeoa5ElGHG/gjEgExpTrNo+4GXZRTQ8uPzhkvpiICVzKNwnpyPMhtQNSK4LPC/Fo
crhMilTJ0GtNStG7zMbiGgzy0gJkU+G/uwpmKerZ0NMwFh0lsqDNbMGCoyBzbd6f
jX8ArKFA96S1lawhnSn9JV9URW4rACXQWcNnsPLn7znhfBH7HW8JLETcJhH9eOnV
369uvOzQ5z6B9z8h/YeqQXSaxIQNRySaSCsbgRJ57OqAZTFNFvSaZJYHkiEQBz44
LiYyZsz5l8KgbTfmTKz1w3/+yQjEtp+zwe56QP8hAHBS8rRSdrnBtOeoA4qDTR5m
D8dPW0PSUA3w/hJ1m5MgMh9qvpa7Nqlfz/YTervZVjYl1iVb781cltH7/cc+bFjL
KGzLGvZYEh9ViHMGn1XWPhxzLn3T3OUGQDTZHiV6Y1+8cXO2hIXdeVrhdyCYYaZQ
xxgMwc8ZhdbH8jBHC3b4QgzM9jJ8hSe1ZTaa2v5RSVaSO2y2QqVcZqMLdKCkPWnD
IRpVZAQChp+Qj07j9+Ysa6F9tPJEdnDUl0yB6zvpsAstkEhLFdpUrAAHUIhz62Wf
txsPL7GXzOjqBNtYVvEQt0dqP3sqPbNjnIZuNkh1vb+1Abk0PmHYsWvMqGCwFPlI
6WHzHSKgpu3DCPYWKkRV/1BB9oH5e6BbkwZu7oQ7ja0pgcteFHn4YuNbiNb5zoNw
0og/UppxCqAtn58VQQ9rw5hGfo5Y/HR9PkqOTd6jGxsZDikPIewJPwtMO7Um4wyb
mAGGqnkPu6H93TirPkn+TlxQf7dA4HTT/w8PxT2dQrTx7D6hvtS75ScVEQBnO5E+
jrBtD1xA8zNDPIGWnQOrwUTUcNfaCKgBsFcGC/38QaE0//iY+CEvDSU+opeAw8om
1fHCB2yJrgivlEVODsvObG4qAZtHdSBgf9ucDFtHV8hMnGWzZE9J18aQ0eS+T66t
QptFET/kK2ywE/C+mulb+Oxh7mUQh2BclB97O95kAV8hpStCUvCQUHJTBVidVXBs
5pZn9id6HYB5ni19jNDb8wF74Cu68KSWpeeG6CbFMw2O2wlYPW2+U1ZUW1nB5+w4
hd53wHzZYwinfaViEFkWKyOYabYXixlPhD0r/hSUyBk2bYwJyUTlKjb/Hz3/zTxk
LGiSftWRlMlt1CCnnMfV8g6EtChj8HJms5V4sWJPGHRrjR9tUKKjZsTkrz++w57p
l+Ds797d6amvtRvlGipIvIokiYQH0LPlfjDY8hkBsjVk2dLvOBFEa8pWpqfhhjMn
yfaRzJwlbLfTuq8ghQkmo7qE1bO2iHqV/KlLYeokgnpA0ez0+6QsrIvAEE+57AAJ
Wqb0e48TvR0W7q3UmnJFZ0kk7iDaNMpk5YeEgw+M+7J/iAhPjIaFWYrLF3xIgKLo
AoVM3/+zmpFsJelBessSFXk1/OU24IHfowH5hcg3lv9K55n4dpI6N1sc4ZU6/kgI
q2uUW6F5rqHq/4Oli93OnWvCgLuezCzasEBpBzXq289k+h4ko+poITd5B5j1Zu25
iWMF1/CxTthjDEZf9nX2AP7Vd2c4NslZvHXPe29bmIbYrYjZsOAjzFA5SHPmVAIX
76gNLA/5GgWQgvor252DOfY/x/TdEEJf/2tqIu+t4GIPZZw1J3BXHpdaxQ631gUS
nGAZyNW6qLGo2tVUUzeXNZPhIIusgo8YizwQAht/mpEIkZo++AkrMJ3WSwS1McYF
ZoNQD9HNq6gKmp9tOXz9XToOyff/Iria54UvRqwfHQKlA1uCmzYxF3HH4IDXhpEh
pNhptW9Z5zHiuqNQZ5reCSyow7sOrIbyqGM/FUcfpGYTfiBHDc+5cTsTkKrZwvX4
M+60PlpLSHuFPnHRtYkz1VWi30wIUg8iXoXps8TITVZ/H9KIqnGJZNyuVS7sDyVe
0m4ZSFGf/nK29YHDBNuYc8YxjIPpOB0MsW2ax4fryINpdamI8e9tPNYEmca7Gwhz
7LtWuFH1qIqGlmp0BshYnUC5gu6dnV6p36Ipcv5Neoiiof3tqKJDeRCO5mXwSGEG
2LMg3Fc4Gv7BX3RklmdLzM5hTJUaA1C1eg0n1S4DpVHP0a4g2DIVa0cb0prEPKqq
78gOz7uZwpCh9dqUlY1xADRZuBgQ109r6Vmi3P7suwh4hP0YfLgxxNi4AA4nXnv5
RGpUASN0VJ97SAGsad7A9iyld16aQSfMvjVcDCAX/kw2wNiCsCYymxGTn5cxNPDK
imn8PmZuaBkjFWaSApwJzHLSDdfsXKa6lE2UwQyqDg98CZnhamT6fhVVzy4iu5jf
APcE/8wnXiPAeJVfY+TiocMxUSzgJHKBQokdkcWnTOpSegac/sPGpO57A4t839TK
Vu9vJDIBwLi6KH9Yz31gpZhtxIEaOVorXpcIY89M8ktirYEUkZfP6/dizPBl4EnB
DToqLoatbRFx59/OXOUrUc6CvcY3yn2AwSP1H8YJ63xaowVTGWf9aUrD8okStegI
cJc6Gf4WGtjKnh4hpLPgOuTEhGNW7sBkg98Ja1Y9ub/QrNHeIja5FmnivfOn0yx1
7STdvmA1mTK38OW5Eqcsa2lTHeCFSmoG90at3stz+P9TqJxb4gORcbPnt9i55vih
AJPQzzQxIVQy/mr/B/9a2efaFSGUDaly4twg+lyNysQcY8eXMnyeUI57WXvDIs6p
ofsueyzh/59d5DTUg2++LCbWwl3zUmqUa8u3bhEtj+32wYZySzmic5MnD+ISPZzE
sMERMBeSYO64Z1Nyq21dEOmmD2kgTJVxlVNaiMjjEdQ8zS3bWwGf0N4HUUUgS/Nq
JHMhBust/dAOhI/rfPr13L4ddTaCwN+pufApOyQxXiIADVhsOKSe2MSqlkbaQPc8
5vykBSv5YU3wROTK3sfX3NFyBO2t0bWntl98P0CzxyHAZV7lhn3FFfKQaH4sCa4A
qvDC40EHJ9+jA1vzMRk6rZrJmXna2t9yORMVTPX2Cu9HfeoSfhaylkwoi1UBVhgR
I+KpVCNAhXU1Anaxw0Qh3ADwoLaiIgNL6qopu+9oS7QHke0s/cwo8lArRAmKvDnQ
DybVWNJNf8kuRoJfLJVN8oZvO8bCqygYSHI+sNlYIuvE92hOAJp/xZcBxdGwrGxW
Gh3RFWL59o11crwa0sCmtg6/6r7NcmEg7zUfTAPF7PbF/3PmxkMylXPK9hzBzIw7
E6ZXPITpjglXEDjzieZRDJPoFDTOdG7BL+9VDJ9VNiUEf0xrsqznjHuKNMielraY
V6w+ukld77xPH7bzm7zAsz9tOyioq2rRyoYVMeOq7+2UgId4bnhAntagB1XYlubq
jlPqeduvFuk5w00u1AbL5H/W4jo23ClH3eur9S5fNUoYHc/zjkQpqjWw0xRi8jTr
+lXAoR+LPaiO/Uet5aRgoZyVMJNKi48ki5yhgrffTkml2IksfzihHy3Shw9bNoZS
wctCz9XUcuBqNVD08wFEfh4WHgzjH43v2FjqcOfnlryqfYo5sDJtJ2yJiSas8YFq
cUSDO1GXCUFVeLZa9zhSrOTvJ7GyS7Py3xwWchDVebynUBANU2fCG7+MUV00AsYZ
CJWsjpKU8F85mj6mTR1nRkX7k1qq1hPpDuEMWzJ+64IsxXRsZj+egBIbY2DYbqSs
F0PQcGw0Rot215+tpKyU47nZGnAyRvS6AaLXCwUpcIWeMoZE85jMS3ZGL9RUjydX
g2mMPrfERC6zvpxCUWmci/0KHFZu3tWx6RYWi+Ack+AoKpgsPvg+l34aZ8PIBBZ/
+jDNUzWqqMa/PdKvbOMnMyW2wxJrdAvJ9bwBU79N59uFTXisk4+nb2enoAVhmaC/
ArCJyqKN2e9e8INJNnMdxFlzShhPPQmkCtSoeLTuwTZ247GeCRSe9vrDEIhuT71d
7PESuYK1vd57lzCbzNbHd4zrMgP/F/e3/ifcX4HKs++BzVf1+fwIw+H4wb0MpSGG
kPfUhzhx+I8gPdCMUH1VHh7N5Sfk+8RNrHfxzU6ksOkerPaIbH+WEVsewju/Aao0
GRsRCIoNg5BcjURelQANvbIyubcqrJ127pmWhw8gVN5zKCIyLsrAjk80jSoPXwCS
Cdms4Pizyad2CaoLyKLWGYy2BzugEoMhOj/dhHYL2TOeSqNnnSzC3MzfRKiSyXid
x7uBoyJHbt+UUZXn9WSdZiFk+4J9EP4rouURHfffSB/MYbRBMpmlIbidvA4XystN
Sg74yzbOg6Pn+zkUL6aVuQJcbD4VZUZXmL/NvVSMFFW6LWDMoR44d8CCevplCWh7
IKVsfr7coQgEuVBlF30SVykFtDVbWWamj/PmvNEJwW+VOlvxfD6l0A2BhFJy76yo
BQ3c74GdZRExnDF7M6uULZfdzPiucp96xQsEjdDNaRMZuVzdswq8dpYEVsgjC4ci
oWsraBDrXffaMGYBNAaKHEvslj3EF7cOFsJFoaEIA/PsM+Sx4nRDsqkTS04graxk
+WL1R7pzkYvt31fathpVMhfuTTmMo6Viyv/XGkNxuT09bD2X1cffMKyFfW5u7y2N
KzKKk+Asyr7To3YUxU0NEMf5zevHDxFYkbpHLpfX8P5ZYzxKFD2Qf1ueVSyIl6Ri
2RfWI8mcOjJdVXehTAVNT21SohrPH9Foo4q0V3EsZ0Y/eMvfWzcbTqSxnizmDeC5
evUAjr+3RSElB8R529GZA8ppe/+oZrWQFjPgzKEJz3a1uG2bWa/Xxsi5KYOwmiEi
f22Z4+UmlQdVZCjq66EwG2MewzD9XYkGKI8up4s6im4rOmAPYLTHfu665dHyyHWO
1WYUtapKZrbensXOkCgmWtjVAjVQmh98zSHUHBLUorAJ77la+NZfPGyT9IB1tZBs
QSQuc4LnAv5V86UA/u46FMGZ8njPuZOJC0Cg9kg1HQy4L+VDqb+maoUqLt4rbzVA
L9H1edhlfVptzhOYgY9EE/X5Sj38ZaJdcUsMA86czd/VO9OdO96Kc6hc4hcVQp6H
wFeYvMfupifV7U3ZvDRQInLb5Dnzx/21y8j6u6kBurYLvUAiUUZC4gHi7rA0K2XB
Zua6bgCB5tNNH+jGObFP1yWutNRZmkm6AXnuAzkq+bYH+FkoEPTxT3UIKJmxpIRk
WPLReVqJElX4Eg3oqGf6BrvcQo/a7UxFq7XibselN4uY2PIN91nTvZU18gnlwt+T
CyryI+HqlA8gsph2czKzDGrc6H9TUX1OOlBYUNYdSswb32ou4s3Ba81N8F8+mHNh
l4ap/UW4VLEtZL/j8bXWC10+vetFrvurk7dZewENZXKIxWarQ95KlVT94IW8634s
b8DofcAgtRJagPC2VrE3S0VdA/NEFO0UsEDn61jfzj3GJso44bUVBpK7SJY3rbVY
bwzwwszew0MWMsSlBUH8pTSQCvAcfOwV1RVo5OBAKaTRxqMqB2ZWiBUaJlTkuUx0
c6i9PFvHvzMOy1R1SAfihqJ0JLOZrWX44SPA7C380n/EH40VCAr5CopP4ajNaCNi
UWFSn7KzZATRfdXvhZyigWhalXEQOueseZ/IRpbxU7x52+VgIlq4Y4p86c+myOcY
C76/P7FRe8hwJ5N8c6ck9TIgsi+xD2UdfF19nNdfw2EX4wL6P52CrJPT10rM0wYP
BFuEr8RwvlFZo/Mli6EQ5wDlnaJOoP+9pHgvbRH6ZRtoz/P+/Zl6llLol6ktG33U
btOlYdZ6HtOGrgKn1BQa7hApHzf4Jqd8Z7b6U3JHcRe5jwW7kxXFZpId5nEKiYfu
VfEPEeOpB2RVhJn1nkMqx0RLYGXxsIKcJb0EZv0mxUIfHXUCRYsUVseWypnRL2GE
08XouyupRbeqnn9DhLjPg2NnOv1g7AJev0l8cj5eWxZcwx1AnMTYWQCTjcEZGOWk
Cp6koT+Dep8HZkMKW1fPreRZth1RYuJ38sD2yVfkC8UqcQKOf/ndXfFvjg0GEmcu
RyI8aVnORbHFhiGEMu1HzyIvAmqbIhODBkQR2bfNhTYAF8guYdiK/IScnTKeP600
uuhMvobunTkbuy4mLlTOcG2XZdV9kHj22e4TiaE2ltF6RUr7wosRBxG2Ftbp8Yea
Z0D3BZsMiZQT3/EXVru6eWoHHP7TBbELdRM2O68qpCf32MAzZNcqJJZkA6BSl/if
ZNFXQ12vW2oejvDcPvoKHM0Orpyfz9anfZi6X3PMo8cmV5fUUCeSjPE66EzJLDhC
E6lM0RoVlrpnfwgrJwtiKAK9MYX4yc8rMtvCCDCf4ZH/MHmGsnfDflA//869m0zY
G+xm9QuaPwcndS0gn2/BpHcIBVZy/CQuqubOonuVPgWwyRXbXHJUjG8hruy+x6PB
nZyCDHzVtpCgy2DugfH93o07g5M4gHdlfEXKJzsvNnXumF/09pRaew+wuQwkLedC
aJbjSOFBdoydkAn3IlOjsvJ0M+6anRaiTZ0sugUtFINv/giZ0TYE6jphnZpJkx6X
JyJUixeMcBUKe/w3l09COZXVBpM5YElUUAHtwtp3//sngeWfJwRvrv7r/Yuap4Yb
8Z46lRK3tJfdheq0abkJh163pMgO/GS7w+HbAYdNfHJh8OcZcV8SJscPSXbnKA6i
kWojLBt2ZZYbJjRZPbJyALUWDVHi/B9A0e3hhCPqhCn/SfpAmTSlSgpWqUEoqQ2h
Hr/SLUdPLWE+T2V1ye4oQ1lskmWJxmluaHUZntbJyJG0/ctpJic1/CwHk5lIYifV
GB58SNzl6F/zSP95LqY/qXAkN1bMUDsD+LXDl6elREOE7YFpzdRrAmQUntTLMg0E
l4qblPIGWekYvZ9GQHVN58MCPETml+hljrNlLqF1L5Mfzh+/tM0dUs4uMde4UQl8
avdepPI80t3fxXxq04cYnsOgGnRUbI9mkhEF5iQZAH4DrWNFEsFGgbTPRrZ9mHWJ
KJcj7uIihoAJjcefa1oRkGNClFD/jY/B5DwOkfH8tPafB5ELNyBZDjdTq7iQmR0W
SjLrXlaiYQ/6f3KFpcn0e3DmbOhKB3NrHH1QtkGgEy4DUIGPpC3/ECuqBIPZYTQ9
BqRO+DLCebHXyXnCozGExwRm2vTZ1FY0iwYYtjEbZCOBqMzheZ75tYrfwhDLUPVB
+le8VmCmYMuxMtu+3ZAXgsr/GAQyFkJI0heH1e/tq6zGXPrymLgJd5g15mar3cNo
rWNifHlFtl3WgoGQzysiec4DGh5qBsD+apE/Yhj+jdnQyT/Y8fXNNYrEgOGZOo7s
L7RpbVVE/bC9dzqHYZUuCgfeQELmVXg6Xlg9OxeyrgQ9MiBFgPtNGnMrgCn/lRv7
fIs6RLv82DSaRrhVQ+uZkJN1+sBBDFzxiaM+WOkRaRyR8a4xfjZqS+ZWQXC9KA2h
FLLRiCIl84q1DqfNU5WcSDYbA7XNNr+wkRGqk7ZUd7OCoB+MQSm1+9Kxusf9aUQI
+l0w+VEo5lg0hI6ayWrzzdpYDb2W0Oc7c9t8vBd+6OQdRoXRYngLq7PiOPjSS19W
ntSZODZL9Q98Qu+JDcNhv9Lj7Qu+Lma6AHX6D7S3KB6muTPoqVAkcH8XJavVrLg5
W7GRTx5C2USEqxNxgu1nEakW7yyHhrnqYPUBxnLGBLZHzw5cqpnBhP4DErwqafxq
9EyYhtyAu1zCaBjy8f3uonHVulJ7XTmINQ7RnB2e84bT8pVrYiZbEy91zzNkW2Um
u9mOnJq1Ibd5G1At570/lSRyLrqSXuOhOmb0sppM6O9/mHJVRyd6GvFuPc1Nn6MU
D2+Wv0INZ2pN8DMH7Xpsz3fJwM6Z1wUpV/p+EUKQ9LndOUcgD/iX0Q6L6E2qLFjJ
l8X5qZEy8kkeP6PsPz1Mjps+y+SBmsGBMnWQIFM3Qi8JocR6Eoy/Q4giAcirw478
sPUhXzO1bKVVb+y3jWRyOoE2vNJB3UjmPkEP8rq823/ntB3i/246EZFCCS1UJaFV
aUiZYp5uLMshGCWQ5Jez7iX2Wamgng9lMIVIhj8BBDzInAeGf/lCQqZFX/ZfpcPV
W3fEnsc8B9o27gK5n7s0PX5QtkcxbVoQQl5d9ily+xeh3A3XTjmw2MmVS6luYRut
nDGXZtE421uKJoYVl6wtY/CBL47hJs4hqg6NaSfnOOQSJW5rgssZhW4PnAtPzXVZ
IHcs+WLaQdTPtWqo3KqAjbBduz/CuISw9XZo/hsdS6lsnM/GTgZtn9oE5ja6bder
eXQc+mibRX6RVYa4Fd3QmgPe50qvHHP080Ju8sER7E1nvDw2f+s9wgcriyFIV+Mz
XRcsy+okWF7/j1rgUgaEa0nyjTTZRzygVqHVM49WH/gCbn6roxy4TeDX18yKM5bM
0k6wQyJiSZ4BO3F0po8LTSLLA9HpS5ss1d1r2F6EjqTxILDHSfGZz3/ZNnC2+RIu
9FEpbdDYr0UL/cnNMU8fUB742hwI8lzMVadzOk2qkyqYtxVrNSchgDSI5elGx16V
pdeKOj6s8Lzx2STisrDZ6QzAyHLjsSWwa4nglerlcSIZtFIlVdVOnLLrXbXL6uB7
DQXW0Lz/m4Bjgn6NtCONKGI5WDkPYAXMRqPAH1u0DmiijMPrKpU37KlkMLZ79vmQ
Gd2Jmd1wl8948cd3aOsNN+2lJjdEnJBXw7cil0F0WMru9w+kl4C4o8wQzG652LJP
CFon6+JA0anNkqXlisAlMAh/rFuI50XrGJ6+bQR6kzjBUH32dw0tWlXFs8QSeR6Q
pGurxJDtGXy/OGPs/HgF5vJOcsOCDkyUaQKuTOpF2SADDMp3yIhRjIZj5oAY9f88
vDZCq5RvZTz/X3Tb34diqs8sYZPf/1+xwWC+fkuWYg5MTpsTBk1/WnCrnSPTaYK+
0IhXLpjV7jK3qWyqw29sBGTQvtcCnlYlF3aPJbFW7cGfQkpotlYDVC0452ELQXwe
dVKlioWveJhPUZdjNBE8zr6XjhgYGcukrTpXd314gn/NE4ZzKlB9qACdGq/4LztY
BmP8KDY7eaoEdcO0Av6No3v7D6+szW6uxm6XtpNc0D5lOBUF04G6Gx6aej/r1br2
Q1oJ0RFzodwuMMWtJxpkkuhpCXpftFzkm/aAVu8jShwZsax5E8ej2GBgzFk4DpUq
4Th5WOOVyyWZ29H9M5MEbskQkkf7C0CB++lkjZSpjtg+N6qbwOhozSlg62jZXK0B
fH5QVnpr92e2RKdEBzupwhCVlgH2h3sA8UQqGSoPV5WEgo8VCGAOzaKr8Gj4oElp
XbIUVlyw/GRimuPgavxoECPzq5MXnIUAuiNSo4o7/JoM2EyYZROdWuD+rTS5pXD3
z/9l8HmKtUVl0Gbk3+EjOmU+L8yEpHS1Lp/M0zRrSavT4AdjzjxDEqvalqIsCIUP
nYrpfUYgC+Dau5AXoedDgYMnrkQi+csjDHDh7Om7ICoYf7x7mKsINjMcCpUl0Qur
Be/RXqSpIHmQWUk6gEXCbHABOOurbBJl7BQumjh0BtgZlpQyHOsqOY28o5Kskq0G
8e+CLjpXm9r8v8LVHzaUrYlA4pC+OqLXk3n3IXKindSCvq22J/j1+7rBUVXVyohH
5ZuNjPqN19/yjV3eCl80fJk5OcWEnCc3P6amdpFm/0Bv7npWxLYxN0ya8P4DYYRu
y5FLKc7Tv/QyEx6NKBMbcVyIPbmSxrHd9I+Xdgs+6RPnrjUnIodKscI8AvySgnZK
O49SXUbGnmHt60+yh1Pa2Ri82POUEjxqxcQ6ueHL3mDmHTaLX5jx/Q5VhkJvdLlM
DTWYCXgXVqwrkkOUt6oG+arTy2Tf/VO/Q1loGKPcCLqx5xOBoyp1nK2WCXbLGGTm
JovAHq4cQFg8yF6gVSu5stkNIc3usv+vmuBEz9VRwnURkIIGE2TMpSB5DVnnYiuR
u5Bl/Dq9v0bPJKGUk1FCIVhjVEdNBC5Kh+1Lmu0uQbKAfbtrbu+C6BDQUBPafhOq
GyHv8jucjPuZ/MxoU0b6FuA4NGnXo8N4GFUMZu4lkY4OHhEBYgVMFBDJdlnnxseO
s6paV0ol3L4SiIwSnNMNUkCefs3qTW3J//98K7CRBPGDEOALUXFiHIZWzqA4cy2T
lrsObPBCr755xNCJ+xJJnZFys21lKvnSfTbPu5FjdO/+d1a8cZqTRIiTL7954g63
RgU0OU/Phngu579uptu22dSt86qpsK3rW+cmqaOoD7ptGuSYbLGcXTbCSeOCrIMR
jSoQjtoiY2Evv8Xf1kasV8k51vC0b7ZeB/ni5LJlMTWNJrQySqUnYnWZWh34nHxt
0fKLgkdwbt189ovuaKLuComXTsmgzy1rnMLu6H6i1/xKju7SOhJOzA3/atYMaYK8
E7woeo1sXi/5f0CTa15x5EhY8pWfmX+HTAfHV2FRd8e9Z8NqYSOp7BiKa3B/NEj/
ivPmU6C80tPyqQXsHMs8NKXMFgpFmL5USB6YErXND6P8Ocq66Zr7tNcWlmcvdVvf
A5y92coo8fYjQkR0FMKjZNyacEZISAw4OZVsHVu8aOQjZRzZ+jX+xyeeJI1H7kxi
UTSEjEP5YmIAsP+nfotLIu7BsSl+p7VAxDHjKxNY6MVmh4j/ZOqwu0MKl7hONUS5
Swc+zHnIQj202rdSmG3oLtTAMUno5qpMl/vsK1XKBu6J+mN6XbbhSNx9rV+Sd5JK
S14mxYNNM1ISL2RAHYOHcajXPOTVtGCLT7PozUQoI01RoIlJlugC28A3TkGlRTVE
THGgrbH+Mzd8prPsVTX7xEmdQiZwyL/2SIQEJigDZdrIFHLulUeI74sn9lSvTLMT
lMCT08FN8UgnMXDZ3ZNDwYhgrV3QPZtMVUx5Jp0YncLtBWjzwNkFc4zDgy+/1gSc
IycdIywPfuvFdnQ7iz4Am4HmainbVX6vcMs4S/xu+APNfDfhe4ioUsN594KNLp7I
C/lpMZ/j8wHH+oArubICGMC3K9k2wW5DX8rWkYjh3TC7dWZ7Hhfi+Q7ENeS4ntcH
27rdyUhqOo88aXDK+SZcese1zweSZrn4P+/K8wpE0mOdU6gq/83NPHS7+zkkr+Nq
US/xlxyNQfHql8DX5iq/ojIwK5RvgmIcRXaveN2Pc/BlqEeI1l5Dv2k0NmyoOUh0
XERqs7OG068IIfhLItsnJrnwHOMljjr5ZogcpBVKINLCJeqE2EsZYOizJANnvL9B
V+t6joZF0xOrAKzIqz6EBzn6s0sQnASV0G249x3k9D9VxwIVIOF+O8ZZ2A2U3rjl
DTo+5o63SYyWk1uqwSAY1z0hoRQKTTtSD6vinuKx9vd9N9Hc+djkb2QIsg6CB9Xm
+2zGingtsLdBQ3o3JKHgQvmMmrg4gApK0Qd7l+3i/kOPxiEPE8+ZSftq2U/QA7pR
Q4uFObZDvtZvGFDcsUOziNQpXsAimjLAcSzisJPf65v2CEv9ZRXDq/46WsRksGuS
hfQ+Kwstiny+9QjqckPI+DCN1QuhI1NSTLLinDe6sG90LJdO9KLWNKwI9cnLW3sl
OtstBbVf7XqlrRIiyk7X1dmdAybXNGrlQtnmdG193KtC9aEZ+UqgiSUu9/yyEd2E
Y43Gj67SzJSc9DxCybIK9Wc9ucNgiLIEpXTbKVnltqjOqBcHnVUXaNihYdVLNbbL
WnsC09kLQvA6VCBq+bPktOOEssbX5UqF4b+H4ksKCWATpVWUcefrvYzy4RuUAHdM
MlrxA+06/cISvPHHKE6afLBXsBmI9UMR0d85QQTKnKy6+5ReVU/qgyy6IuErQY6K
qrk4AoyoBdCPTeskxEpyPi0DwpBB74Vci98dffQAyRlRJPTTVOh9EILlJgfqKzsC
Z1ROIlYBPdnL8Rktqh8m/m0IX/KfqY3Y0dWD46hsC7rgOCfiJsjpJOT/eSFQne3l
OEwH3lJSC0MzXJP/tTQWb3FkM31rhxiqcDJmIM9WVoJq/jfdlmf+yhCX+BIfdbWo
HYtexaboLXsj9X8hIR/j60wfQRovILpMS5AicZb9mrsTwSjtDlBAYQrgUGRqz3Q6
lIDXn7EF0Q7AgN++WflSixBRAQPVZEkTQ5fygoICFzOov/qkARqX1Cnz7YDf4sV3
vAS0HFU7Om6iTb0SI5xyOFtnfJd79FkGRwb8wB4gAAcXG5YCBO/G15TJcasS2KS2
xz5P+/12YsJ/9UC+SUuRh1Wdlzhek3vTFx/l1RHXdem+Kyqvr4zGO6Irz70yGyju
h7BaNEVpm2wJDUnyFOh+fjBRxavmmw7Sxy98HAviA1JPGtH01SsVnVtlkhW7ejOX
YP+Enl1FgYBpaCBaSCzbpAFuBKSQKF8cMD7FmS1pOp+lT549W/CuHbgl9YUhDMNh
uPCnj9QMDvlgShjGaSJObdMv0HOKrD8/8gl6QZGhN78oCgS6hsNOyM5QLSjO23Hi
wk1jlSZfKc6Nwd2ZFpY8ueuMDyCpaD4cIfl2SlCoX7R+4sCcyV307udtNJjWR9aV
d5J/Kz5Ihod7Lj4rYve39N7k19lgaCZCiPdxKUJXZ3sH0x73+1XLLEsMSCeWK4YD
IbaAvO7uT7KUfQgbB22KpZJjdDW8zxU4o4PB5wAlquI8ESjKI0xfLqd1vB2s3OZ/
5c1p5y1YxCkGl7Hgk82yOufU23dRLPnsHgRfrda96gp1AH5V1gGkGGrzBze0HZBb
Lq79qhuen+P29QsQG4MijoXD0rFKAbZqAuf1y5B66Y6ho6NsJR5rQFcaspdHCmAf
JL3GcYYk0tkeubC530xHsilRBB6BOvCaq4l5ioNWvBH9fG9g/PoqNf0xrFxeNKcl
/9WFpWTVzCwxQ9Fxv+DdTeyphU53tyvatpgQTdUZYl0XBLP7+/mShoF9qwV4QlFe
e//kaa1Z6Rutk422pHQWyD3lhCEe9pLoso+eLqO9z8GtocqumSY5Dw4MwduBpFV0
NkyddbXNQFRIZUPCn2RzPpmdGt276nFKX5KHdn7gw7/GSwGJFcjy/HmTYKDoZijT
CnuSbdI0r4G/Smwcw/c1DFu77sS9b/By1D+7MiRGZAxtWO4wwdqAmP40PedcZ0pw
trdYkDqOJ02/5ePGBYgDvk+OeFXQhGdMTK+5jWOvfubUPhQh2Ly4kf+A59FufbfE
mMyGE/YfFf63Tl3yUDqEL4c3/NtuJ9OH0iGl97fvdjJJ0SgvuUoi746uXAtU2je7
0lVzCcMqI8YmyvCePk3/wnqRI8jsHNnfYTK8uKzVdtl9dvGu0/eFnrjdbqP4UKGX
evssCtAJI8VSEuXCw0RD5KIz3cwx0mFJ2h+G7JmCwSouy3PKpuCsz/B9MmESArPv
f4/VHnz+i3D7ySI1dcEGtqE/hQswfCSvLUt/2RECd7/ZhtFjwccX5dHuyZqFkX+h
m9ohTYUbMstn2d5UoCyGLYAhc0QnsRq9zCVBy/zTg9u1jNhEyyDWgZfvG0L8yI2A
z+icpGGEXfij5HL9etMNkoOzf50rk08MtdNgxzIy6sweMopqP93jfQB4Na40BEPI
nNSENXbfYCuZoyteh0Ludbs7oTZiAIaHMJ+OpBjW4C+H9ez2ayF7/XPCP98sHvlA
/W3tMXVElsbLhuKnsWPUXZUkHrR5JDEzhBR7TVbg604xxlR4i78oOlAEgB5vqGQH
8O6az0zIzjw6B4RfSXPMRW0vWnBPF+TmfL9N6HQXWlaVJr4Avp/s4N5W5ggoKrL4
jyxxeLTwxDPPECmESmhOSVSev3mOgP0UrAuqnhVC95Xex9DGVQuEBMkSoLLqtVwp
X/k2PKoQvPeEyuRHRukJ75ZHsZS1/Ddg1X4Z0gN60zXgwnl+O8lje6RVCql+1BjJ
VoE4uYrc62N9qHGGmVulTwRRmBecsy5Tpilv2aBFTr5iD84/vccmhEI2qp3dVdrk
XnASlI1/o5uqoNNr3F8nTlrVcduwNW/92Ch4uhCGnYJyhOv47MuLyEAFLyR/5typ
fNStStrenZ4n8VzmhwpUy6va6aAog2JF4tfJiqbCcndXzzn19VWgIOKmL2cqUDuc
nUDpivY09S7HkcFlSQWU2/UwiLFlKBCe0kUx/Z9ubKx3rkbgQvPXm85Ei8hzvkFA
H+632ykdBFAcK4RefWpa9NCbeYTeFhU59PbYXCAZetFebLV47SYUAwgOBhP3ngiW
8+X1ds9GUJ85wkWfVIXnRmv7wE4xLU1QBMp4l4crkGe3MvTsZi5Ue/k96LZnsBok
Ff3JcgfznTBdYJEaBoNyFpCAQ3GPx2sYI/OQGMUXbYtcafxI0Y3GMnnIWY+c3b15
8TnkyGxVbh7oYJjfy5+Wz1AF4/xvyoIyjhBA8ltGv7PY2raA/+lPgfebXUvDHqDQ
0xjJrkBXBf4iMvjNUjbld2PwFnmLDJ6fZglvYzoAyQgYMZtxzJKFHxHcGPesJgI8
8PizgXvr1A3iFJhW8KwWHjbxY3rBVc2BDL7AooXWOLHF8dp5uSKbSXCOAUPXLms5
+WxyZf1LKi6CNCEnXj7yyEy1oxmxIuin1OK2v3W4GWhrKwVdlE7B0/Z59oKrFBlW
MPF6rnt/z44aoFh11kx5/xcwW8tr3NrkwKGsO+4487ZBXvzlbYXaJKegaEuUlf+c
EDAb/gThlHFKXFMSRVVONbBPSJSMXYdUL9sW9F5In9lE4KG1us3WqJnyvRyv4DAa
0e2/xeEwdRSCt8IVzD9tinfO17KI0rnURP5xn4wuEuVwcbYiyZ4cm72UnQLCWJHH
htVihpXJjHFsHwq6o3uLMd+53wVOSV6VTlb+I5SJXlTnh4askd7UtkQWwN4M1tXX
nvvMgy7oOc9MPSU69ClpZlKtpYWQraRFsszlf3jqPUIpVqFB8JBNsSJBlYOwHz8T
pRbFFupWOS03Bz0jMGiE2bsZ7jMDNyWwbPikExg1dz3SYXTMk33D7j+Fc6WPOfoq
dPpx8uttFEpPv41zAjXqbbpo6/Ta0fVOQSuMuP+Gfae9RHIJdGHt9H3bu10rReQp
J9VfgeSQzR9/mhZvQhHSr43YCmcGlgy8QW/bcUYmpWMNPRJwBUhWwaSHlVNzDHMu
PNBviO7s3VQL9CAIKhwVjQgbfBMO4SI3frSAShdK90dFJpWDUfNLuqy9FXXanVqr
nk7AGuOpJWiba5WVQk/qhknfrOhswifQZxsdSLGWNtNSSwX12n7wU4BxFBya2Fkw
BouO3pe5IV7+Ep4calaqNO+SoWgWL/kJLKk4SEIugEpwlk+uZiKbRPo+UNYtOLlX
V3KUYcQENl8KO1gtNEU+QLNqD7euNJEW7PWAUCKtWB3h7HN9/QOJnzH9qKoOUVL1
2aqNuKCnQadbPpmiteW6iZRdqknPQsMd8kNKsWnouwgZng3y0dI/9AEzuBBHssQ4
FD6sfzAc1GraUagfvrXOidjUlFiNtyU1tW9xHZvofTifmfHt4ypVHgYxmYZaLduT
CLimBJcpOxjkTUT4c8jsxN0ol2dnJfcCpggOSvfop6SUl2dYRCMPOJjpzKo41Y+s
HX98x2UmAZlA4CnHhzfA9IbHyTJs7OzHzAvZVh4D83lNRBGseKU5KBds0WutLFsg
3XauVA3VSf718fR3RMjEtxPuhmHJ3ebYAiAGBpjRfcXcqNCiYiEbh18TqEqGamwo
hwIr7KlRAjdWShdc/t602bAPKWpGPYw3ghGSfK+yzVUG6mLsZ3iwjkXUtoxZOEzz
eKW+ufAi+3hSAh411pV/GPXdb6XJi6Nq4KsP1vLb0mE2yylB73Wfalnrn+xK/6yp
2ftYuQ36wyjo5DpoA7xWn9GdLtJWccXFH4DLVHrs4pN4QmmSjKpOivuar9U3YoyD
pNxx/UHyUFI1dOIC0f5oC6vSnG+2NHIV0bKkPjp3Ncw8G423lsSGRW8ovQbZZkzV
LPrhZmnfWP9JTaI+3+/4yX9LCWp6ofvhLIAXBZDL3PN7rb+qtjTrJfjCR815Zkah
6Jk1pXVMCVmJGWj89JasDV0NinG3JU2Sj49Tq0FtiyKMKSyYFgTt6dQfgGif9icZ
wK+rbh5ETEkr8CBf7a3x6jMttSmNkJvwfhzWwOw+KVKQHH6/TYzOt2BlF2BYgwuc
Ikf4Z1Cg742aLYDFgfcLkwnhyKNIylHllVP8CUOSDNVV+vC/Z7xPiU3JohZsFb6O
8tBUsfmlLCwZ5Z7X1B4Tv9To35jW1dE3BSfSrpw3bZM394+TjOF8Bt0kFIwWLpVK
Quwk/SAOsJPNgqcMtpe86c9aX6/Kd7P+evCPI/MuQ7Qr0nHcNT3qyR5XYM9zVcyu
2L0ojeNh3ms9n06xnC67LqRJdg2IS0L+kInuvm67G5xslTH5DT9IBKh0Cw/WFrwX
odqXIzUpbRCIF5iApl1z6MuCebJykxS/Y4Mxg9JItxlEZJeMUYmzjToKvfCmHdLf
BuunVgN37cBk+AzKZrTCkBLq60jH4GihXz/olZrAv1T7BB2AiJGfeONNvGXe/mlH
Gs4LtGOenGOfZN27rc8H7CXxYvQkj/tg4IZWNeM8OPzZB7nVdSNiQu9oL2dIu3B0
ww8jCt4GnjkgQ5ojTi0Q53iNdcz9uY/Siu4ncT8syCqpDIeRmuVjO7qZorLbQ+6e
OeL5oMw/A9xZorUF4Q2UL6laT0jPtAJq3K+6S0yCFqqgk82idrUt9fMRi4we6oj3
xSVbMnL8wWudePhQII2C7QSjGfyLSFoKza3v24Fvs8Zlr7PBRdlwqX6jwiaWChdh
d7rpsWWIfTn7CWhNTn1DemBSwt7hhBr23e46x//D+J+P4JCCAw2/eWMag7T6rcQN
+gKMDbCkIZwnMSTtsHzCOVu1bLB2PdTRmEFcgB9VNdf4NE9es5e+AmJ/IY+UatTR
V3ieeF8fwQWUx74jHWidP/CCH9yjGQU0u3B6flRqYTqczFuUUc0WiTA+Z5VgxGmG
qbESM65FfQJO94tYu6Yf5D+I+z82PKoS6Ej0hhh54jnxeS0cNimmadeL4Gahdo31
si76ks6LDXTqh3oW5mvQstUcnSUstzX3NxAzgXouKIjFieRkqn2q0IMDvv5QmAcu
iCD3O4FNNQpU5D5ZNwd+7PDTsnYYVsVmInTC1OPTOw6R8LDqC5zUAZy+DjjC364s
2OmzVkLPbtmq+Du/Gfq27d6pK2NT24rtGr6GhQ/djd1aJDwi66goLTRttilcnFdh
/qefZREU8Ik3GaIMxkbVNraJ3pRZKayPjfTsCbkt5LcRGD9d/si/7hcaOcE5gjvj
SiWEDMaJ2LIXn7gaX6nGTC/lFOzkfX7ubNKaolPfsQGvewRNp0PfJKaVtqkqKB+T
xgEsmKIjlGHEWtoIDirqdYvlocYXl+kuZYm+opLUlfP5GNYs8C6tIxWOdq2JOrJo
RDKgUMlRKW7HhoeZvWNvWSlA5r9yu5Q+ofCP9A2wz41kS+sNGUUgla1DJefrCEmi
73OcXxIMgfIf40f3+D8xhxG+sSDNBTlXNIPzhVdbx5B1WknbRbQwAyJ6nyoL6/w0
8Efi0dJbQ072a9VXcM0aEHEche5d/7kM6JDksYSBmRWJE75wHVGsDLomBmnAqqEp
sHpn2tF+KEgVqBSh6rEiSCcCggcf8DoPejwgV/6MncDW+reuHpWCppd7bFKesHTH
Gsl5z/zqTTqaHvsGIdR6skyRZ7kufOH/jjCFKGZxZc98JRfPPa//iBVNZLgY+aFV
JQVjqzQ3BTHcmfLXtBb6iar9n2Ju7fgFKIlugWrJ8FTXwYBnok2+zo63CIwTmaZJ
A4S0PPyCTKaQ/pVexB/+qls1KAnKD+DgxDUDLWR1xxVPvaJ+8g5eblp20f+EFLkC
2IprSbd2jMdXssBh4VlT0kkBQGXBO5QXaxey7IGM1/r60TJBVCNkuUcixDtnUObC
iXeJVJ0SfdW54R1QbPyHHXdkTR1nIOhR8tEJ5sSww5r4CgS/NRD3v4O4CY+P/5VE
bBbK5indNOKxK9xyadQa5eghInORZgAXyKfx9HOH3DohmqP8v6UHACpZULaVuF/9
JJ5KHG6qY2hkZ4eSXgDicoa8nq7xL8CdZ9lxHc6nxJ7eAcurpYlUR9iEyWm1+gif
gvFdOfGm/8xm+tzEF+KziIjl5sPDR/gjXwgg1huFcCQzh8hxc4dKW/0slqg00BO0
GRaQh3Z5MhrLG0LclJ3gQwEQDBBJg7PW6rWFPkFFBK47mxTfQEjlxs5d/bcy0ozA
j82t+JRoOhbT/kMCrxETOXNsuY66sPlcIkaqbx613n+nfZHCusQhlRF5gUNUcqSS
lmyz1RuDQJix2OBYg43BymSDtJ2igSnUEuCOy7LSwprftAMcGDEFICToUCys9b1b
NeVedSGwODx63671MY0qTjEsbcvsvVobi2opBRTFOFc4iu9gc+QQcgWp7F4Mu+jS
ABo8IxUUxrAPbuw2NZO9duxrrOtaUk32toyXf6dPBd+cWcERBL5ZxexMJi+LgqXN
UDVvdteN+Lc4UsJCOkVeSPzAzxy2wkasobDPsPb2+GgbDopRb8zBPwno69DjDIgT
1tE5fz0JDj4zWv2YEhTa0m9sOAAeCFsTGkj3dHjMFN8mL75kcGMbA8olt6GNwHOZ
zvbnGfvjpa8vO9NC3fEHPU8MZHZOemCjaQAYF3IyA501D9+klm95MKN0BLiN8/Fz
GfJkJeRr2smOQ4OFO42bm5cofQldXyDGhqavHMIjoOI493fFFR7ieL8OP4rs/WG/
O8UcImdIp2B8w4eIMyRn7MDA9MmvvtSFe7b7t+M/D44wm42DbTY0V+THcWG4Bzzr
pFxbZfVk0TwY1rPvt3asFTArwoi2WPQ5A5sL2Fx02IbR2SHJlahv9g3TremrNYUP
MNVsu6zuZoOGa0lrTn2g4dJ6/KDYlPm+hSht7DiXO8n83Mkk7vOr06tFlShQZ0TX
mrymf4G9Va/2DXwsmJWpnFp10EQzLgZjP477DWBQ1Nw3vcibGO9jobTB/l9pWf8R
NCRK1BE7neBdl8Q5UncVTD3sz5Rt+svRIhUiDFiRUZGTG/xs14YegdXhw5JLhscj
zLpNKtAAbD3cJJC3FBl4p8ec7+bfSC2WomrrLOBzrNIeFaQl7A0SlFhtEy9+MN8G
xzmnNloOzMWgUY5p0MUoTI8zN82BnlQ35UA3+rMQw7CTNONO4EFYBSQLP+a4sOVV
gX+4ibkBN3uwteiOJoXpWXHgvzEfw8KUnWX/S4PETjnAm6+BwU71I6bfZmUNY+6I
Ni/jRNMEdcGf2KSLz+hvqYxBFW1LbXAs8K8KVVAOIT82d113zix5NIUdN68uH00u
ED22NApezPlMX7ecWPf6nB28GOoZ/5aarnD69lGhvCTEkLdoXyJMV9teGCl3O0uW
usJQzURXZc8fNMWeKDiX48aXBs3avhYlrn+4rdrMeFjkNG7K9BciDkALeO3oqbY7
MXC0MN+4CFNODkVQM616Esnrb4sClSCLN6mOLXgUNOze/QisW6I7uasUkfIHiVvj
1Lqqu/m6S22KvyDdmBZXRL5FTNwprdYteGV+AmZuv0pmZwG6uxlaOV0nXSlS+UNn
xr++jUesQNghT+1h9TX8e5a8F/Lj8cnG4TUh3eAwozZRL8BRLgOig7wqshWD+7tF
aZiQTmW4uwuInQHVCeIOUSFZh+vpETY6aHk8lPCfycXWTPlU7OPwSafRK4YtsQXj
dvsmn8DoFKXQuEusP8Nq3c+7tuh3dTz+7CFxPTG2E2u/99ANex5qB+BznWOhUbCb
8w1LMBC8FIyOZiTmom0F8riz5WSc4n8ZExCysewrV3hRcSgMBnyAwUWK3uyI/Ntr
cq5RqAlG4nqE68Ld4FflUT99UkDjSCJ+LUQCTpqLti8C1sWcETUQkyXXOvAEZhf0
tpCvK16Vnu/m1FRfcrxJz5dJJrcTTixNLDfuYwKp32ehOLhtoBRi4gJekIsN0I6X
ULZGe84yqEgv2A3ZoKwg2uRKd56i7b9dLi0xQMXOns2rwaUSqo7fk9MVFkX4kuk6
zSeFykQYuO9Wnwd19i2uEuKYZ5g7oMITCkOmkk5BqiPB9OgEJsHDZtre0LLTbDvM
wXTFLoKc5HXYQodQVtHs+ZFecEgmnrFowjD314qPuSmK1pzWrDTuSq4OMyZGcDWd
jkrYd3haCZIl2xcSqmlDrVfoF8qIA7J2j9GNNlxOIRGFmRLLtG/UmKqwTzvHLJyw
gqMd4mFONH7lcJeh3rPPkD7/nlHfqq1V505YfvqdrEcLYTwXyPtpYAdUPu0RA53O
3iiWyH+I4oC3UZ3eeY5xzkgIoA6j/ctfkURIgRRXY3fJ4lf+iCrsPCCqNiARVeJ2
CJMxwHMvCL/MZm5usUoJiuOxrIqJ1p5T7ifvAQH3YjpJIYjRs/JbMYnFuGGMXSKf
YK37pU6l6uDuPs0gxIYaM7V5abwBAv+PVux4GikXdSBxzV2TYN108AX6qOeMRgeq
eU5C2f/U49Lt69fipRyiuDbART/mvkV0qSPweetBTvSl6ZVSqjZp5m8e9d1I6sxG
RfmPXdQOf9SVUm8NUS4BjLWqY9wGEapD1Kje1/KEwsUDcv4Qq3vi7NPgFH3ygA9S
xMGofx3tLnNmAg5+hucXfgrXBLPtKGM//31DCgAYL4aTg+Gfr0QRCH9KGvF3OqXy
vHtD8/6rN6jqmBFNdAj+qHooJ2oM0Pi1WXuifygyTbL6RiVTwHx+auTM8mNseOAn
+a0tfLH3Ec0gWUQgxn6MTq9x2Tqm+3uH0vPINo5ekkGxHEe0ayyKQsOSNh5D+TeF
6MRbgqGpky04RifPqFSQwrH6MWKPh8wrpqb1pCPyjd0V77fS69GCnuA10eBZOzjH
eoYOEln5Ke/6Eqs/bt6/GY7Ql+6ednc3geVFWAFrOmIZnNxHsC1ymcWjicg6Malc
4lWTUdvnzjM3aohoDVmPYLheUsY2xgCXxEOzqFkoGOwB7TP7VqMV49grVxaza1yx
Dx5Uc+jy/vnWeB78VGdzLxnhqGhIZSN0CrOOSgrOMMEEx7f2QCLN2ion58ggez5c
jY7hf0Lpxz2C0CjOj02F1crMSY4FHB7S6GrqfBKEbcXQSX3Q0S7LykbslcfQfVRZ
/RXfIt+30UFpFGmRUq0+c6KkZLFR5Wt1p1zWbQxcUIPRpGjVc4lH0mwzxlo37nTd
VbCdw3yktzEPgrtqXOOkFlSqdwTHoGGnZwlplEzPdkpVrc1MAuWlUQS4Zr6DXvKu
ghaUVCTksnhJjU1gpzRqMTaY+7Dn6HATS9di+Hu04ZAa6EzeK7I3/d+fK+FT/biV
PlK1f6aVc1jEMajP7m1lHs8kxOJAmOCKAGVVVM34SepQPDjQZwwLBX/fRyiOOj/L
52e7v/jQUWUy19d2GXm1BJxbHtN4bDvirtlq60RHOhh2LcHIl+X/1lapZaEIdICB
FhGbEdzXhNeISyUl98btTo2aQUQD6P4ojPm1cyqOLbp6aSr0lYTC4pjoEmqizp7H
YhvkY/xlXhc4SBB5a6i6a1CZe8PFU3+TRLWOTIcCi6ypCMegT/wXeruejMN1Tl6g
7TKzupG2zyAFFYgISzZ4UOD+bxtQGHjHSz2gXmnO6Uxb5xcD8QWNLOd/ivsUv5zv
R+2wTDSjeaSEEUpwhb7yQPQhYAFmiVi9g4+w0dJFp1oGdFEHjiPKQLX/X4kfZEmh
ZxjvN7GCE7TUPfOpmOcymLOwAJw/ppqq4GhdIW0eoddzKUjOKTHOOOiEIeN0cf0X
BlaBNE4SWJDnXyeRSmHtQa6nhpVPH98tI+FtIVrR5F3pX3zexshsMjt4RG6x76xm
06fIjehrteNVIMpvHGFhHLl+OXeP1uUldFG9QQrMzUXtZ8m9GQcBnD0SY9/nPGa+
c5oX9Uftm4xu2tCO0e16z5TQkrkBGYx03NVi6/Shu3bbr0Lu86z3a1y7tPm5W/Kb
kIv/UFUn6P2N3WkidkVB4R6u1bB5J/jYx2XTe1amU+liasOA4E7UgYaeuWOalbgf
0ABnS4qwMokTfgn7jex/SzucBK0JZkrZw4UQoSdwTET0xsHge3DT64fsaa3Nkwb0
INZuKqtvfxcymodhtyLI0xmOMC9OmyogIw++8pp4i+HJ74jGG+hsVTEv2u+BZmtY
hcVjt+bHOAedR0iI2tC5JBozgsm3wE4Jc6eh5nHbovlKBRm4eiFDD0RWtcitjvkS
IwD5KT8CV/FoPIav25DK8v1NLtG5fits4YJfzBnHxfCA3T6tiPoVUp7ASUDeqCoA
PqaQLQSqRw9e4sgHtxl+3GZYr7BQ+O1jhhm7nurcdyd/GoBF2CB9OLcF7mzqeGFF
YgDxViJ5uuu9VcfV4AFgS9Kb8uTrvppVl2n5sq7DS/YKWHf80UsFP07oSgvDKk1N
AeHMOg1bo0EyLN95XKxPX7FBDnGKk/sLirCsDAXqsZXQ7bassLr09Edl3q+ba48Z
ao1EP3cleydqyqpPsTym5ynwG8aEjy+GfNoWntFkpBTPaUbyNxVsEUSxB9my+PFK
sgqpsL/dqcms33ZxRGpSSD/5w7uRX3Rth6785PgfKko7pYS58db9ihxJvKgOBjpl
y2QcXqdxkkeVOkj6KbeVRfnzqTdZlEJkfRJKimSdU4AjwogN5RElc4nalbw4BCqN
mwY+Blh2VMI6YxfX2raj1yOtPjmN1FG7tmDtyA54zQcM9LlPiwvmlROECDmaY+84
bcEj2Qrh2lJi48BovKzA/qTf6AregkrOsgwWmXW5zeOW56tFweBUyPdpkQmx+hAh
y1KMyGNOQF/b4TDBrFM1UzvqA7Ku2O07620vhdTj/lNxFy/VkU69dhpp+Tv3nIKz
/Eqh6yRxW1aN6CUL8Ku94Ql1nFlCpseXWGrUiEplqafQbLAvce2c2LDHk777/FH/
0yy0+E+ejwECLnRK2deCKCGTF+LE8s/ilGVrZzPUS1KG0IaL+nEubUy8TpJNfHYw
dN5XI+KuYb7DMk4bXzoCaIX2JOuRo3/47MwOC2lzIMVDTjzlx6dqugK23xYlesd8
hRrKrG3+gzjFVM+59XPTB4VMyZP8d4aRTKnTFZWLy/n4wFkptaJh4xZF26/ZPQkr
AeFTX33QqUawhE0wVJ5ffBESb6MHF+cvT5NFGw1zURtX+r5Row/gkafJcy9lIbba
LM4MVs1OwW+ZPcUvoEOppJz/+PDDRumf2LtjuSL2AtC58X4F1NbEARFxYEwW9FIc
ZwzXQS2qH2prOqByx1ImwdgASiMAIY0sKNrJoqkVmUkWUyVgVR/9rx9XFpOF42NI
r13K2tkCf3ElWG7wZfbksaAZ8hj7ZW2j1Suuw3nt6+haz7GrgrXddKF/zXU8Fm8j
QchKGtmYZ1gCf4K+vBcJ/vq5ZsHzR6TXzuXBJ4IbYGM/LFqTSveuVFnXApv2h+iD
vuaEoB2rXvRJw1kU7SPg3pWkJzGmU3RXxH7Q/CQnIc2XTeoXx1C7XEdvfgwpJctW
lAHx6Z2E0kejsz67yVLCfi8wqD8LxSnT0WD9HYTA4eBeJSB+qULZ1ZCLMp/PqEgy
JcbRBr+KPRH/vFnoFsagy74hRWNvwqCOOSE3uMb8RmfKqcrGGRk+oHizggyBC0lm
hKXbIKt7+vUxY+iDxMuVnTtieVf69jqCuB1I+5GO2z0MZmOGl6MAZaH9z/WUGClF
zhvmBegUgFdMCN/J5KOpgzQqm4Yl1sHL55uFiYy7z25Qd8z8tDQMkpSJq+oGDxlv
N/K6niHe5R9OF8UpI+DxKzSUXuM5yDd/1hj5l3rfKBIevcQyJ0yIupEBVIFv/wTS
k5RgpoV2dk7+hPJHJrtZJEzWi+YIJt09tMB6ic/73+nnRplRiaSmyN8AxRFO8tif
BreiToPUCH3pkbdQylhddb4URMlQoY6ptK1HHKj8U/ouhlmN0MLiuiFvYiJXtBkz
INQOYgW7zomsf9VHhJJUqQlWldpYspOr5bLq8X05cdqy7nV/epx91wE+cUyAU9Ql
OhDJa+8XFftQ1nxaqZziy3+FkTMw8iThBJUUD3z/OSlESo49FaEM2XwVTFNikq/r
q2OjwJ9QhYan1jCsGF4ap6vpUudP3/PpriqGXL6sbTF8zhXO2Ve9OYBtwDOsJUWQ
5G1eu9lPE53XDV648vqRSSkL2S5QBhGks8nfhkwjOw2SV7tWQnUXpwlWvSv0+6Pl
tIECXFuJfvO8N+U2JmF1i4ttCcNMkRVaC3iqtJnQrcQ8TRNqIsW43m02YRwWqCiQ
dcZ6vsqWBpm62mMM7CjL9V6ugUTx6nr6MObjQ/lpBiPDxPoIDkP5kSlIz4jYQBRm
5E1ttNmEGTwTRR6AXrLHAP8SyRL7tu+4BnfMOSeVcquJRlu+P0yTpJq43UGaV99l
J7BjE9wG4+QIQ7MhZvQQNtXlNPhU4IH9MPLqmN2bBxdHsepKLB92IvZzIvJqJBP0
Cl+lS61bWYOiYTxzAzd+tbzPFa/3THDUayABP1tKmBI9WQzvXOJnAGJRfTCaQK3p
muY7iH57h9GOYH1bZdp0iyAf/cmAQBJzA3R0UX+5sx8XtnfMdw89gMqF3JD2a18M
qQ5Ng3M6Mat03OAtSqQdWtD6rM+rscWbVE0pOdFdLGjKPi8yYhhQf3HD5yGLZwVb
qinLDjYuXUHeoz4scsaLQ4rYYnadZzPufPWpsINf+bHwxPv3zWI6NpAmDLBcodZz
xwK527bPqgbPt0N3yYTPq19sjssHYT8dyhqYMThYRbVVnQxINr1QuxfGlD+9dTvK
lm702I5anQW+WwZHX0I22hz6EFbsJdrK7wKiszIQ4KRNoi4K5f1Raxx1atpbmkyG
q8prL6UV4mzcVHsgoMFN/iB1mE/Rw8pw9x/brE7E3wWLHAINSfnS5xpNdGGDeMPw
vD2gBRMUEEi4bZQ2LWFnLB+5k+q/3XNsc996dj/8Wg13RtyoFqbPfnPyYutdnhff
UI/yO0ta8eUej8pQ4UwtUWykCqyrVFm/bjU8gyHmxp1rOHNQq47h/q7biv1icKce
LoOAxC9TXRnp3EqGUKc94mG3+J1RuzzYwEiLBcYF3o3W1a8ic5z4gTX/x7Wr3nlK
EpOobtpyzw1vvjjJaW4fHr4yt983+XBVBkwKsiwAHhZceZJExFRnb/2RGOTFLDZw
52objGXNMXAEXYc97EIa0cqR0OtkaxMXDGAGLaW/3y905rylKJsniJ5FrdeVrrq3
i78jmbP409qdDGFFu8BbyuIbJomPnWxHNYa5uJkQOfmhV+yhTmFyPWCPbyh7578u
PFwerRf7xqSMflFBgCVL9/TILa6KRkVLRpYj7GH6gf/LO/JuuGBi6eSzhHJ21hQ1
/dHayTy/ksM5qWnP9XCkTvwuumIuiud97nmXnRa5uJQWYWtphS+S9NEcvu3xvCEB
9dXPcM5iqW36gQB4b8kz0t4uLkujl0TX97BBDKuK7YeN9TBSNQcp7DIBGcDeW7Op
KK+vgh+nZycSaZ8Q5aSTT4h3WipkXu7KiifgKkvabmucrOVwtoAmFSgQQsvCW9dl
pXMIsfp634J/b3BlFWGYuiMd26E/J2TjvnfANfJPZGq0W9+vGJexqkTAmnoEkP/Q
zVoX2MFK2lLws+y1Lm7JTEcFi6kY8wO4KQiGVGG5iEt+4//DHj4agmQtmDaJLPFf
4BqHP2dyh3Gkp+6Lb2HkCi+5wFLi3Da//WtN8a1pf4JMV1DA4/GVA7nkiN0cOIca
gRHotu6F6RXL8Cwq5TNjx0AMD4hqS79BTmFYpW7iHS6n6ipXdt/4KG0FzmZTq70m
azru9RrcKVdJ4EOdqC6fSPCD+1KJS+9RNYLeTL8gpwB7OVXgX12O/XdmE6jk5ewx
N6xzquzMqf5IAl7PByqDjVlI+h1QTAVHf1+qcN0Bv93TpXr5l+CGzNDNyN9g3XSM
dDR+iN2IbaDsANz+SDS1BJS6O5hCtslSXl0tXBKdGxpXutMF9rURS/haPdALE+YB
DrVCXTkltQliO/Mtv0K5H8Y6FIoH2CCaLC6fV8L4aJ2MQbASwL83mZG1DKasFdDJ
Y96q6GyIqV+xjmMXUaJYXSaOpMIO84pIZVvUQrgwIxvAuDZuLSPnaD9wWg3cL/8a
L527wk2LymaWueIvUzGnzX9LoSWRe0C9ZIPgvvsz7n6u3GkfniogeIv25M8dmXbT
7Ey8afE/md9t0dvYibJCzeF6STauiuBfeFIQjyy32uiOfFnD/5/CnWXSlqgydPR9
+4G/68dVB6g6gAezsHiwNtGOMWFMe1iKPDLXDc/VXkBenu7S/ebm4Zcz55D2Xt1W
b0s4xRfVjtm1QHYRxYUE2/XbA2SBrlLsbDBWECISMjkk+M8qbi0AfvkaWJA6TF4c
Lj8wCuElN8NF8e7AXyCInQd3dNllNC/1wYYFdl9u/oC7Ix4WjFg6DukCsGuWVpi/
z17KEKiI6nWO2sR5eJ3irHwdA3VjUD7a+k4GP8cIxugXUpuFRHBgHHhwKzyBUimG
2nIQcztuq3WL++SIHALccAWee7D3wY/1DzCtyrgLi1XKdfgCUr78i2qD9rVOGml5
jfKCqdCowiTAYkIOfK8s+7nbUyUtUw73mr6YjhXHuYFxGuMpSGUahCPqo37znVMF
37ikC+SHCKy9jfoaGIXfw+u9IV0i3Xbs3+q3nKUvSCCaWFIyMW4y4VYdq7Bh0T6r
UaJcT8FFcADakZo3Zm2uuftLS+j4sHaoZAwyVzV4PAusGlJPNULBjJeR9EihWHVM
lTecrGdcYkd781DDZnv8sx2XGxz5F1Spvg7EPa615XCrTFGYsKo7K0ajidQQY+qH
RE6hehbMsaaE/HzKy2rA+3Wczticpydg7budwTazFhQDqsQFq1vTH47yY4o9IFlt
w2JmugGiZD6jx3FIdkimK5QUWlwjtLZOXhoyAHSaOM2HM2+vFjhWQCJuHH0u54Lk
OfjikWszRI/5e/NDcwW7pd/n8MNIYs0tl/874AoRB9RIdugqU3MQSFjT2bWp7eD0
AQ1nh8oirKVirpnM6YbszpRQZvmUOyQAWerjyFmbIl2T/jjo1Vo7Di0FeeaP8OcG
w1PBgiUql3pDdoCnix4bnJ99MNW1Nd5ndAk/0kWZkdUn/EyGuhocJ/PTkzdwIyEd
ul/px9RsmsSPfragTiGMBWz2zvDxyojSEtnj5m8AobnwgT7rzJECzW/aZvrW59sZ
BgME/b2s9XuVopaRktquTbXqJ6lciIwRgd3934xvsOqUcwt8uECxyD69+lj+UNVo
9fQ0n5w34WAiZ2cBQk2thGYKu57g6R7ZbixxXhaMXGci+ZCHMb0cLzUd2MBbvz9Q
CgjGel2OgMjyW4q6qju2KEIzsFLo6ONDYWMaS9GuZSGZYZP9D/aK7tSvy77a9j7X
y6H3Y5jWGY40vD44ktiZ2GI8jL/Qt+izr734d4iseAo4coRXxs6ce8J2DFK8SxqN
VerenuHJWN1yfWxa++Y5LifTJ+iPULqq5QlSKVCesk1eBsOEUqGt1oW9z6jKbPBG
Cwki+mmPyHVEpwP9o3SniBiULlozQSC4X6JYmxW7iXStmVJ0UfhNiMJXPGN3AOLP
ccUr+QBaO9gfjhHGO18Xg2JoaO2EyXpKnR3rRA2wEKZELpISZYMr0zqPtQiUtAMU
h2Jm6BPLQk129rXsCFt49Z/FEULB9XMTCxqRm7bbI7A/I8Qu6Xgkt2EJDn0rSI6I
035s4fg/loQRQi2Xl7Q1zBUXBlwbHQWuUNiCdAAxUDhK26VleVYMQMK7WgiGVzd5
Xj8royWUKr+yml9IYRbc+z+ArB4TrsfYPy0HZIFU3MVXoWwjh54uZ5pE3h5V31MN
CR/TXy3lxd10HhV1Z0Y90AveqPbve2fAR0ulQLVV2cIVYjJyZvszWcf8PwLtESP0
4J+AkKDIwo1QtcsK5ehihTHWuktHmcvGeFq8FO3RqaYu5LLOYByWdW6PeGnkV/Ca
/jLIIiBu/dgBIJhDbLVs2FkPiB4iePYxJedth/zP6SXT+vrhNVCseUbe8r5DzJPw
vfjv4KD6dSwGoQPL757wvLbcIqy0lRRq97F+QC0zcGHNIxrFxiAZBg3Pz2Yv1N8U
kIDOkxOUM/FFSrKbGMKLxUarYQFk0l0beVvb4HaIpImZo22QTo4OeVNg0zi9uEvm
rzd4Dlir7+uNCj+Jgy1HyZ7HfF56VV6mdr4wQdAk125hsxOavRBH3nzSLPp0cJzA
TbPh41Omu8KOw87i+iPI+wbiFW2F4z2iavfFdmQnkqHGUDqgtN2wpZYpQ1BemaQb
nDldxD5/O9dO6nkkUyxYMBrh/H0HH6YDRl4uBNoRg+8kmRaZF3Zq+5BHLKJFtETz
/cuSasE/ODGGoM2TlEJ3jYePOTavRZWnrFLtVgQMQ2eWWbj2l+cG3QbrIJJT4VYA
aRhbMEQ3ZdAtCxLQamOMDn+fsaz4dh2dIA9BbGnAphY3PKr5YmceSbQ8eBJLDrnd
nta0CeLSivE6jfhTAuFUd26m5i5ZJL7qavhfh2HYUMZ04qS5+mS5O7cWYbg7LEyQ
5G6kAl0K541XFhceJ7JfeTSLej2tMxeF0dZTGYBKj53ZdRrhcwtXRp7Y3po1tKen
eHqAJMMGUdjaW7lP4eFzoGa/f/W++x1rAX2eiS4BNts3Oq3lpimuZBfGA43TTMW/
jPbwJL2LJbVHxKBssdc08Q1BuMtz2Ir3ZijMCarYtTKCMz6Lsys+N1X4xIehXxEN
YgEawJWqI6n6ul3F8AYDLIbIgPXnmYvYNEoD74P11k7xy1pshS5BZzqHBxAxznjl
2AFuT/RFN0OyR4HPpU2VzWJo+ewfqtwVzq60yv4Lg12yavre0hh/EDV9ML98illA
ulswMgCdMwGMEWvnGRnxRpZkOaZ7lEHxBMUhUvgU8SX08uKfTYoAOeVoc8/f5EXb
wqUeOUFeYOVawrWQwOOTy5wt0YHRrocJqOKgrwKyo3RP3G4Lg1WiFdIBzOBT/5HO
RcRttNU/HJZeqWUA0frtDJ3zC0Ajj9+mnUelNgdTYx0WjQPbCfuQ5l1ha19o2q01
nbuyB5QORKinJRmeDadSTMMicm4O7XN+5f1rwNq4VgVYVzoDcTvcnujgD924Pcsd
uJsXBfxxUYGTOw3LNrG5yqYIZWjbElmtedi8grQejS2xLCsZ/gU3bHbc/Lh5UtUK
TQHsrgq0whzXGgqp8XPgSrT1/sfo7d5akU4GXsMVejUrWecBJrWwu+w+F5F0gLAB
fvyrZKyEIyTWhmXtsfuzgZ+g4vguBUVJxvftQ752o1U1k1Mky9fS8Ob8SjPSFRFY
rod81up/PBgAs/XNKyYwEnquyNcOfa+kGTR/s5cxVh0ADDUH0BkZhOSwCtqqZEvN
AKzw2J9sBQhLtN2DObGOHxqg3srqEjySPeCzP3Aj/yKzOa2YWrFnMu/kX/aBlPM5
TZdwLZKbVgKcuww6jJn94tMsafUGLOpbOXo48KqvxQwDaUW0OyXJvE4XX8x6wrA4
+3cTySx/wm9Mi78cZVggj7V1rxHcFFtpCEs3nHM4ji3RjsqrVfdet3ZwWDJhRMlL
CBiPHYCbRY77xFnJ6F4GQHVHHkAiUTS1FRg292k4u+7nkE4f1s7rcXoRLzTuLMnr
2rcWUFZQ3VjQMDuW1UCAaZVu/LNSnP5hY+JK870rnVQAB5Aetn5/VAuAPtyHJfYR
VrMt1yQxCIpu5fVu8xrBYNWIuwkrFpWqPWQuKLYNSGYKgaBHkVKh68hwT0+CHnXK
Hh9Tnp75hcrdtj5CoQeho6JSa193zgdanfUWkl58aRJ+FDwExQaUwqyirj7tGhnr
lBN6LUnXm2MR5PQY6/lIUpjXttDGoByMDfD1uVzi6W5sm9XCHBlXD9ak5GLY7hG/
DlHx5gfB+2bOha3hOBCMOEtSSH/q4dkie5GNbrOjdu5YtfNbZDDUoKa1YjaUPAsv
jDelN0DA5tt95eBbeoIASBfRTVR08RZJSkPJ4VK4MtlohAQjwyAAdeuzWdYDPFkq
wTWGrayxcjkxU39uCqYNAMKrlaXvBRXXmduPhXmSZ9cgueL1krk8eyQRKfKKDK1i
G4N6O3qavmkdLLmLjIKpGKJ7MzfCvylmeKmmzqA3DFjvyifezaAQY59Y/Q/WhS7B
G6CmPcBWGET0d+DtABp2t/uImgUb8+TjPTNs8qjqDwtSGQEvouNgPz9fCwj+9cu6
x/l87qe86bDTmSmLFlI3L4vXHTsSK2CbNXRW4CWH1AA51nqc6uyHo8th5/duF1MW
zv0bfguivzC6VfbGtEpJ7ZQYgjdNTxJt7esJKM4KyVgn7LVTaYsDM1i93nVel7b9
d4aKHaSSi29J9BIIvcrPhjIs46en6wjr7df0Zcd2qr8F9aOqwzUYWju1XQJihKnJ
U3p87V1L+F5pqdBwhqMtJpyABqiFcKbdpR2MJPSAUlfqpw9THQ27VSABvvGKcf9t
sSriZhpPQMUslWE2JoSDktGjZ1C9Uao2tNWhwtLQBzUCyz6mu3yeLuwNY4GS3mmZ
VfPT9n0qqOI7yHPf+AHKMSm39UHX09QbMlYRdtkt+/myass0lJ+hHul1K/Nm0++S
zpeKVzDwPOZLOTrc54eEiMn/97jr42zb6ck5c6UPGzRi/+2/+j1BKxdpq8JKGJNo
YSITN6DKGrywP7y+8RYB3HTQEHbdpw6S2hxfa2IC7O4xbg4TH2A+HYXImdGfFTEQ
AAnPY81SVLqgar7RZqbVJFAo2ykzSq7RFuMKpvwCKKE5hxQ1w4gFLFyX3O+j6ZIA
kcP9SIrmnMHB8No44dox0egZ4sB8SX5Au2PpA2WdHa5YBCBeNNspUa5OqjXF2B9i
ykQAwrn+xjCS1p2g4z4Sm0DxzsC2imZUtv5t4HHl66Tr2mO6ZDH58nEsdZrU2guf
3Dz9QfHufNwE36Em69vVGSAXKLZa8DInAx5HT1cLZF/Ry21h4cahAHnioSiJaI0V
bOMjfjPPm5v/Yiy58fBXx3kxdqP9vFSECOGGoaLY1vvjFoNPCxEDOCbK9ykY8WHR
JWOCIjxvf/nZdmQPdZsPB4LZg1ydG8fJwMc9u+c3gV+L52cE+cvnXXfhJmHn7L/o
Yk7OSauE7TLWW3SlBDZ+8RL6BSTraFi61VqRvIAeuZwahtDsUOkn0wuhyOxA7Qdj
BtrS25UZxA/43fGlUEQ6xPedPHCZwXpAPDkS8ufUzOQRLYz+CYk5KYAijr1jdfPT
QiBEqxCUdRtLGqgkxPIFwKgnzyv59o7/vruFEEUnSECbFLwK66E40BXaIIGtn52r
aI26X8JzvwmNjZUB2NSnipLWTPMzisRTt3dw3UPn8kFY0V4DRONqv6kIVtsTR149
lTVo7yqWRKw+tI8sKABe9AoVUGVt9V6r/4XjDBOw3ZZy/f9M4dru3X+EfObgKUrO
4BSvRDJ8zWoT3mjyiHBTbGizCWQ/an+K44BjLdlqUk1c+dC5kaJ6KKYn5ZvPAdl7
JfcA5+hg7iNaq1Y1EvsfIBwdVjMVMk3nIoly6ugv2ppJugvXcrDNMSLCDbfZf+tf
3XZQlgNmpRPF80Qz2cGm0eX8X0RExWp8IQIN+vyZtJzz4bpy5ciFSAeDGgA2S5UG
PyvJOwcZTsw5ZehPLuD9y/z27PsEiQzG755sg99NF2ECxHtjmxkMQ15sEHllqyCU
9KFw3okb8YGUuquc19MAjIc1B1LOHJEJHyoGefAKDbQAk/en5DTSKhCPEEAw/Ts7
To28oFeUzql1hEeiOzSWaSaFO64AODXsfpyq6FKaAE0o5hBojA61oLXMmTvRvWoQ
Wu+i0avonKZFA3As680FDNhZcDokpfUcD9Vp/AW/ITedmqAMK2JFL6Ios/6eIFwh
KLKcq4LUa6FjED94Z4cAOOHtik4uwKDw2YH+AAsCB7CidvEFqN4GgzVTR6YCZC89
1jeso8dQfZlSVicFnFaSxt6Q81cXOczB6pXgGZ0C5Zi9YG2rFv5N0puV0tMDkJqV
U4BI+h2LcctOESzgOQZqMgby78hMcV/QkYaGbMW0t4Jlq/TE2azmJcvIHw7pkRRF
C2DIdqNPENCK0E6i7D0XBh+EvE0gv+eXnYACLTfIzSZGhtEeo/ajMa+hr6g7A3Xy
f+k7LPecwy+DdYYIM7MzRn65Ts/Q1CBX9g6DbnlKkRbHBikUfsdSDAA+e/XjGpiw
D0MN9jNEwV77/rQrLCEzD+HQDEVzSbgTK3AJ30MTn3bBOg8KRDG5E7ekz16/xFfz
wxOeMGrdWUZlY+bjtAqX4h5mWG1L1yUHaFmLntVjwY7OWKOhkmoew0N2aZpVzQhf
N35Wm7ebZBSRfjdzZ6hS8B1ApVE0oxjZdXIJNfFYAU9GZpZOo/fmY9CVqXkMpgy/
s19TE4kE7SsZ0f6OXfjKlo8pJa6fSZ9C3LbzgCExGJg1J2qHC1v7KA+4hwGLAk+R
09oOY4CtJMIL/3ouJly+kM5ipWV6GtPytzffqecyJjblm1ThADaZAfeJmmhJFayJ
2EJZOBPipLH1YI3CFfghsT4K0igbigiqL4+vZTSfSJa1N/JxvjTZ1FfmE1eCBB/p
4VPuOxepiIn75llvtu14bT/Qz313lZP42g1/nl/M8mrFaSQ41IlMga7caXrZGOMX
BGP9miDBQupZgp9h7+TZsaMVFG7n/md2RI7yYqTWLGnydGcL3pc9FOBRWdOdOZgW
tA5S42VplAVsbiwqdbQh+TejNsLu/NdXoP04y1hsW0QmFA2s2SfvOBXgVlGkyEfN
O4FTgFnYzGsFz+e24OzmG9WfsOkJs40v+XFQJ+8Qh0ncHL9IhsO7TiBUiQAY+UOo
B7Kk00jtN8UxeBixPt9IZbsX9Bt0JriEu5nc23Z8J+EfB2MsLutvPoJApRL1VoUW
CbHg2+NX4S8je03SsLkpZ8M21OxHlr5rs3nSoXyDLo14sqTPpGr69ur8v8J7xvvd
9ST8zK8WN+qeMmd7S001/ckCq1fVD+3uyohXwt7OqFiRpMZauJ5bRBxZBAPH2iRI
xGDBG17jp1eN1Czzx5/1LjaMnjtoGSONnq3S8eRCAz3jk6acUUBSADCN6rFv4Z7b
NVM7uOL2pwBpN9WdOAW6Wcc7o+EYGonkMhR85WMtFqOK9LGEYcsdek4XYCwj+CEN
BNeAjr2oB/zBHTn9sMnBG6Qr74LeC7Vr1Hxcw2QzPCg3brO7ZNykEQD+kCRkVGc7
MeQNdbdaX5Zvz+Q2WmQ8/HnI2vK/9itVgmAeuMQ6ZuurqfmyyUXy/AkSRjvb0Eof
HS7Jhbcvn6m26PRgoNYGuqiulsG5B0DPykHG4IOcU/LRyf/D3v30S6zG61EU26/h
tyGdsyZTEM+rGMINcN0ZYp7zFgbBf5seZExXFTP3FogsJN5WaVByCEpuz1k8qIfO
i99lAIBikHzy32aKokK859QBbKiN4lGVdyW9bh1Za2JwzwV9cKtpjO+m+oXc2B4r
KWR+qEpF3ERCDiW3sEvByzTM9W786KZBUi8NwCHmUc35bl7a0FAmloYXKeB+vzEp
uDi0LaQzYoWDqpDAmCGmZc6AxhPLHhB83jRlEPiWo10W3l7dhm6NseoxYRDoPZdN
B7fR/ztXGlk+F0pLdrqsgvAjn/DIyBe/ehm/xmLWXNGEuPt+7GcVpRYyZ65GDSLX
lnqL5neYCFgAX97TZ+jIpMrKb9gas/VumU067GXF24PSgljvAMpoY2SYHHoYgBZh
3LJNJoCOZ0PKJGCLUfFKCWWwfeq2iZ6O66ZO+fulXRZmYqfKqR2GtAH8iitzCwyY
kn/Z8auH9LbXyk0vJfxCTUpp1mg5OE+ds/Xd0SJDDHRIGRj5zJBYgIA39IZwQC9i
yHfeDadoLk+od/wyjcwhHsGGvSfug33+alQXz/PifSznG2aCVmH/0HBll9y7Nrie
Cj7eMeghCFJQRCxHn3b37t/2OP7vZK0Eks5npPyFFsyGhX7WDdeJk9aBdduAEUL8
zEABHKmLho26FzYJcFBNwgOxSn7dy+VYU435PFEv6Tr9GaQ/C4VkXCQMvFLnXz5S
exDblc5Usw7PPwz4uiZ8vangGduHqi25YegSMBTVM+iEsZIuAvN6jSgzJetYI3xO
S1uM+r0HXYvQJOUQBtUbNC5H6Tc8WMkuuuEglj8StVy4ftmFeQwqQZdH+4fIwFNs
iTFQPj/s/D/eGY9UifDcbBcwl6W7DpR3/JufPvL/5maOLAkQ3jWX3/P93yvaBe/R
jwcTkDXu4GSRbA2p91QelTyjIjW8TgmHwaahuyJxcAgOZPNP7rnJ6GGFIckcetK0
RKw7AkaWpw6uw2BuN4R7aHlyx13xaJrynbjV06/085QgZOigdBJb0pejQTEYB6s6
VSF0pQhc72p40jgHTkCv767zYLfsaGOHeGrnIHTqm8/a7xTtQ9PBZ09pecqBHHtS
Y+zqMakUO+F2HJIK+baRB+ieEYSm1ALIAt6xGuXNqiJtGT4YOL2AHDM5HqE8CDBx
H81Bx/mqrRfR2QYGKHTlMVvkZY/64S2WsOpBj78hsNebQTJLD8LorCQFIrGbuo1d
5eoFzDZ0Xj+rGQcX+JMxDpeFJfdbVRJN85VHzdWuLh3fv7NJEe+dPa5lAoGp0jce
fT88xSTFbESeib88jIkQ00UJTweSm8JhwvYorZPbjYJIBTKedNSdFpBSEbCJkNeU
hsONUNWu72pLEFVcQEf2C/V+9edthJuumhSOozP/56fo3gFVOxUGHBT9lsJk1lIW
sdCUfoalmY2GA7IYnUi6tUTGFV67j9LY7xcx9vL+XHufcEwwnwurRvgj1WjhFOt+
VCEtTXgB1leemcw/YuN+QfEWHIgOKrOjJXn5gC4AB2i5n/BhSTZvzFBQo+LFSMRP
1+e4ekCqzMff46FK5MumM7kxTrUN6RZ4b5nQmuU/Tzp7MeOnGSC2xkCDop37iDme
X+4vTif4HnzjPzziYQ2Am2C8My9Pp5QSQ3Mit+ZVCsEwT+8W4EptooNEnpDytXCp
xzklauQv39+tyUsxrf+CVEYAFwQWr1ZQlO3xw8GPFvXbX8V5x6IsAgimvKFzxDjo
yknsI/9qOujZHDd4nsNTN8/STnn0Bi87vKEm3oMf18XJa+1M/G/SL9vjhhhx8Qzv
w5FaMJUnxr83CpUwayqzGJk8zB0BUNTdUnXA3dtRmoS7zvYV9hA/dGLLzF60cT5T
t5Wf/NIc89pdG5IB2UBBIEh5F8n4leJVh+xCGcsOcoqbDD34Zzw4WZDNsGSioh3Q
Fiq/4cjWWgUtynZOCvjO4QiDR+eN+C1uT5HGwwP4/MX1w2KaxiLrG1nfMDH4UYmQ
yT1R0CkKhW/2um7UJwrJhNfPQL2G/E2KIr6LaYO9097hRb1N38+wmtF/gEinLWAp
HsEEu/cDQFgu+r0+6ep/LoHtxYAglEK/5toqR2hWEGMunxADk5/ddQuntOA/mHxx
iq1nRNBdq/pFIKmto67W7dXYY6miLgBtPWScF1z6LR/OP4gJZBUehHGRdMPo9lI4
raInz3ICmR8Y3gBQxq1aFXzN19czq3wAPdSk9eFbYSh6tdz8Po7TdWz/6YRjKQwO
zzwL6nipzorcf5vLlXzSpTmefwsjfy0gnV/z8bjnyCi3/MFKRba+nR3KtU45VQdC
aM5SarLP7r630KiMA7QqqiHifVGi3JGkRYJzSaeZxW+ASmI9xOeSWpbn5cuVQIWH
eoXnnNY6FO1K2/oAopYJnkikiNbd9pt3IgPIPdjv7de4ke63Smm9T3seu7STxxUE
ZYqmn8hwtHwlSAu+WaYbOy9ssrYbYqp4GRsyeqgo27fy+ht4OT+eJB9UFbLWPGi3
go+WjwkTjrV+LhJ6kETRPNB1mEivBR4WwivLjKtiVIneSeosbwbM6znr0s/qhzqX
5hkXYk4B+C3BeZ2clJesg9LPTrw/NgGkbf6PsfHtPXBpxCWUBkE7zB2PdRJvCkxW
PrKsQBUNQ3ImTkUCV0NWi2ie7eMgXQ91xx+DZsChleELnawllC4AH2vOCA6tG/K9
1JlHih+xpJ5m2kHeAHV8LERo0Hq7uPw4fzUapOYoh4FgSd9dss2Cnb2QidYG78V6
zvwx8iDjYnIf9uGPsvtlECZKveatOUhmRX+MW/lJ7p3k7hdtvHDIi772wSY85sYL
PCOTE8YVhKQN7UfLT5dIj/mGPtSzqj5Ayx+P+kZFKn8WZfBnkpNuq23Xeh64E9Zu
gVEhZCM9UuiledrWEQ59EsmT7Fi7x5TgpgRZuF+9ZaZOQ57oAvrluFFpqxRcJdi7
tikRWfj4M67P49hqDVVF90BwWxRzrsdxbQD7UCXzFSSi3h3P45Q1dEc2VyrPRs5d
DUqz0kwOqIuf6JM2XvIUjSSCKb71bICV1RYCH7Q8PBgIqPe66TY5GgjC/MRJFVN+
oYOXcp4xdF2aXyQjNcuCnhXAck6DOh0INPPn0gdf11FtS4JKzNXUvd3OtPciSSf8
9imXCfpn1CFAhJoVsKmYFNihJDffyDWz62+DD5sZf1JCsMhGPUUQF/CSCh0MJlt9
2fSZgl/Yy6gJioebo3r5BKxG9FQ1Bsc6M1MUZntBQdU0jXS/1SAbIlluWD4Kn0fM
VQeVmWhzq+PboXrwyJ2Yk8xmmISGzE0Gms7kdXhc3XTHYGKZEhhj9+90GZ2SjYZ1
gwA/P/GCItOnwF1e/qkDaKFfBf/VY0dusfyRs+dPultwvfViqjfWecgS9LKUIcG7
aBR1nBWl0zeqfav7IMOzpUT7LN6hLZ/0KFqlw07I/K2ayBzONkUL2TMhKs7HAYzF
ii5a26VM/nxoMx3UsGfA8vDbED9C1JRg64EOwwqbhpDZMz8PKrxEAfMsIwNNgqRP
6oLFGM2slul1dCplknV+9rOSQZ5h1Ny3tx1QO6DT8Hm4iEtRGb4AQ3gJ1GhwgWaF
NsVX5sI8k/KVAfh2G6xW0Y9kvx/Uo5Otnzy43KlrEHz6l79KPZhhKUViZ9euI43t
qZl9MT7ATdjiGiNFR20Su5PF/yERcI4OC/JRy1eVSZvv7+NLwVNIpfgNuhp7ruWE
rZj4UM90D7tlyqz9kefftyDlkMkNGQHSU1cgsR99Qx1YaO7T6wm+k/4cWv2EBsc2
Xt6a0MoXob6if56UkqRvO0nPQR38OAABeFZAHFiavjI7lucNaANBOwUMYv/CwbbR
2HWJyJuV9qLNeeDMLCx1HnrsjcXKM+nB7waO+BW/kdtQXw/r/CaiudFiSs2zM0ka
dX2Wo9Z1R+P7L+pT2JNilH231jHzvmBlXaVX6BKaO68SDnNWKGI23K1iq5TeaSyE
ULqcBldzCXJY3MUzvRxGWwUK3oz6BtrXOe/WYs4A1IyqE4SwuA5X9Ic4U0mRyjWq
vx1/4TRnj4tCsxUyF8vtKBxqjWR/y52ROROIY3KJIPPWB7RuGZtVzYHTasn+qLfE
6m5b2R+2d1/YMb7Xy/IU7Cs7ZBbHVWpi0Kz9IGIOseRyRlJ5rifjjVFDcyK+d3oc
dBKyonW0j7igQ5Ks549KQHDscUr0SDZLigj0LDzo4UM0CBdoF/PifUFa+6XZuit7
+qHXq6kf4xNFj12OjF73yZFPvhqkjSiJA6Mf5cSZOw6kWa5YgvI3vGnwRCZJRIzn
Auak/lT741x8LxS6D9w7qo6PoaDtQFTbiNYth1ww+HlkFBfqhzM8zFwMogulArIo
Hhi/UXYtXHk9S7djdzExl7NwnLPZqWDJljEcxRubqKW6ObDMMu+zDLNXM+yV9k6o
/JiAGqrzb4twp/xQwGqXk751PRincioUpJnYWlwS4tatE3Q8pk2LeC9znPVLJgwr
S5fjALBKXETep5lXSgj7wHQtK21Xv1CrVvOuVyys/e0a65VJ2gcatv0MLDTgRVCo
ZKLVBBRyt7A35HI8YjjSYG2vB309j3iZJEV3JiNZxPPQvKCFFR5ydfM7OKBR19vp
9ADW6xw0mzEjoKoHaKXHNNamtHLlDC0ol3EhUKV4Kd+mNEd0hK3rLAd2XwebGpOL
81eVTIr3spsBm5G3sqltk/DZpGuoinMLHPVrHh4lr/7GH8TFqrdq41BHfNkhP7FR
MWcWXeWjdMPTTY268DHKBKI3ttIFjgslyPNb7jKp8A1RJobaL51QSfiJStkzkCDO
q3VzZK79gFq/ZwVncbQuoYOMpRxPhfNlyP9dIM/ZRFWDJZg+buVJXMX5myxh+lfD
0oT1C8sjE/RYmO20BWJ7wdW1+UrHa4jz3rDKWrZvus7vW4/grywcdgfm+E/pByKl
ttKBUSJgtlo1eoytE8IW4vtYgqtDYgblDnqG8dioHV3CA18SF+1me0KiQwCGSdmX
XEvEUOegb1d2HrgyzIaabV5KSbh+MX39isra2Ate+VRPFy5z25i62xknkTD3bGAC
ftVc9TLW16JKxxTSVbUOi1xV4iE/5602yIruudTMjgtD+poeKMy6NfTqyS4ON32S
cI2H9jb13vUCs9LZueDblZrK03CTddCi6OOy0h3aaQZDOKcuNdQQZje7PUNg5W+W
JfxBbFJC+O3T2rBJz+bjSBZvF8Ba8VuuMVEUADXGc6ecJCQ0vOhMd0pYtKQW92Aq
Qt1xE73sGCZkTs21PF3kB4vlme3j5CfxX12bsLwM33VYU10yTM+DH5AChGcv47Xv
PXmGQyiYXhJXsSNlZJqho+RY8FB16lxVCIj6jy24b/5ScEz+GGBBGP7bmZo7mnb0
Km+KzbPIV0rvVBVmYK64wAsz/qBQbGGLs6AcynXOs7OgC5QfueLSwUTJZVSAKDSQ
C1XLqnMIZc40Ly8WjtG/rHD5ZoJmTQf1aZa3D1NnFTaC1nFfo0/sh3WsKBnSPmzz
o1flFmq2u63ZDbEh9th2A1T7HYdB1tOLysYNovOuGHFS0eVIZCXC8EYuNxm6zHVB
E7Ope/q/vX34Y5F9tzIgkdHO+8r1QLEXxIhapjc4mJwWt04VmEtSeTaoy25QDLbA
hnkgnZZeowsZQNC8hl42N39WcFuukqzaJHCaekIavcbYE1T30U4TpD42HE9cToRU
+7tAcKrnyZZLzdG6Nk1yqwFVK7d4fcO0FkCN2sGVLnO0cecroTOkgASaqxMfs2hd
2n1TFueAiDhn3Sc7kp6y8yh8YFhdQJZWZCmTZZRv29qqiOt1OG5sC6yCGUAjuBnM
1yexq5i6Ue3u4EKxhMfnmtcidlMsK5J3OKwChQIyFuaQYrzTmUmfZdoDUQfDynKC
SI8LtUuwpkPfVj5akZxaOmskoid1F1A/U0Yft0sOIR/5A2Fj2gVacj4rby/zJdpu
DIaGBqcnxa80iicsXn1iAOFfLkGHMA7O+4MrtitOpxhYEJnJTTvMHLiBm2/9jUvY
CegrjfB0pqt80+zLK0iUnQeIjCnI/GZBVQmk0AHirJm6e8En+fnueYANSHUAwZGE
WeRe96JL12qQHYzOW2eLTXMW9ZZGN0g5+VYdNwnjD5XsSd30acNAXvktmKEbw+zQ
GAcELHkWf0HDybGKypSjj5r2hAoqDiOSnl3Yq8U+nKlc9eoTDTr1QlyhLhW8afER
lKGPWOZ8tZlpJTHDVMMe2bvTtZaNsprLE8xOuqZAd2J1yBXj9R0WcRfI+fCMYfGS
GGiM/dxgtCYo35z0ujJ1iIqu1ZcnaIXOdMu94cccc5mghO476RhU93ShnYWfR/jS
2B3ElVDSwCRKZr+9O9MevWca4ft3edxqNO4PaU+umYrgQSrnhanVeGuhzAWX9vN2
VQvi+okGyMaYmYfsafrh5vVbAMOk1upJI3yiYQ9TznAoV0NIMasH9fO9Ct9GyUPU
tLZtNE920iBTCOo/V21RR+48Xf34G/6vTIkYd+PhiPOkuqVz6LXbJngB6MzpqbUs
A9aH+hKgcVDC6CfcIZUxVGNUExwAnhrANxTKjocWph+a1AkK1Kq2eWEJyDqVrBax
czj01z9ogLg00DwfUuk9YOu/U+7Xqv9z4p5XcQEnBmMRYSAn1NbjTrBJ/Bh9ZrUx
r+4FAcHZAZxY1zQSBBrWgSxCqC7qsc4LDgVrAX/1YQM2wRD+gqJglTsbfGLePVxy
giS6YaMqEG2WvtK5P19pODL+prUltoE0zxOiLH+tIIbuhEB52Ix/16YDyO2roDC+
X996AZuIwUZWQigbg+mSFQTk0HD1XCcuW9clgAkefGn3UJdpbzWu5Ag1ZHvQKat9
2BmQrRqZi0WvEjijhvnvYwwR+8Deea1Mafv+V9NlgZ9GSJPbthAfuP3wKPduypLM
kW3N/XcG0iOfgZftLz+xrfSEcC02GYAJjj7dgiFc6fxgc2njU/nv88EOjJASo0rD
8yykzeD5KHVKxZHXTKF1EVnW02f5vuGK/onrIlmlyQ3el//vsLCTJXNni3aKG7iY
2YdXWoy2MOo73dzuPk+kAS93qss5XHdKxQeyHKVD9XQAfD8+a9SxO5u7Wd9p7jsA
TPekbmLT5+CYWOlpmBJH2apQzj+dJZrJQG7qaxoJpQFEHro3Eef4hDRvcaQRQ7DE
na3GebNx9Cy9LqApVXIBn8wn2ZkwhMN0zbbU3wjAFH/frP1Vu+/UnyE1++Ax36iM
EOUXdYbbXYC5vW6e1jeJXCDJfIAqmSpO9IQ8/86FFNpRHqgldQlcqbI2qEiA923Z
g97T1jsrhnoAlri1gPPW3S50oK9f+VLgl0zAg21rimQb4O8xA4nQbbGZkypaYWjR
mYYXaH/Z9Fm6Dfo3Lj5DQPrT9dOu5mpNFSYdQ3FvTSrybWPunqdSuU9ZeArJFeZ5
xrqVrdJTUIU8i0sBV771A0YwQmQ1DpUeHQbD3lhU1ObBF2yigMowD0YLMurdDqhB
uzCC0fDF3nI4WhGu9uNHaNoMqt0rFAc1JP3gSocYC5yp44sIINg4WOwK6ZVWV2eX
YVcDlfvmPNAXglUmQL5ZDJEEznDMcRUyAvIy7ZtQUBIR/88TaGpUj8+3EuAsbSrI
AM1ETH5xT0mSZtmm64WLoMhnhbiUmq/CGsuvm47QwJCA9/GnZwvkJCJa8llr/a0F
dV1rua82s/U9yuGVk1VVYdTLO73qMDh5LC84tIiWRssxc6OlXSrQZmpX1IFi7WoS
CoiGah6D+1uTH95I4Wgq/EVNzqVdo1Zb1Aj6douBz7WAWEDmhK+MMHNkbVoqdOb3
7zEkV7izSMwmyFN930R4b1tTXCzSTDFsdOvZ5xViauOvgBIzzS4/spj6Y6VBdiDl
BqixYtZgdo+vOSZNPf/pnpYfsfGTa242O/QlC6KcGKzBByRNWLtkz62rMs4K9XO4
Zke77clWSjLFOgufQgreGe833yKog86/4430BrClutPbVlYdMV2X71yoHCM7RCUC
fa5crjZoq1Ce9ViLGZAYZjy377TM2YP9vcpJMDL4y2urIztqwm0Jlsu1nrfb4wog
kCDlVgkk/sLV2KvXAY1rhtfKyOlSMMljUc2jNH4P8fNyVRPUqmbRs/gpG7c+XLvb
RoBYIKgDPgal9su6TmyJvKhp9/vPj7RDNl85DVx1MYIR5WGEVX5yuGsFjP84l3zZ
roYR7O150lvNsGFzDJgHDYpD95ZJfvPNDWv0oOUTBsOadkh/whDbIYX5/Ikj8FMe
vywlqqwQ8oEitieBmFRNKc6uSeLAG1A7iychDOd7kSwh+jcXqpk9W/IW/W/sv9Tc
0h53Ms3+XASMTQkM5yTNYMAJfejoES5uIjiSk/qUHEGcVCYLPN4jJu1GbGG77hH2
BtFiM2aAzhIz4hrygL4JbEbfTv7FSP4WDdsUznWz8gdj1vVFONt2ozwIknuQMYox
rWVkzA6ghUbdRY2QGupeSDp0yt64Ty+Z5Tev5DveqQ9GxgDmZdX141HsdKLM8ijk
45SnKYp2PARyphYfJkd+P2p2a1Wfq7c0HrHomVeS+voizmu50oD6RDU/h94pohPM
a/eQgSF9KrsIDzlb1abRrZq20+LFLIKHJRmuy/XLpiuM4gXw5wEQ38g7bbfYetp5
+89tF9D7mvMqMoK7w4EIvb5cZm76c+mgiVYG5pfC2AKWOv5RMD6fAdBmvTlcS54W
5i1bgiuT6Ygx3n7WuMGJWRWBLkaPSRSjnxMewJwTAj5VuUZ2g0yEQ2VXY249knfH
/HgLNZJbn4WQjmNxikGPEPKQqPjSoIcQi+rXvzbG4IlDLwVw3YDHrJ1iJ/16JQIk
3xug82SnOtrqVugfxGAjJcIN9sr6pTrHJW/Oyc4NbdYKX35foIcwSuXt/V1gvdAS
KP7MPrI68GIiM4pSWNqha5dHaFmh3zAAfLyU4q2zsW4uXluvNx/uw5iXD2PPrZqE
B1Kdp8khLGUbZcoWEiNWIPiUO8EgZRE3WoNg38tJylrRX2A9ESqO4t/qIynU2+Zu
1i/3OwaQrq8Nb+rxqKS1OXLXol0Vt5zwjPTsruy7A6j8CpBxotlXKRueqtzSQn0P
jdObsQonz/PO2ViHDVbSLrW4fBLHduQLL7oXic6jARhb0gwTPczpdcV3i1kjMr18
WI/dikHfevxx9Fn+bTpLfPdjHohnmuUdV3Zk2FJT8jqAEPcBFIMVSBbLnu5tggit
jhZk6+q0/0swBL4n1gmFiAmeoLLwTbytqW0a/rapDKyyNX1piMo4CnWYnu41j+Zg
XS+MaRw/ak4LqgrcwX9yxQfhOs8k5APtrNLenJN5DApTJpcPChDm08OMKOj0dTni
114GyuArJPWtnbwoOWDa+1bA4v6mHQp+1AdgstrMMHdT+6KUk5UMmML85pbrzde5
S1aWz+uuR1IcpejrBQRu0AJ7EZ9Y7a+nY+qvUUUis2uDoqZ6ranOs4yseUbm4pQ6
zsXq04RbtFYD7HEKNeliETuwjEsnnbTjCDcuVWmGmtlrfLwzIVANNNPK8jJOLQIH
XOtfWjsckYEixS4r9xmGZerC6cBiprThCDc2osKCKXAsrVvdAsiSvUPOS/QSRzK/
9NhHZFpoeCdoKwgpJSqtbphMTTOoSrxPVo1AluPy5SrNq+TGqAw0sDoEvXSBHUol
r6bTpJX85/x+r2TQIq8scBDCcZtsMEGUXpwZS8g3jq/vw1WLnnz0XVt9wze83Ddq
9kWoguG9yfhqYwTWzrt877M9EeunjkWxJ5cx53kHOb6gXZ6YuqAqxsv8LiN616/E
6kRlLhvRbX9dz8LXHytBnUT51Te8kAoaglErWG7Yh9VUVunW5CkJXD1ev4hzJAZ4
5YksNEIA0e+7JsL5FrP6K7djJWiIKok7bxcDnvhdi3gZuOpCCMIHmj8r2Uv9rptM
JeZ5Vod6Ke9G69rSX2WvtUuG16ZU6iCtuYtghKMYJuS9LOuLDhQ57gZnDCCSfkQ7
+AVyvUW7yJpRvB+vwTWFYBZkgmRolRBJU1XecIRgrMyB0EaIMTMjm0tadIl9EiVb
4wpNz7hdrjXJWJz/vfSiyKMCI1BKtZD+1Mlz3qRButMkizvAsG/JIZl7OASUREHt
73AkeJc9v/kKUPYUtTozaOSdMFVMW8pQuEQ5An9WuS+e4f1yNp3SaEFP9rndDe5c
Yiivn1whO47BtXUmmXJzSKSBOMlpTQNHbdUJ5oZAG43PLyN7bclJFPLpDIbPu9xY
1mfUChtS5Tu/CJtLOCyAjL3lDxt8vikhy1UWkJPftMcq+c7I27oBcA7eid5oh+KO
eXiruPxinheYfDPcFpnAtrNAxgtBGzO9w9HdINgzxCyz0xjARCI13mOcb7azIhgt
d0vnXmkXbAeTSAq7e//wp6Ho6PVp2uVzTet4bniA2miFZufZPINkKMK7slUZoqdZ
WaiUsG5sG2c1aQDkbnWwAeOsgBbu72qYZINNf98f07O+bFLNUoWs1wXaGIPH169l
K8Tp+6Y2JlhvsKjEzBSGWIxsb6BXr01+35WeY2Gyifu28cfPBgdTqRjj94/HaZid
LvmMO5wz+HDr29WT6gRyggUj9oFkCDe8p0Y62pK9k+EFh/WPJBJINT9I/rxdBIaM
UGO2Y54BP3afkNZuNwdtDD8h52rXXVAl9+IiCpc7r0EYo28gR1k8QSWn15ijB7kX
GpvI+O4OjU5524rlsWK3To/xJxgUoK16f1gfnuvzh6mYlp5Xi73qgJdie3R0VRtU
tsPuy2XpDshOQjWCuNsT2yDVodOzSZfI+wyxTGmOYvRyASyJt3pHnAxSDrQFPljh
8MCb1VkNkPgTjqdWucUwrgB74rrYGIFLCftV1MHHWdgfGfIeNjJHah6NerTSNJhS
oKYFpq8GqD/pb4u/PcxugsXKeWBSmEvHn0prjp0H6nfw5ZuL/8ou519/USNRqkag
l9cHnhdAAUBRkS14bpu3L61bppr1TjWy939WCdCnmO6NXV99OanbZo3HsBpXVFcp
wrpAu0dHsWtQeuhz8mGdFjidyyWFu8IQuJqxBLj5A7A/1+rLdl0p71p9vRNg74hB
36OdwAvAMtrjWo/DrWPnW2xc8fg8ziOmajFQ5/C2L5v6eJ3XO01V26KaQSc+WUZK
JUDsbXIUCmWXaxgLIQgeervefn3Jp5iQlnQvVFJHEyU22OYB6RJk4DwDW9N6ulsp
DT8tQdjWrsSaiUPOtjcOpe/TZLDani8a2sVd362lpc80/VOM3vaCwdd7WJc/LS6x
20Kx0o1vuf0X4McZpvEnjdi4h6VqMspPyPLv/8v8U7eCi4MhEVzLQsRB9TTyZSut
LQU78C7yQTy6zg/OWMn9x01XHTrGsFvDecUJK47cUUPiLGry9D5aZD64KtS9CJPq
9BqwPFw5ZBjf4HG2W4UaAUNhIhitvHBd75snr+DczcJOg5O5xvYxTzr/YA/DswvP
PVUXJtALVnF6O0rIp8eAoLdNobUc/LTfz4PgmIuCbD0OoodTaO+95uqVWW7xjkwy
TAdlP5OnZcS4V9bnvsJLR5TbroEfz3cAZlu2hL/4RTXM/ssXQfZdQ5U1zhUifPzI
ucl6RtyADBSEsXW7qv+nGlK3P6TfMy0y2ehVq69APEPHinL6RJZMzsxIv/mb60AV
qXBxqtKp+3tqodpeBdw9Ic6bFqVsonPHi1s0o8Ho2tc3voNqczUOOhm7OID37ljX
yMu2dICyibxVRK5f0b1Gm4iq54mJu2hUFbnJzUdQ3Pf/Sy+/AMji27DExekhV6YP
GbN5GHgl2c9huvPvBw/y4+o6lluLrGDsooQ+3YzyhlTwCwD/LgcrG++A3NWWiGVC
+52clJ8Uf2gK3yaW19HwVopzfVImBz8THX3fp4qmrzA/vIbovDyYUzrf9EZErvLp
PftaJ6e+goLZckMJevxflr8Y8wTIGOxZDjGUV/GMeq+OvDI2haA2p9v6CP/iOxIb
Y5J2TipiWIat1jULYxzY3EiG0Q9ExtPwYN852vc5uLNHCu9+nR86wwsq1sptQ1/G
DUhhqdB6BSQw65Cg3HaR/sBh7+znX5inzYa+OueNHFhxoCRIvqh32YWFpwMDZEo2
YQSvzEoPr4iyU7GkEfuK085WpJDa8Yw5EnfecZmNN4SI876lfEPVoBpvXGd21U2M
qGdARlOhsd07z8ihylUBuaq0rRzaBLGlfIbpEOPxxgwJ91Tb65aoYcb/l9tE738F
OBoIsyzBevk2vT95b/aBH2KPXjaoDaJCpt0U7loZd/Tab2q8YZ3/P0hVm7WcBJZ/
zI3auwentW+0P3TkDLZ5CA9yELVbovSouhdHqASosktfq9QCfnN1y8qpKQcGHJXU
oAjC2jncNc1CdSZGQDuNDF1khDYH7m6/XGBHeWVI5rY0oxFi01yVxI4i8QZzP0zi
rsIQRA4BS+qyDwY0DC1BCRPLqXyZytn9V5gPtNCZrvVB3V14Eq3xy4zma9J35QBY
Ea8qcBFVvAtHk+i9CSN+e6geWPNxh9CGW+FlOXAQ8tFeGzhUXD6XnGHWZh6r67EB
cVTMIJ9WQ0NybskAzFWNBXIDJ6/hbM3b3pDwxzcV67YcKWQPeJHL7lGLuZPfQylT
jei7P0KfgBYGjfZlGy6jspQVUs5ypcRDolq7gdhQGAQL4la10DDuqvXACXZ0hl7U
Cywe2UO2tf7dhkD+39GR/1OaR3TGbQdfUAZwDuFtycetrvO07VysABHC4mF2YTcu
84fLdSL3/9ny3J1u2RhKYSFJqvQUK4OPKFlHyLcuQuCEnjVBKF3jD0pwxx5rijUJ
oqynECga79DtQniKd2HoPkPfD2wzVmTBXtupDoh2TeFLlxC9DhWKvG9k6skmBaew
N+Diz2R2z4ehSp4eDjWTG7jZPz0nkA7wAJDlh5TwIweH654ODzqu+pLTP2cZuGrb
EUXZz0p9hsYjWLk+9SJnynmWR4Ti7785rlKRn0SMvEWfqPlEx/jOL8dP0Jth4+MN
WO0rYZcdXp/YdxwA6knIEANyTAQlyL+6QeR0Q/vBTyR6e2gvKJZ9SN4dDgCfcaCG
cwx9ZPKw1cvo7VDKyiRUIflNCYwKZwgOyU7F/TcsOT+OktWVQYERcl8Ws5iL1fR7
uswXB/ae4RMQA/Qp1pCwOzKXXZGhIvEstvm2zUEIna79t656TdkM8zlzcysdAu/9
xSKsoRD8dsITwo0q5ckqXn2QxGzdx3aieUYpQzKiDHUkKeFBitKDX0P1VCev+p4/
nkm1UO4myY5WSrAcImmV6GcRZGR/cBDQmb1KTCIkyVG6ZjFg5TWFZVNvFEONt15D
t3xwTxgnrWRBeyQDrlsVl24Rb4Eu6QVB97ms1pJU5OWIjFPOmZnKiEkeDgAc/O93
gFri1j4w6mgC3aTA4qZ0VYMc/A6V1AY2YZrbHsYA7MHBOmr2sqkev5ZjHKpVJGHE
nMdrKqr+qO6i62kjKz2hjH6Pt/bn8PASK6gq5rondAEfNNv/tx2OPX3NQ8UWrMca
1amYp+M043nPor5uU9aJNUg6t1g8GzMoD/+IK2ivyh+obskpdEo+cj5IHEdApKCY
XK4hgOzX2GuVCOf6PvL5izB39W2pMZRP1Jb7k1pKuRpTD1LnXgImkYjA78xzarW3
BpBDWQZ88Rwnoi9BC8+zQUtQdH+FYNo7Tbg2IrnXcpcDHjGk5AdNOvEWln2QEoLn
CuJi5sK9qQ/nNJg46+c7jMbKbFg3+OUpHb3c+seURFi4DJ5ANHKQCmNRm37vP/re
kw53SzXY5ed/JKDpDMsyyl+02IJnqUS5Z4h8aZAlasYOzbqkEgK1r0hgQf7BA+uH
i+LPFgWtFQsODYcS2FhenycPGM37iUUX6WKUfUOuu4hSAg0AOebgYR0Gd1hTH5EB
NOxiw2d3s5N9eqPi2AJ2iNUuJaLzvTcKrA7Lwe683sW6RIJ5rNwlryt3FDa9zljv
IE2mry1erL/XEltbHlcQsZ3ZBJRpGFpZ3z6TnTXlRpoGR6L/Do2WmXKawnnfTP4i
8MctELugcVIlNEN8dSoX+CDfCykoEfbodyIReV7EE+YEQiCZEar1O1AVVShNm+ZF
tCy9KGMVpA/6e7Ld9Wzq70gbjsCw5osyeLfJxXATxi3PXrixQSBeuuJR10vVSp4R
tXv0XvjNPK2vAmyZpCiBqrvgRRs9JpGH+BOzdwAkr1EBTcD/OwM9WOuxjVpOgGZw
8FcopWH7u7uopYsc7W/ANsXr354RA86QLet8iSeMRC+MDO+xjwTo7Faum+dm21qm
itfdA3pi34Or8vBJgxo+W9sfRBjuBIeV8nIHMTpboc7v6XPyX/CXUy9l5ektUcVW
xwdJLnrRWw9QoWVYlqToWlDn+oPSXN2GH9a0bo1hv+CxhX8QGu5TZVmp56KcmVNT
M24ZKrCpu8G5xqtlYPO+dCXVCejQWdYHOG6PBYj1broAZwtYdNwEhCNmmSFbI26u
2ypMiUKNHpP6p+jbp+cFNF1juoULG2t9siJK4GzMzCtsz19NfoPYextTqxdJL0XE
968yvbsJlrtX+fye14BAGbiyfDdw1rHd9I2K//zXm+z7yZCuA0hlflp3ClXMaIVe
2+I1/2or91EvNeRD/W++f48qtnlVPqU/EkyvRP0JQ94awY/TWVTUGucng1crla/s
xBG5yYEvqQ3WvY5jcxaL9hHyvj0NsA5XqQCAq/x82dw9JDX89TLlkxjxfZ6wQ5P1
SimToXy2doBZIMe84+t/UE4tpZ2lBebyJfwkdd0Sk1zySCUODT8MgwzXVMtByAUi
JaSpzUD6ukvmsrN6JyDyf7aIZR46CNqVLeT/893IeUEyU6v31iNjdy5y3+9ycsRL
GlKGUrLSgsCNO6wOAdQP8SUDNIfUO7+H+otkakulHBitDB8DZMOsrwjFDJkvN2pw
uoTQCrEvfPCa0lzhOf1SSepUHLod82J3Szrwmd7rP+Vf9U5UuD6iJLIVS30EXA/m
dh5e14vOl37/HS79Cs3i5xlk0ZH13zoMW7X21rUol6WdjX9MIRoa8uDu/6PqeMcs
oEUdtYlKZMV1af1KzovZC1ZLExXGfl7m+/G5FqZrKIco8JZVqaui3jISttjJqqul
Bu2LisXoUawIT8+o5ffP9pAefWTlLcwNFdd+d84VclZbsKfPZxY7vYobEa7W9ui+
1RqrSD5mTJ9zD9Ua7dwokj6Ab7TB03WX0jIncttuwQ4p6c83Y8ciTXpygpm58iEB
UVyd+P3ZeTZqv+dI+W6rUCmxotGQLZDXoEoSFBbot61jDcGK1xVDX2asXFv+2cCn
2PEuBhqoLRt/BCO+X29Hnw1HvzMPSCIKk4Z/TvK679ZNqZCCImQaw3ZgV98AN35u
4cGTimWnK4AMVoDn9YZ1d/uOCYA/6iK7rOSrURiD7bPiMpubn01zdErbyxp8fO8y
CmVgd22z3EEqN2vN34Qw/erkIA6y84TyRu4nwKs7QYXWg9N6cDZwBq8jzAH4vEdA
yzeTVc7kGaH4FF75YxlGQsZUaGhSq78131rw0cjs5L/ejVd+4wC5xZ/V6EL2JZgP
UAXSwEUbg7Dwrc3G9ML+1And8rYlhQUJcrDHZdqC01nD7m35juAvRSppp3CuFpJE
SKcAl9LZzo12K/LWKFlPUS+DPH9S8D19sYtp9WTyxJgpcUeLi2/3ysYcEqvUuw52
YxljG1YFDhlxylhYDIg11rQDk9o+BPF0QwkYhY/W70ukDzPjVt21wBHT2uII7GsN
JqUI06bEfVE0tryxfeUArYpw+Bn2S73uJmmUWWDaD3+tbs2L3oqwESjpSUre+uDn
uornSc+beQbGxeuVfCa/DiPh8YLSzjmeZ9noRo8OxLoilwZo8WBXSw0VMuhPPy31
wu9NbZXaEYj+XIJ1QIffCqqd+MPR0+j6I9yRROVvZvCarTsrsVMn5dJLAlYbCA86
k7CzpIfb7IeFMHUDTEeEHkzTf8GFpZjH3H9krMQtdtBbUUyWAOI4jIsJv1RHEL8y
SIDpXvuxjNPGOaiEd49YxTJd9kdd3PSyIMA1R21fXHyrOZlCDySZo9tz8QmMsaD2
GV2I4pNIUBryWahsFsItKUUIWfZlJVrEE4Xm6e8XtXyiKjoVa0DtVPaZNCF2akOP
9Xhi3de4+WZCQ46lKWPI0jJ1ZJaoePdMw+lQQVJ8zgBKEaU/9jZ/BK9LD5VPBaaV
0bUT28xeYYDTEQOQz4APEbMbf2BwGOL+vpjdWyCYe9Uss2Kf3FuzNcKf+8xClZiM
jOuaQDNDaAWz/jGptpF2G7Ne54VjMKTmNXnuqqzLisX00xJX0Hc9kU1GIex5TMwb
QLCkefi4mXk7W1DiQEQZwu8Ih5ax49v8TKI5Lmh81B1pferX7nfD6EeW+cqj3TEL
5hChUIDKkS85p4HdAEIWzX1jtQrmZCh6XvUw17tl/37E7FycSpc7z+ThnKHgEupy
Ay1l/fYADsjprf5OnJq2VLju63H1KKtrGvC9Zw8JEpsykon3Y6fHHtMH1gUm5F5e
IQ5ra/B9eQvX+cjNHNxy14lqN76UCQ2kgE24+76dWypbuh7c8fnfG4aTcgsP7f6o
yZCIXzKWRXYOEBWZPAUIhB6Sm3ZZqqpVMvm20X3PekASaCsGvyuV9fSzUpl5NS7M
qyeU3btr41SgwbD6RpfiLMEpGGv3iLLofPifYsGz6OooqHyiavy/rQcMb25SH7ll
8tz75Q7+veqChh26koG4nGSCjr4Tn9z10CnA8BfFqj3ENRpDJJiahuEOUo7YnmCB
ytJ7fB/qiQFioLnkNxcSco1CrKpq7rqkcqjhHx1+degxxbv4yoraqSajIqQZqGUR
kSsdRl7X+6nA3kiIzIznwOjKFasVArm8uUIKErnX6JPkunSMOTRKUvPkzvxFGBnh
AG4KAJfIITnJL0jCsjtR2Y+sZ97/4sRgfitzuh9Xh5lYlRXMmkdFzIRZPFiAwBzl
W4VEMr/9F0AH8oowZuoV1r/Bvkpo2FTspuIlSDNiCo5pUlm+KoBREYZUPIXI7wqA
YES7bgw1Vf9e59xd9xSB2KmF4zZWDzpgDzImo9puAAScACY9O1+vMYn3qF6Pz/bM
133UsNO35bzFm8OBUjuYQrjoujg8nvGjRmt4FeFAwqU9rs/b1hGYq1YOBr90MvSR
L/d4X25unahNiJY4MVWl+O6WqBoopoiU68suwR4yzkbjgEQZlGOQmjSJ9XTTWDe0
qBjo6TRfNzkHz2tuJ2hWKUMARSzalM7YdsqSZclzWJHjSRhAfRsf7CpXkcnDcrAa
1bwe4lHzfv9ukBQGdWUSqMFd/TG6adGhWbS+lOuJm2c+7f4sMw8JMHQ3OT8IElko
8RMJKpm+quUtwEFh+AEqBTUe+17ID4Ds7uHvSahoKWCMxB8XVY82abyI+vuku4B1
cr5om8PF121T+mjSvUNy8Kml/nES8gS+/1+TJtA1nDDi40tF+aQrj4yKV/v56lCB
Ec0JBSoLJ+0Tmzwi5Cj4JJ8ld1jQ+VcqYekluGcZqQmQFif9IXmQ+QeYE19KfWAw
hfS1ZLXxGuXu9xhMFnBScVtEuYslAF/+wNgebdpxNEa3k73jG3J0BOJWMq/waQPw
1zU5jw/Ac+/5ju7+pgVJMZMraJgsY18VH7tSK36I55ymgnCOcg14J5K/wWLkxNIT
5DRkYEZarakwOYm2EjLE6F2QAn15FLWFjHtKC6j56FyOFXHHkqMJVP5NBROP4uIq
XqVtSB1VGsn0zQIaflsm0+zUstCuraoKv1rdRTdM53xCveQRPno9ed9R6977RT6r
lTcnqeQgBqvOShznkongIBe0FHOcLYpP/QA8seNNnPgN0+/7QpquYEOt01utcvkt
d0pDOGuM5bOEjm9VQGfN9JPWFEHTO8ZbZ29C6l5crEGTrv7MCu02SPEcEC0GZb/E
3rFv73cd72NFp1skEnBQN26a7Iw6Cpl80aStrdPt2KWNhaPW36T3aKPvSTtouKfD
ZCxqEFJVCLgf1PEtS34p8myOQMwNH/zQKlf3JiUz7H9hV4xXZbig4LUymUy0iIg2
1Bb70e1VigX38F2yzrFzNQATYbt4wn0CXfrLyZekBs/K2fdRu237fOmq3PYfxUx2
aaja7bmR4I1F1fnBNFiTPxzI43bFPyj3WGAwHilOL8rv5m/qJS0APxuP6rb166Vx
8mppOuw2hxlRf+4Gei+Z9L8wDaqP8VbIRA6lK5FAd2VkNzIr0z9k2f4ficDjW7Vr
o/rMG3azjKbPHMymkEKrvg5peIJOH8azSYys81YF2KbN+SBjpFlIYr8rnqrZjkXA
D58yPYpN9n5aX3gfDyUfkqMbACtLfzyrz7ZklvN80TqCO/RaaawThazQxjpQA8S/
A41xCic4Cvn7w4/p7yg+nfroHzomtqqatO8/KEkRthfmCiADEpwtYat96lNu13im
Ar4GXpdsMOcz1sGIUMY1mWsBodxZp9PeZkPA4+O4QJ1/ASYxeRtViWlJRU77e+bW
fK9qFoBE9WSlv6rxn7aeuQ4/+pc1gcO0K/OgYggGS1iXBqsArySqMW8B/pS8PRDj
hXFWeqGFheaRIJBEdYCZQGaCyBOWdHUbtYcNgoinscfqCEhKjyzesz2RF2hZijmL
YBKO9atmbVOBaxeZWQk9/tp/tmqaisLrdAMoiDiceplYS3//Phid4jtZ/ebwkmFO
OwpOyRLjT2gTZLg/7HARJ5dx4187i2fCM8NZs6YjmVAzZgdQTaInbeUjVsrPpdQG
J1ahfSdD2GbopgMVYNV79w9ZVnsquXeMqLB7G6HwhJiIb2ux8RGMe8f+35m+42WM
o/OuaUW3eoOmRIyMRRI3xnDaET7YG4o8dpDEfPDnmAhJlTWRkvwpAL1qRfB8ary9
jzdaHAZ6oIh1h7xuBNr24MTAKRkPntc/p64NmbNtcJUmOKvBJXWYhY09Zt/1WKCq
Vezf5sprOwVwy6EYO9R6/XEH7Timk+IwwEzpDw6OnhlCV9WzZYeE2wffVO9A+qmS
uxy1ImNHXzZ9bPm/rtXndSySq8NRjCTGxCQeV//4QAPv0+A4+8dQN9s7GG+h35vu
bYILp+A1Vipi8meQWSQPUFehCPH0Z0DpXJ2Q0kxUlnW1cGNsmnYWoMseHQpASGwT
M2ReO6Mn7VVFNdQtcOHqkfFxgcQGIyngOCmUMcXMGovdyDfWviXQb5b37/1/qRSe
/rxEhokJ9il5YM48lxZTcY6JVX7llXkzrasz6qDJ05+t54vLigLm9Xj4xNuDupQb
kE6qMc3TrLEA8GlTjpxMeqgidO07kz9hz7JwuPtvMffaqyIa7sDHmho/KUfXSyFL
irCfgkeju97X1+YHSG+Cu7OmEGjIHVDBTUioBlYH1paziFlRFuE4IlmAm4rGUkMF
rZTAwuz06mRRHB5lQwe8kDvpX8I/Yq1gGPSHCy6Vu9xETfMUU7MrPJf2HVkUIyfC
n7qd5hS56ripxHhsNufz4GGQRGlT7N2AGOhuS86LsuMZzJW2cO4TyGr9tEgrDCNY
Bm1YnzYkkBcSLGyFC9IVusuiV0j+U/X3IR40x8TUAJ84kI++R/7hwuJYHJqVQG9n
4/nM6v/BcAAeYiS67oVy8uosg6Z+mImB/W6ZoPp7JgCunR0+Yb9RqXub0DCm6DY0
pGrBVHYFjG/EIxmlYQckVYAPljNwqvQD7psBtoKCoQ/fWKSmCbUCEK4B6J7cTRMq
Sa6IXoQHThyw6m5F2dJ60rL3JA9QiUqosOgSQWspxXLnvh9OUxyS6BL7e+8ZlKJn
/WXN4x7XfKC3MqZULafAMZx+fLMg5pqZone7kBuDkSW0kOPQ+lEORwLOL1wg1+X3
Kz3p7omd0QHDWOgO0JOeN+9t0HkoFTBVGJNeoG1hJBo2IMwmPMOuu9ztKr1FnnZ/
Yad+tuhGqLeoCiDzw7ugqvS8SGbhjhqCv7OD+o1/41iSsCgB2rTRmoQOBU/EyhEb
YHqlMkFwld+CUgfKOUJI5qm+Ri6kI5CEf85CNGLFtm6ht3ZsGr34gPyw7Rjgn2Qi
M5/VYw+HH6ZrebRD02EAg91mflGbFd15HdW3ZXVRMQPhoWsDN0IlliNzxkdv91pb
Kclvk6LM0aslix0eZV8gd7Geft1U/5UoEiJo7lyFDL44T3upDBslaZwCLHpNX3h0
BUfLkzmSQ22iUjiYYnjgMl/b1rPM9GZHxB3hEydmlEdTKppYIXuwUfbkwaLhlJf+
eHsWC43P26bIyw0XpokXLbejbd7bi6WkhHTKIjtNjb/vq5C3s+ygyNt+huGeqt6H
w6FEK1BHHmGdkjRQ+ZcKkPJvcmd60bjMjApNaDs1WB4Z99QVJMGDX8MUOfEkN3KQ
NXuro/jHT6tg9hhymkXCHEOlRt1XuFmg5bfVm0byeWsrBEcslEIeC9bGrIIzKuUl
KY0bpw8MOBr6Qm7kxhKZ+YRjgeaMdycnOk+Yq7NTBbAxkrVQZa+kvSBAbaty+Z3i
uXah9G8LD9zfaYwQkzdhtWMnt8quivTgx82+pgbeK52LRR+j1rfzR3r7Ukr8vNM3
6Y5ooJVvSgGGpXAsSCsjv79wHFX3tYhQB4zI2CeRVisXE50NgeFPX81s2pypErjF
QoeYJh475leanc1BKjz5j04wuE6EmTocWXlUJT22WnROURoiZGUy3tIRMeurvkXb
qN63xV0hX/NFiWW6bupMacBuzki8enJwOamDcG5qa7I5P+3qSqHWTLkhpc0ozsbi
Q3tLwceOp4Dc4XPBmJ5t1V9wEmNiWRae3xb2DMXic0ju4sg2obE1YhgdYkleQHoA
7EJAgVtuvuGMa22qpfT59+P1dqskg53+d9RM/GGkuwHiQOuryGZwzzjBnr9/v9zB
eIWfDJlFd8H/NvpAZ9NSx7CQT7B5AcoZh/zLyZKmk/CxVaSqLvm/25IPwNCaTWwi
P6WpCv0R6k1k9/NNJ8euP5d+/Yoj+i2jNe40/VO3xF571fi6OqDmxTaYR4SBNnUN
6WWPxewvSV4ToeCdvNJ3Jf6IM/KLMaZa/JkqF0JSo7dUuziyuZBgbYw7eenfp8d+
mB+sBK0HJOJWkAORhs64R20ssuhm3xh+zPDf9kSkuWDcOqkUiuizMaPgLh0sdBA/
HKGoiWk6zf4343cM2pSP1U8fShWT4L+N1kQ+PeZyCoUITF0CeKJyj94/cWXgR/G0
BeDK2YsyJi9KtHFHAdw38jUdT51BQAG8qok3wSLTJL4hnVhrKssmG7b+mI8VfejG
Jv3+WAUdnKMZCMhbw3Dh7kWeaO978zd4kKfDUF7kVk0GFDdWzkuGXNmCI5ets5nf
zHmcsfidK41eDJSGeKB73KiErYToxUNzECe/CLMk4vMTb01u9nYOzaXmtvELA4sX
z7Bj1ITjPlyrdBv3AqMiF4FozM3vfwZ+vJ8cMI1qrfJh2nsa3Mea3rrNWgl6rbzz
N6fR0yNDImPHNdI7ykvTVAPc6TcQrruV8TOHirZB4GlBI1xmeSzsN7bDS8bWV9ZX
lIaQqnUXPilh47grXDtmNK8GIuZ7lv7sIJ/Sru2vGX5X2VK+lJpEq4QHVtxpj6kz
hcLU/UqYBXPY7Ddakeq8MivRwNHnNUbqwsHf0j5enTHju2maq//czEWNDqmdc+d8
ofcbS+kGTfulxU0KZthbunDXjOLjsQC3cYVl1XK/98Ll9ZYzpZxuq0wrfTKqG+F6
5uY9X4VOX2fOM9mARCXXCucSXw5csz2wT0paNdxohoKsPVzftH0Z8Odh0aPCx5kI
webA6hYG2WbQe5Bv9gaN755ElGDcS9MND2nbpkni9uv8DnCvEi4t0lxrZmSxawpR
9mkJCUzzjepkShmRgFyJleiTjtasm9UiTmIsCB7B7HhSOOnKg4sEdld0o0g9huwM
uwhOvyue9Fk2LVtvK5Omt402v7dVmYBJgGNswX+zgannIwHWHNC7cQxUM65vF/10
rSWaOwWAxWmrbADEKC9cGAXHbmlEFA1vZhWbm4FSqLZJ4lipGTtmx7NB03tw6Hia
u8bcbsOrFxZxPPr1gGgqwXr3sowIQdTGkivdMVso0JFXrcCuH8gjw4klkZ5fAFek
b/FX8kMOxybpjfg0PZf+Kn35NS5tqdnlb7yHk7ueLxu/dGwDRp4Tf3HZKMLYkoyZ
LkpIFWmdBJonwQXaR3z6DhJqztzpNjDdn2n+diJ3l+XTK/XxjTFPMd6k1sPOT12J
xNJr4LQSQ5xmvQcj/lWAbwDUVtW4G82N0zNarPAzOxJ08uhxnHf+YPM2xJeDQUNT
zZYUFqmsXI+fVBaQYTgEvzkXTt3RMUyIo8EPzoNBjxsN/Pobf7CXwHdDdJiH861j
d0OZAwjDTdb6zJCmA8XwRYocopKGfpd1YcudFhxSBgGOon6SbyxdROPxHZYkPgfq
CUkuSEF+XzAR0LvmOFmdW10QLpou4glvocHx2hhgUPiIvh0bMsA+OrkXK8PpSm72
AZzJZ1m64xqIDeX1aq9EB7DAhfLMp8dRKVNvz/Htww7xxCvJqk0lR3ob8nsGlwo1
A6JGHdIAe0/ygfKJjkTPyVxCLcp8CHL2+sJD33qnu86L8wNTi+2BUpK0ZNdJ2JmD
GYd6HRFVtCqDejtLu0QVgKeD6lgto+P+aOS8ICG+0oh2oZUSpUQDseAMG7bpjRUX
d0YSOQEHy9luyEGSfDfU2dKF75NfWROd0F6c3Mbx7KX10MTjUpCGLiG7kkROYmMx
XGux2Mn4pX67v92WcYeysjl6RUQl9Lc8aVFM19XvB3aS90eC5Y5MEj9uicvBUDqs
8hAz1ROf2lyihPnuRh1A0qpxmfay1Z0i/eEdciJxee/vkXekE9fOrsgGCzCdOltD
EaVAcAFNtu1Ia/eW/juDHmHwaCiC4GySMyMeKt/u61EeW2NAmjLlf8EJMPZVxxt7
r/hPO/3UB/z/dQMd5ycBVJ37rXZKUM9VeH2Cobe3LN+WIWeeihmEMP5nrr3T4qYa
gIxnLXbdso3HPeku7nbJfaHP9fSteS5wAcSjXLT8h5bC5eoRG83rJ1hKXA7fPhTg
6t91u59v8ReS+gYeEcXpnS3kmBSLemD3fSprpvDCC4uTfsG2dpr6LN3372bKpQPm
jUOiBRSQSTE3MNcn09lfAjAb8bdLKY8y8GMBSDyNPwbXohvOLRj61yXdqxdrIvxF
5XMJvIOrZaK40mzOQ2b64L7OH4PzW5CyrtC7987W8pxAPQcg1kxaxqfY0Uj5CLFW
SUPLjC1HG4VqIYfqxGMvKKwmYXghkH2+V8rWLRyAKleuMCTNRCm9i5P2EpyEpc89
LHvzuhbD8Qf958/7BjzgeDkeJIbGiLZTLwvTIAJuHtlxeuid8tu97M/ldTcBKIKw
60wBEe+Y6dmkQVa0/r/1LFULg6y7vtJ4o3tSGQht1/ZeKAhJVT8oLTRiKRp8Qe2W
QhTPWhMWEFgpXftFLBMfsGAeww5B9jv6o5jRk7SWcB1msXQUCydFpMTuFFsJawUW
qIcB2nCDNw+DSis9nYYbC23a5Rrq3EuVpusDNzHG9ZnmuvVgMzF++wRryfB2XI6v
X1FZBrBPdp0N3VPbsdOCPJRomlQrhPURqtPxOdMmMIChhGz3irFpP/9BtfWXDFb9
NHJH6no5zsAJmDtPVYwmdd3nfF0f24v8yUXDI7ku+mUHOZPqQmwnv30Q2lIg029i
/17XD7JyFv2ZQkfqgyA3Xs73j6P2jYUxDX+sR9177am9UPl1ihOaGJmSjSZaCf5v
vOAe4FLP804g710ThDps5jyiYhXFPHP4eMob7Ypj8z9s/hX9tpvpKmRoHcqv45iq
zpl+Dl+xk9SXBPg+yJbyR1K4E0ejqz6cvgwC+1Rjmjsg+9fBcHymz8hqY4LCYGyt
MyCLTc25pirI3ZUW8lNhrZxB3o+dnEoU3CEyZgbxl27RMFRh02NQNlogI7HGKqSU
RtuHQS1fG88MCMho6OhCXCIzv8EaTvQPBwNere4bkQCtlpPKIsehj6l/KjAqjQxo
602lhl6v5FccWil9VRBOT8y2C1vMBTxPJNtYQ0yX5tSYLM/HzVEE7Jg9fHR9zgWh
6Wt3Zu46blkzAVfD3Co9HCKejepTs8Mdb8m8xX+V3Hgyp/aCAjYBtxWve6rk6KXO
jGiivXAFh4boFluQ+vfgteouKR6GjS62F6f703zLfIMoECVS0Kv5jO+zXbQOtqcJ
lGu1smGvhB0OsLB3ypcSwO0KV4wvtQWnSGM7NCDpWGlW63nD3L53XQK2WWyg4pg2
6KQHSaeppVJn66cPQOAO0CEDA4Nl4RSLAfDKIKxTpzP6RqAWkU/WqCNoy6vz79dR
MlNQZVi5hdBXQq+GCvUA4QMlGFor6DzMqD1n06lY7oMYBl6dz2jofUw+P58qcDJp
sxd4S7D9UMuJSsuYL6kk8iljl9ci5dKuz8QcznXzeXwV0Q4QVD0CA56X8VBQiaDa
YbSNAnm3vBlgfyd/uuiPX79a73dQeLWOcjw6RNfBa/2skV6WvoWUk0HEa/W2OY/R
J04ReOewxGwH4wt5xt9GyAGIPnH9mhr7/PqWOh/o80XcP3W3cD3l1HB8UVSZSzdJ
fpZK2wdpQ+RnMbbzRuqcQOHzxCHBkltDg/4qIlVS4ZWPhzil2K+QhJJCk41SkW6R
cCgB/sDZqfiQYWX/ldATriEvn2mdD6jNZuIyeKJ1HhE4uaJaXLJBygk00IQvqEfr
Lo2AF1+TCT/Yj2JcKeMC5+Z9E12WtykhBlsxOfKcJxwQ/gQP8mAVg8RYvz7K7Vok
A2oi4DKJV1a5gtemMIU6vHic0DWoMmvq0Z/IEEyNrB4VlwxBymVr+LQTaA6+g6Bc
l/h3H82DPlmrQDO3bYZRCw1Yp24QxCQ56Gf/9IZCVYGoZ82VzngU6WyYchvvzy8A
gPURYwhQ7sgyQv25ltrPiMXafweMCSrb2QS0cZEBzKh1Ont92cDMNZavV0geyPHE
P/r55yOS0dCz0BFwVHau/+aWXhNiQsGbXJGKdfMSNHobEBfhGeWEsQU1wqiU3B9c
DiNbr/x911L6pRNVPTW5y9OaCW3ArSawTCgvF1NjD39VBBo4Bs11mnQzN7qmLk81
bBiGnf5/obbMbtBy5fSLOWjJ/tY98khYP7l+UAIVzKIGJzUgJ1LDMLAxARCBLTSk
M2cj6YqW1YJw1pVWm9Rndaw9O2vmpV3C3CvM+1PXGATBPprt3b9okS4ZG+XYFkB4
vqxSHdt+hMpwjAXj1MoIAm5WG0CaT4UhawZdI7LewsKCgdKP+Zv6b1qHf2Prsn+L
jSFulW+Nz/mFaCeuH1IctOzY2Ub2Qr7mPpJAYaUyAzaRFf5anQykcmy69RD58eWp
AE8Ubp/OxriiKL7KM4ouj+2twn2/3PEzinG/EirHsV5Zpiw36EYm+CAMZGmSuH17
inzRU7smRCMF1R0c46BUu3Ad/PfSQ09G7OQKcnkBJcJ2nHEpbcUCLKNFfBuYVCag
lVx2fpLXAWPin9X5gKwY6YgdCq858ZNnlsrCouADpV9pwBiib2pPXPWVj1H58bIg
Sr39jvIKFoy/fqwrXuyTKAOjS1YHZW/QHf+/tFKuqF9BmYY7H7/TGDGEpv3d7kGg
HpuJGrNi72YN71G6DP06j/4fmAOFa0N7QmVrleJKjY8P0jusIgqVsgbURvtcUhH5
EvaM6FhRHpt8pYEBJy2X+q0YryKeRVaei7g1CodVqZ0hBZWqTgPk+J/ylDNuVjNE
bYJFuMVGqbJL9oQOTs/gWs3dmjUB0/zl9wlw4cs+c08KymNtCH1vQs8oXbu7CHAd
2Ih/FI+4n2Yge/d5EUVlgM/NMuTrdy6IzIU/SPf9RKuLXOiL3RRpBH1bhwRvbJu3
MEVQ31NSsCyk4mGwSC39EuY5f57mo487/Srxx/3WCvP4tMrnRFCCs+UxanEMXoNN
V1m5H+1x1i9W0k2H885swmK0UUgcquteArOB+VX9tpX082YSW0OIqKRK2GocAKqq
l1zzOsEHd7v7ESUCLMJFtTjQDA2a5fC9mzUa7fhImG0l02XCcfsJTS1cLY/hHLSY
C/m3fiELnKZ6XYYVnF+fru1BFfx7s/HkmOhUt5kyxeaIiJiAhC8uA5CRRV7xhU//
LTuDETHAdNZe3Cv9x9twCYNhYaSI5vJsaZjR1/6Y2bNCUcg3GyvMiUdsV8qgbXzt
uB1vLlwmeequAdlUEQBuqIRt3vMGvbhrW4tONrstT8sa+iGRIaNlL7nzTw2E4Sg9
AoZBM4UnQDMQ4vD0HoKTzJ4SR8428fo7SWlKEY6nVXqB51rMNPtP1g8pNdu2fq0s
nIQflNzCiQAwJae6w7oPD8NNUeeFAWwE/NOD/+Qt6JLcF3ZYrNzVnt1u938STOFP
RoQAZF9rl3n6fkW3icWrww2JhrEK1UsKFdWPRic/JL3EyWGVmM/jm+y+qUktU31c
Vx6se3QRmcRvYfgEF7j0dFObzPNj3rY1wlP/uJG4urduHD00JYT4LCl3TqaULsCU
pvlaFHnarrcsr0BvVMrch+b9WofRrmIGBybIE5o0iQ1e3UfZO0sSDTmqqYWkBuTj
m4JRhHhwrk46I6iMFanwbUR0nKHTJgm1s58U6UPTE3OJiRtZyw7VbsrEfT445EGN
CEDwrnyOfIxNQIr4umXORxu1EpaG8HJJ7QhjlVBMR0Sx3FXeHWo5iIT/4a3ZY2vT
k8QPHzTOKVThHBDM1ZLfTyABXcvAzTEXb9MyaYm3FwqES9PZd4MLP5H3k1LF1d3Q
usAZYNltoKN4rpiN5QIZtNQnEN5+HUj2nYgiuz7ZZ719O18aIUY91OH7ztMHR4Nh
ud+dF+8cMVUwdSS5LW/G/wixbbufOnievOlyYDtSyqfH6QfkSh+LPoNfOyVb/FBd
w8byEFtEq4ODU8GP8V5kF5/1Ws95agpuGB6wVqxjxUiKXEy7q/wpywWQZ+PEk9YF
fvKn+alstOlISWD3leffiaANrUJyq3eeKFWzF1sdK2dtMBjP18zsbo7EhM8bTlRA
Gkb2lev24ZZYTRI53xtps4ZSLenzgjReL0y0U61yeynBTScCDsK4hqeFxmilmBbv
YxRv4V7a7UBuD2djz4LuqTjxeihdG35NJ9dDq+I8oTc+uU0FJ0xrQs+WsJMCriLG
3dPC5X99HOMTLgAWULjl1XuCO8+X2fhidR4iR175YRH4/yoR1oT8D85Acof/l4nM
6b21+fHz35SMcz3h/CRqzJLx6VsGhNM+HVwGc526I8su/VtSGvD8gE2bLQAN07Hw
y4+1i4QmYlbDY3mgd4GDK8PChWSCwH2FyF+eHQAo92FcuJ8NwwnFv8vRdzLQSob3
IanG9GdspbBc3O8rz5w/9VNG2fN2XdTdIuTkJ70RYSbYHROH+WdFjBCm7Ym+WhA8
xHrvf/8svWYcUw9zkci4OG+wpnzbPv+G/c6xXGwfgdd9PEY9sHtXjRmzy2WHUndE
jP0RCt8LSz92ZtE0DLoSJ8SoqMT1290EWn3NcDZdg/k7+JirEGicK5AsBts2tfjh
DX+oPgHAIfC3Nn4C7kJafyqS8szWsISc3FlbPsymIK14yoA56+alUKzD1I1hG2Xf
TU4uk5FgDxnGx/J6u0K/euZIVlPTZHoYauzxyHy1PCmJidpABC6cg0ALRy6mr5X9
6+FdtN+EEnnONjluKXo1zfNW9ESG7cHMkqXF4AI5zJHs+ax7CwJih8AzDv7IDBP9
+SYk9iZWA/IsRoHQE50vzk/64lv0G008PWjEZqGW315lCFne0MDZWozV10K/jhEe
uUwIytXcmXK9C+VID0X77IDRjFsL4mJb4VmPD2pFLlyq2GT9ieE+WLb3cMCwRRa6
+PjfbokEkBV1vS4fL3qmLpIY1BqRzL2ciugKR8HN5ObX1AtZSzvQr/EMyYxUmTZ6
LZE0khOjl/K1XPs9bSOlMpbJVEBvjP9vlPlIzQXx205plptF2rcyX4neqKN9uOZF
bfuyGbrRt+tI8dhl77XfKVtBpctJiu05TYeSS+5YyzTocaLrDfC/5ORc5fGQqwkw
6aT7b7nrIR9SQ5mYW/UEdXggnKfmMviFv7nWyIYeHztCX2B6O0Vdv0EqsANJcyMc
osZCdSHIQhUQgas6vfXylvUIBMUpqdWaGVrSMQ+dM8d1EWAqpsHHyXBWvJ83N0Le
QRIJJatXuyVM6JluBB31J8QMa55hEhyCCeU9lyJXtrbU/9GG1ZaMq5i5iwe7fBqt
0zNg0uSTxb0VF3dduGQIshBLxVa+SvW9j9QCOAAtGmEoWTz/J/lYF+t5mS4gM0Yv
m3Y21pMFW2LUgpztmfTjrdGs26AQcIWGv1C8iv/psNFCWi3JUMYXQsMZi9cibIbR
rsLgfJ20mWBB29JCZUWeFfl27hseDx8AnoH2OHB7VOurDwpo0YL4LjKE80hBue85
ZOWY+ICQb5nV545aHQBdOqo88nevZflXU5u99DHVWxDSAaZmQwejzWrEx0ccZHfz
osuy9b519kc9VmPTox8UfnNjxDX7vO10bHKerRmMoFseXls1lLKwgii6CmEou6Vs
YMVUyZEmV8csBIgj7aw4qsIa+w7EpDx4Q8Z5AcWfi/uLS7Oj2pjtSjSYOOBL1WFe
88dAk78f5oswQ0kbwoar7HFiiNj7daVEgHqpyBE8E0pke4aX+LFe9IS2rGIt9m47
NVsQl1YmKcpTy4xJmaAozbem8e0H2VJ6Yi0PCbYUjOGej47dDtzN8JTx7WVv2pQR
TYWYi8xI/AjCmtn94mEJ2CQ5KusoMmpjXkfkf4S9LkIYtkiBbvDXuugn/Mnw1uBn
B2dMaXJpH/l1fxUDU8gV5dla4qpM1AIcpscwB5bG/pJqzIdMROLs0s5iPE3E+Q4A
CXPNbvJWh/UEeF2BtIyCZBvdVfqhBMDxebcEIb/1AVNN93Gr5+PCmZfMAMcf66nu
vhT8KLYVXKCG1tHemMX4A1yFzgUCsD73nlBn7vnI7bnUGvFs7YztSdTS9p5MsGiu
MTPrafa1qggDqgfTIvgcbGY2ri9ZUl9WQKtecoO2D8DlXlt+8HOQR7C7vECSibwF
jy3oxndTYBXjGm9nERIn00m1k2dSytuCwBguX6Lxq+G+nELmlOPjbnzI2PzQa1d4
356yX2rZEK8g22qMKJi1EKW/HLDEuGILHyrHYWgIheMX22COL6q8dVRi9wFQx4Zp
76j99tdfY0MqgzgcvziB5wVoASw8TsOI8T7vhWZ3gN5/Vj/vratP/8pxFSaoJbgj
ZBohOeUtjdFjmiINpWUbc5CnrkwaE5Sm0mBNDHtMyhb9DE3Tf5Jm1NmR/6HoI/mQ
dkQGYtImMlA7eLoma5a9WKrFVNpyI4XBq8P4n9dCn+N9/29hbTGtLuVjtuSAj1r2
lC0mPQuwA1e/6NTyvFUqYtlu8ChMOGaqbNukWbJHzN4JDycL5pMlHK3lnzy7Mc/x
RCCFVwU5fkIUxA8NEbTlGgLjNs6gHBR9pLbZmrgVwsNFfKsJ8gU9EtONRxD93jhd
FBpC83aiVczPc8g8N+GsoSjXdojrCI5jtamgL2yPxGYcXWuswlKvp++aegS9veqX
bea+vfGEcPuFkdFcD3k+EiCXCdwoaUMPRJzFO44NOjc2nVLkt3un8xMf26gX66Y7
6RX/57goeeyH438qe+C0O0ud0NP/ErRUhzAG4dbUgSI9KBvLx9KDYxqaXDKjPiCi
JsH2+/kq44vU1cpt3pYAVTsF9i0Zp8gsBbMyFUxbiNW/jV1yrGQnxqbTU/qKy7HK
SYAyhidFDFe+lBQbwHokyx2HheO7zUU7ooOmwbU6/neKARyuTx2MM3ZRi4VRKprW
Lf3kdf23bat6b5Gs4lJw7yxBueymY4ycP+W+Z6XPwrwX87Mv/SRnyAmKV8zEPzx1
J66egtr2XY+yll5Zn3yGxCYqDMvfm2SQLMR1CdZPEAJzPWh7v3Z0s1CRQ6jGBGJt
vtvL9yZ6rn2k+hejTfo77s87LlinhBPbvovDn15w2ssOZjh6h0922EwoQxrgdKfF
Ersi+SUjDMY8LO31uC581JIPy01Z8jXhosdNAp0AHM3920aDmbjvqiPt3Dd+q9JD
YQkf9prb6OfOJBukfT7PHvhDJ7ruOjtQoUZelb3piVenakTAZpgqtiIB7AsmAuzS
OUyqR2MuiBUY+ztdaKTyO6ENR9M635yExJEvUF7foPhZ4Pw6VeFxx8Tv7EyAgIf5
D+g3K9kiC80uouWTxjCUMpKLi7gDgjeK/+CUyFYwydubxB3Wy6GSrkb2sDEzhawR
rpNA5j3KGAStyKSoyVeyUvo0j0ke/FKSxA9pPpWpK14PgxZ5TY6MvFBeu0oLDprB
W7zQtfC6K6APYFwu4+uaMxf+99wbd9g+/aPnhZH9Und6LGl7Jh71/CUh0wKcKUuG
b+3M4UiVlfn7tYIIVL48y7pos2YorF+wurKXNtvZYKIAGT40GtGjtqPdvF4bjPKI
jCFPODWw7Wb1ATbP5Z+UNdhivxECH445DQl/UP9T85+bf2RzD93mpa2HrqpPhF5w
yRJ37KG5s0aM5Q2TXbjBe4a1jCd+kZVFWKhonxDptaJOryjfeheKUA1mP1LuxNIU
wXXJ7s+jkJ+4NJrG9KKsngfNFNKEMWFoi5WHvLFvYTYuZ1siJzzGynyIjlHSaIzV
2QZMQt1Wh/qv2YSrE02vd/Zbdc9H1PT7mqF331/uLNV2klUPwDAwpsjzCeKWb2Cz
06KBzjtNdGb2gdV0u79knO0cEhn3GH/65P0odeh7p9AioPHearnc/CdoLYM4lR4g
MAkyCAqxInoR0AwRPZUsC1D2MBMKCZ/VeUB4EcEyY17N7VefdsuXLkbUpmpLfhIi
yZfMQb189ixE4jfdzhJlrpKFnZb3N+zF6/L6gDW3Y1gu2hpK+kM6v1H5sI1ehQ4V
mp4gvlFMGn4CG5/TgGpmumtOzY0KEg/QJH5Ou4Jli6M7ArJj7HAvIX9ivlwALAjg
PKGcXxOZmkuKAkiNxQvwBAEpFJmw4Io+0iBwMJBrLpRAWuwwk7jBleedqmUnNkRA
VixmLTelfDtUE1L7BHHFoUkQvInOxKzBVhOhXIwDIXehZbHWU7COqbegUMPa8Qb8
VqPsWNsCMU3JsXVECqS0NjmqWuigl3OCWktKLLt+xKVu/v4kngBTio58gsHochFE
JAYdp5z6xWimrKfw0skhBCguEpEmD3bn162b7tQZukjlzwBxhb0kM2GlL+8Gx79P
yYocjX4xy/BK3hKKEybJG9uxu1qw8qjmDnphocsaJtwCf1TLMKZlrdxgmRP0Tw+A
4tjazfQ5SOzNk6bDdcRDdkqV77FCyBbBdKkfqd8ADBfNEtHrm2O8TAFbO5ryPVZV
UZhMwAgoFHBxQPe1MZtCqa/h++3aOxNBuQvoQJ/UWx2iMZY3PM/da47u5ZmarrFm
LfRa96fLRUJjG5ki3IND2GZrGhZ3dknCHnEn0tpVnfqYPp31whBwpIlZD2P9jsKE
g87ckX8SY3hYsF7xHhBIu9U6B88Pkv3uys/SGyM5w6wmTGpkbMUTNdMv8jhM4Fbz
qlQYRYoHW5cvaELhCsdYuf7RZaECFFdYWsPZZG61Z7bnpt0nqmFdtNYPf7wJzdSV
4Ghj65m74hst5RtzgkL30SpVXCCiNObZC0w+tRcWnwHSblQ7c9RPoh79Hirl7CAU
y1LM8pagtileEyEpsgQKdiZ1q02yfKiLbhAxn4UFvj/fBB/yIYJn6+sEJsBYchNz
KQ63QV+joA3XFs3yxAv21yQFYVY2lLF/9oqnMUTnXSqLBOSio+IeC7ZGaXnpwTC/
3cQjF+bBRCol3V/q7JAX2VD3vd8Z1WFgM+l/506vNUjhZB7/BkJfq9r6gSwZpJ+F
TyT8La70nctj/pwxfRuF0o7Kd3dVE86kgE3CU7HuJbUSmVXKL1wvUUE4AZHXSbyA
0etBZGNbOfkYMgkZr+PvLzmDfQjGSuFXxCOonDwqGFhNu9nIm9yki5vF4qmxUXiP
lbiEnLjA68xyuFmtOMbptx088hi6YFoCTHOqXPtivY7H5uVtMvLehJ2lvNSq+Avx
nreJRZ4lwoPavfs6/qaGnkswj8qfmzuwMTGMh/5mkEIpRwWs9f2jgDj887wyFyV0
1nWU1dVoiL2xNWJ60pbr9xGCH2XoDQ3YeCD/GAb4Tq+ukXp7R5xpV8CrXch9v6Ne
xyDIVY6Vo++JDK4YGMMNGa0vM/V7vbQILtP2M5Fpo+RFbRacREYGLiJB7Psmzm90
k8PtYQ//KKnyhXJc4423YkXMkalXBvXMs/l0KWqqatBeyrcTmQB0636jsgKbWbzf
rk5m0JF0uAoFvLyWR5G6OZ7stSQgDgp0wL+yv7o+f7NP9FteUg2J24sxBhoduuIL
6tAK7ca59XD/RwDRz91XQi39r99DIVUhn1B1hnLQniDjPDL56iO8sngv3FMYZRrJ
gT8mzTsg0CQP16qzCJ38yKORiDEb0jcptjfjUOkZHp9lNMb+sNHWD4T8RulwCH0s
XwI55xqWERMWjVWD0JElw69smxRNcPyPbCkTDPdhdpqBKa0jFO684Ic2AYv0RBf2
OChoe+aaL2obh/ZGmmPAVjxqUwGQfHr3TBF99spCZBr/r0DkpILV7fbgOye3yGaC
j0ln8l90Bvn9bYeJG7XiUNLnJ1YxKHamieIfhkwIFFKAsAtmtvRthAVY7qxVaLvT
AZQCwJQDYUPzU/6suOT9SkEi+sqotreGuoMV6Xo0jasfU7JsvbDcTy9Bna31I+Gq
f2UJNohcmQG/KmnKi8fqJrAWe2j7WgL25w3Ur1CnbUAvfdRMhQf+fYNaBXaZBYgW
U/JL1hpiuyHWGFNpJEtgBN7SsapoQtpxAwxfwQ0xgS8dFomg9iLog3Sbquy3SZgh
a5SfhECeu3pPsrdzja8xlnYjfZog77q6IkFSy9K6VnBr6lCpkj38Qo2iUgEKSvRJ
DXeNrkhbz4Lk7Va52imTENadXm4A/nPES3g3AC4/YpSIiHMr9ff6J0k9N09EZ5pu
uinnC8y3pSXpaE5gMzMjKiUFyy0Mc67e/JH6g2NzBNtVhas1Qgp6E3nuyfPlvjKD
y8a1MFc8M/F4/jjn2utpk5mxNN41ymfezJ1Y409ODh0IATwXwlmqYAieU1+jfxBz
AdSzTvsICgM2sihvQ16RrH20ZBqKID4DFtYUzEXD8skDmG+EYJfptNyy0cFt9PqB
VpHUZKCVg5C7HiQqewRhHGgixljkCY/9piWzgQn+XluCr59HbzPYXXqbQCaPa01n
H730ARKoPE1Zk+ZdSShfYwfLsoumYIXZAYcz6QVBP9LxJvuWAUtdjPj5nOHuuZbc
2L5wURGneXDXdZU41cmkI+3R8TNI97BL/AxZDYYnJ9DM6QZQ5ptcrrrHzFFns7WT
rY9pGEaN+w11YLec+sZdOot7r+4+yriG6TEKG8dZhb5o1bPMbY1cRRXgj60MLRUt
eZ+t4rxEnyx1LZF+u1t/ZJltoULLyn4ahNin1d1tdOadE3Ma57P8t7NjJ2E7GR87
P+rTAwFOvCIKbb5FXkw3M1Cu/jw6RTHlqST1QCC0i7Qv6Z2w5aZrPS4vWbAUowSn
Q54HdvLw9n+0g3qDIaX1tUa71mQ6hvEAvULfUpw2xcMgaMX6qIXowi/BMAKr389v
qrScGGmseB4/kbU9gS3hV096AfGu/V1T5+PczMuA9VLWU6zVSy7EdzYfHLwMsN3t
Dydcjz5N6Je2fcp6BmGsRTUFUa/tb6ejkvMzzltc+3mtK5SpCMQq0DNbvFJwPibg
EghjMqnqLLmbbqGBpHJTw+ktKuaeK6yl+XQ8gmMMKrzn+rSB9nkHBffItCZ8GCQH
lUEhyU2MDM6GEMP0ar7ahPlc+4E31ioFPxHp9lbFdJroQXoi9Ie91MtQAWMwJTU4
ldDc8M9V6HMWpNfKcQBx8MJRH7pYQtHalvFMr24AAa8GEio73OXhMW1/sNNK4n0x
Azib3kowj+ge6PS3fLZ5jaGompah+d5ak8Mvy3ItN/eBbgD1Fwd6GGPQsSb3mwme
XMHEbbzm6pA/J8q190+HYk+DEziO/icOi+c6gS3nxCl7FJHVt28KFC2neaA2P+Is
SfaWnsd9ST6Vyub/K+VDfs4VTaXkVOnVbrmjAiXuDqQd9qqS6vsHfdVXlc3JRBXo
F+qZTsdQF8+wG+v837gR3+izpJY+VZLIO8yNaCbK+Ytxbf2sJUtqmlUAjriNbzLY
OVJFUAgRN52x1BqEH86G6h2n94uSh88xh2IIIQwCgW1v8kLtEHpmnqTVbU4KpOgr
kRIe3Fg9gNMDDcCdMAwbcukoA2TBLFKCW9ZJJFJ5xrTzBtWq/2eBeAXw5Rl7QEP2
qpyOEKsn8tI6mjCLNDkSphth6y7MxefFU+61CQB1ZqwicltF0ex8BK59UnSrvKlC
YZz3ou4sf7rnZ253VL67cW/gJCVzFKwKc9Pcx01UQkgPwja7pVcYGZ3Bv2mXXNYE
x0v8AG3voF6HSCTMAAe8gpoany+U3DYaj6efCScCFCJ1qvxbkmDhgLJ0iykY4l94
k9e67jkbepj95YOqV27Gg109v9+x5J9pidhi3Y0TfIovZyAVVCA11Its+cXXjpLR
Ud3erunUOrCahl4NCGRP7hW80PB7+Ea9UOKUAFwWlsUsUTaip7qv5KYT8y974SW/
kW28RPPV8Fwd7xAr8fheVsPWchUwJYt8tjWhQzi9ui/NK9WQjSNjPQfEJe5dNwzw
lcE9ZNmE42oeBGJRT3ucs0Np6Q74V/k3EpiYy/8Lf+rCdV1eTf/cG4FYGy/7oihx
NCfV/bW7a2/NxOW2lvjPUeJGzLrm7bJZUi7YyB/RVEGonGKDeZ87EocKRQwKUCxw
nJe/xOpwjub/BcqOXEHAhecXgNhbNQaPANIOu/N7HZLW6hxEyxT1557x0fnU7o+H
cXBRRib0e90oRKwycYZI8fQLfWLrfkEDgNqmAsc6/NncqqDuu7xiMDC2ERFgYT0a
IvrsXBxbXGQ5ANC4YutrxudNT2iCKyK0subLTT1i3CxaMo4xltY+DUFqTbY8/6ei
DloYFS1rElo+zlxTSd4sB/y/kZsnL2KMXIb5DsXaeR2yRyV+kUgXI/HweGD0Ee92
zU4jcq0/95fqBeRsmcpq3qJRLoUfJ+C4My2qcgD0B8gAl32niqK/C0NSBg4u6nME
K2fzutW1S/IsXn2D3kDx3uVVibEzp5Sq/ZGueS3C27nmuPkNN0wT1gAJ4ia2w5EP
1Y+VOEe4vdXfegQVTfPDfXClgGV5MaAX5qWExd0VXXYd+X66OtCKUlk4/poO2Zmz
RewqQTdLrXPVx+T6NmOKh4ZfAVMex1i0tl8/KZq3XIFj2SwoP3q2i0QDCPkh13cw
5Djnue3bWnG1QqCUMzgW7iqHFmuicNuCh7UPERHePu1N5MzpxiuCCmAZkcf/PkqY
JxQgx1p1UNRgbl0L4uH/sJEVV7z/T1t+Ccf0XbBb+oImZEMj2Ovs/IwS7pAKymes
Pd8Qg23vj+M9VpbYj2zq2UEzud9GrmQpM4g+z2tNj7AeF6DAOl0sqFhS9bvk9s9r
vQ2sIA6rxoZHubQ6PorizUx0z9eLduZaTOIJ/eWM7wnHPLfDM107ps8j7bjJeeNK
tHG1AkKQ6nm2N34+SIz+qE/s4u2ABd1LSDpsgaWxWMt+idYlBSdHUm3OZHPf7SO4
yqMCjzrguJCjvKDFMsdAsup3kcHsSJbLOM0+Hr+P0LPErq7vUCL4r8TUojCpNh4Z
ngg+XmHNNzsfAWm16BXkeCFTOyGVV5yPjz3qMTyU3tmw3cYr/EhfE+B9La+JtBLQ
WGuxrvW476nnXT7eGJ7ZBR+QhIJ/fu9ZDszKY7iuOlyhl5BCZcZQnDope+w0Po8i
wwru1EbicHEqdEx6cvPwXuhpYo6bspJKyd0fTurzmMXrNhB84qZtPl5AXGqff7fV
0x3V8xQoVDQasd7BJ84/XP7IhuLm0OcT0Q/h1mS92z77o1zh88CUr55jgGEWGXIC
V6XF4XTN+2iJ5IF3cuW/6ci3/tLiFjO/9NpVTxllbSChqeFSFo7dpfeND+yjSJ+3
Hb98b6Ef6YxpzSgRCsd0GNdrKgZ3Ab3ZcJ+5nYWK7XbtfY4lwF/NMF/rHPKe3jv6
Muei+tD1ndOsIhJO9UD6EP2j+5HrntO+xqAljdhFiIe5hG9BefzDwnJUGG4lLuUw
HigI8MJgbsDK2uNdlxkapGu6J9jx8qNbHIOx5ebGhsIvC2+Okwc+Q+yV+hzqLqej
szP09j0JNmn555G1k1plpv50CrTlro3Uo9OTslgtbwGHpGhXvWr1G9O1jbqkt8Pw
+q9CbTxz4NnFvvnV3oXB1G4Gcvh+Zow8ToEr7rxDsu/NmVTv61kQ82Ne0oqzb9aL
Q4KOQfiKDnDFW8QplzL7a/TGOnnBkQkZ8zihGVV84t8GQgRZjWIUzcfaBcQ1LexS
yCDcPueYRsu+5xlc67fmjF7/h3vbIX7RPFSegxddV/LsgLVOtDEWxky4KNNnO3mh
ksIeu1Yl3mfPpA+KrUQ/hq3Qr1gZ7prmk45ttCVq1jCwAym8/CHzPxYe88KozzRL
p/VMyeUuZmCc27VQzF4KbhwDEKmIbY6cEtieT5hLhVzyuvOdqlE085VoCRqvGZ4b
UZ4YCxdiHb3lcms3Hzovae+q/cTdzaxJCQyZLCv2fuTWmxoj46UK1DPB0fsYrDgU
DAaVsdQfvNYTPpn2T53zGhOJjgpz1YvtZt6UOHOoq7Xb395ZISgIvAylleuaK8NZ
Uqs1KCCgtvD8M/5E+JBK7TiGa22VPxYbnZKoqfOsquyCPFS0z2vgYHxw4lMxmBlS
sT5Ep/Vt2KDrgDK44fdle3X5ZlRdWXbmTGAKvvYEiJAV25iJ4WNnRutqhGoyFTpV
9IEFAKVKoAoF3Qiad+MEC5mQSUWCHCoLjj6vaVvz89E7eqUDwYNwMNwa8lKshQEQ
fqzVnimy/1ySvZ40nORRqzrRgP/6VZP+dM1VkDuNZpSbgjC01m1ArliaUnlfV6w9
WpLPaDSSMJAID6guISb/I6XYgbWuJuSUQSaXPEgc/kmkBchej0jMYahGneiOewTy
E4IAO+w76Q0VqxMT8rOCxZ1RPiyRkmU4uSRTP5iPpkweCW6andzlO3e9oxs03yS2
piIkOLPh2fkGdLMT57X7M2vFSchyuFG38rASnG0jZpo/z5/LYrSLJE6R14+yURaG
HHSVcJjctlyRVZI/ZdC1gtfbrsZD2n5MdfCVbmw45jGbAZNIa25oiNbYfvKTfhB6
+snsxiuldRAxtRjZsCWB5sBlcwtIc0uOoWtSBHg0Xdu9Ns9J0O6/XzyZoNxI3CWG
b11edmYA9Jvnsbd0QEeZ9OKYpNCJmrPsdS07dT3pnH32EUbJdJgT4ZfM+cFR1XJe
VBxxsWUFQuXb3BCzsekETwGdmWY39y+WFdYO9pwakA1Gi8BnpSMWsXLdek6zWfPl
Jo7pogZfI5rpbVv5cRvFjshL3z/qzdlqSYX713mQQvAGjuo+i9GNGTzWFcB9v2Tq
pQKfaaNNIk/QRIYJ/SbSrjZdWuwkKnfajhHVJNpM5P9waNQiaVyD5eqcLA7199A6
PzKiNumYbBPmCtp2mObJtHOmBxbWm5hxgENZPDzlrdeQISwf4a2noVEOH0lO2FP8
PpTIMp9PHlPJrGV7RNeoJkzPTbl1R105ptbL+/1lZbsKmO19Ic3dE02WY2UQR0ws
ePXJG5GTxzT180juSNDGd0uvSv2xsaExpZiIurw3F7LbSvnClY6nAuTRDUt/DJGP
tcAsLgoT5qIVyq+JQgDjIDnRu45PZld3j5CQXgFy9jI61b1Np5hl3zrYAN8gBBJQ
iUeSIzmONOm8R5f2piYnTLx9YwMr/o6aYGytovnCdxdY4PHacJ23TptExefmSref
ais5bMYl1EXsZRDYqeO9AF8iXJ1mwGf3bj4KO0mE1ZpSMoWUjNTih2/bsN/b6ULk
pS8QGczAp+DoHuMX7Gs/wIpC+lSMO1vZxcxspLhySSP4QITj/2+90ifaH6bSA1QA
cfrVq0Qtwx5Ps3Bf4l0FveJfkNUHMA9VLQvmIYXxIc0HJC7HmjF8watTs/zF+FP0
Viq5Jwznb2WrWooL9ml4SX5g5vvllxUkqGEeu8p1ADNEmwUseTvtoUG6xPsLD/vR
xfvcBLq6TkI0ZrhUnKjBpiMK5co1nZf7TlJ2gD/l1gNR7iL6hVlskiTnk1SaH5Md
sMNsDnKNeTGVDRO8U3Qu0VQqbhoydkUf88DKgedYNDd+8K1K1HKVVEAxckcpE0Sp
pDGmV7K8ppUBbSiBQi2LxSU2ZoMF4yGRn3eqCzMMv9TkWY2WMq6LaWGWedvCBNOR
/Ay9h3cnMdemhP88442gjscebnhscOJfXlTD3z4FIdKwiZL+piXPyYCHTA4L5gfK
CImIvS6Wf/12OsTFg+HbYzzDbJ/fQzPfTwH5fkaZ9hs2PXBRZdO2w2OlzWxKkWLw
mv856e+h6f2CoRqnjGU7RMK73D9TO3QsqZzQx2YaU1JHK3cbYn/OvaBV0Bb3LqQt
OOphWPPa48khpaC3EyQDKN2sdN3R7hFZtjmTR4pEbEGdpVrcCfc0pDD8at8Q+8rN
1qkOnA4WwtttbSHcgqErvwZnNcSEOrSldeI6+AXbPd7wyurLjwR07csTiTy7Ndp2
Iib4iP1Rr400DUbngnGWe6ByVd8gB9JHxndPMjizRb/sTYl4IwaLoa65JFKpAfsy
l1p6vB2nQ9R35VajRVm3fRSQrT0Tq7jHxWQnYg45JwxjuW21t+gAIjSgIr6WbPBV
qKc95YZqRqQv7c4ndX6ACgtO7JSQX+M9nnzqo4qPe6CjIaRqBSpBnYqv4a7Myopo
m2J86dQX+uvwUpfL9flIRBtHkcGKhByNTXfOpsSRyxbpAn3mO0HfSpQYvOSzNVNH
6OL0pUlEBp7Dd3yZUFfzzAcvThp0DglVfuNr2xHZ4Q4z/e/wN88URlrp4HGpTv7h
ZdiuQmo1lM4MtolXjzGpU4lRSYCuYSbTCob6/WCUddBTxqqdUFwUohemI/UXyZ8F
iAhKSzLFcqj7418xnJFgtEBxWfTSJBewZtMY3FfpXKZBasiA27hO1ZyHc3z6bdsu
WNiQdOvTiNTVrx2Po9pGcrnytB7p7R5OOY/yMD3GMcGbB4aMYLTDrNnaaM/aJJtQ
vDEk6cFxWhNDKe47ChYCZVksvNaCaOhNFuOprxIAmTYfA8C53VeaKcaV/EWP3Kqr
P5kP76JfpcMh7xvGl+HLGgoT+T03UgLsvYS17FP0C5fIcORYVkZXsr2SlMMcR6D0
zQmJONvvCa7sjkGBd6lM4MyuGSKyJOibzcUErBEha1eB0RGkoiFuI8+9IHsboc4x
So8ejqBgc7h+WXgTzz12bzEKxk7m6TjbWJeazg2GydLg1EYg6G51n1j8ao45IF/N
ggylCn5S7jjvgpJ1qnOvn1daj19E9sFY/v22Px9gfzo7M/OY0TnWWtA8eEMQRxxQ
nwU0tMNipmaImdyaXmXatXcOpZ5SIyOMfoNSgi+OenrrxAQRY3+pmvUt8vHyhQu+
Q3RSWbpj/p30bRRQsOYIMkL40qrOGRfd25hAVqBi8fOO/WvBzuDbB72jjCYIl0jf
k+kTwhbwJLFlDOabbwFKUz+2I106mgFaAroNTlZgpkH7O49SWcJhKuF5Tqgn6yhd
otLfZwhhClJQJwzjZM2Ovl0VM06bprfU7rvOtFgzVikYva/KAtXbE9vWQpDsaFJs
AR0i6ISWXXv3S6Mgz6sDM1wJdf0nuQle9zvPihnF/qby0NxKgqgD2dsMmZfAGk07
GBVNKiZH8EJinYDLaC6hdrqhaUYdktiD35T1ZGEtWFoQV7pjiLq7NtY0HiACtLsN
1U+Ufsz1PMu8O371dEmYJmEBcaPtnpxpDfy/7ov7NaSNliUlEMwO9QhJBUlvWhGq
yMpEaaWZwDteLZfflgb3ihMNFvcTK958bxthFWLXLGnpdN3xh1ZOtkUs5BpcZSJc
Du92lI6xLtVqS5LvstQdKykSnJcjMLFlQRU+Xf3uQBBtBq1G8JIBKgT7aBegiV9E
+HXT/asCQIW4N03XHlvz+IIpIAKGL5KGCKFgSHmhMvfaMtmw9cEnCmPDBVbmzEPb
TRWINKqMlAQ6wYVCjegInwBjKAA9aHCJcf5I5IgP8fK6uNDrYDFfYKQ+ziFw/l42
aeCEE3qbgfEgKlTumLKYAXtQCoOlnvgL685RjuIWFMZDanZtNBjY46cDOiFLage/
MjOFrLEApjmT1q+B5bfU/2wJxUArNMlTjuF/BBIO/+CQOGkv5p2BGSy19fcgjl1V
wBis45hcXbGetCocXREnwsq5ljxY8J4h0nE/ahIrbpsYF1RzbvMDsh5gDbi9Gu3B
pr0b8Xf5O6iJJCgZvgesdSR3RbRHkcl89aF6Qe9IsrFYG/LTW27rBDzo8cEgqvpm
0Cu4otYv2BlCqS8cJrdQMD8AYbGTBzmCewX2sQ9OwA5YWgPgNxOR/GfUBw5R1VNo
suJv8X+FDqv6DhFJbk687aaUuTaovPsB5c483ufV8qjfl60IPUL1Bo4pM1aLseyA
wxMNxAOnMOZ6z5qiX7tTZ4UmWn2bdIFrjhiKymndDxApaK7p/GAg9qxV/pyTMLYV
YK8j0qKy9JD96Cvw1PizH53FWfGYxeU7HZF3x+NmwEHK7IIg+2/FIcC2QAjngAa0
2jrs6rgWhmNO2tgM5wNnfHxfv2YfSrikYlcWkwL0ws45FN2RCXeAdFqUkQbS9F/O
P/jAQaI7XaXw4yT1yg1R9+g7u7HJsAPOULsWunagi/6vokSk0JiAYLAkz5Ls+xMZ
8IBic4e1s6ORsb4NIlk5ZwbXhY+NRkdxnU14Y/H3mOCJHA1NJqMq95ARYjSRJ8TI
uXjzaUvEQKilsDf268Ro60UhT90MVp2dHOUc2Qg6E2rkYO+5NAskI2jiQaDrI/Sr
sZPMHhUmkA3o55RerBMhHq6SlEqQQ2bkCZjaEBjqVMJVKleCQXm8jVND0aufcX8l
vSWIdf7bklzVtU6CgyQsLa+FRut3WJp3qyOn961IxIvyx+qvIyc1a1pTWo+Xy8dH
hHsSnuODfXkhrJLPXawXLeoPPuFhLQxz3emnMQhQtiT6hTmdCvFmWS7fcqjj8zQa
l/g8rw3I0TS96UjorCRrxxtO2LDQ6wURv3a2secZbabe/XDD4zpDFZuLbmpcab2c
uHvTBqjFpvYcOcYJaNgwcd+wOEiVcmBVNGgOas0lvjQOn8TUR88XhIaK2w8ncwv9
qyCxqwK3MUUILgvaL3jvp7q4w+eRtgChQavyshCGHA5KSV2gEgSCjuHjG2nT2KDs
UsjmG+3jtNepLyuBoyIolTYO8ljL7mI+KZrxVuzZLSEJva2hPOjB7Yu+68yd181A
MQgPVreVvH41A5nzNwmStvslmt1Z2Qs1x51QEmKX/KquTwP67GgRLPjFBkdtrc9J
KDekN6oWAock9rq/BhPHJdQCEKLOtwHTIV5u+4W9ujh7jPgt+kinc5ypp+Y8g+UV
kKgha4HZ8JDfcptQOcTr3tZaO6P2KC8nRmQDPAl2x+SSeuFuw1wuifIkdXGlaLCM
f2bfpRDNW5VTnu9J09cPOmgeQiw3PPLj9s08QlVWfltxw7O23UjRBmfl471avV5Y
opwyhL3oxACg46VKR9hkS19x+AzPHNxwbu+8iHfLMXBZsHrnfBOillPrfFf5cTbn
5ku3bRSaS7kk+oH40HFjovltQHKQaMIDz5L3FlE5PRg5IjDQUY7v1VgSuIG0qLvF
fychDCwZFKTBDCTfiQPYLMl7W7NfdnxEIxwmWg2LVTZbACkfTCAaynGEJA1SQmHu
aWFOOVXfu/1LmyIAAUlsrQTPl0HLinVP4chGGozMwJhMf7qvBCB5Hx7jBksEijDN
XzHlrRCSfBZrYZGPUfd2vCkwlyXQZcfsnhZOkpuKNp1Kecr8rFLDYXeFED9coU45
TcnVERBqj+j9LnIDZdaWnJ/KUn6Z2hZRk90xUvC8xc3wprxLXrOQcySyBUWqBeq2
tHJ37QkdJ9fCiakcQwL/oMCLEBkY0J5xS8xjl++pj0vGXdKeqzIfoEkyDYb9WGBd
w3GsPjfXkZ2WJzIbrEVjV7nUdqR3PMswouXowBvAgOHOjN5HGOkafLqHV5m5rmC5
8OiiEIRIzdRcVGk0maiJ/6KHbTw5oR0fTGXk8JV7viGXUy7w3mCE17KwmtoMWFTk
6PHC8kK6rtYBwxUfdwTLU69mcXsQ7geaFIE7TCHcjYhyopxak8ukbWQuNzB9KuNi
Eb0/D0uTNweQPwIKROtPuFRSjr6N0uoMRUkohIera8Ujhx2g9TBxcXrzRhALsZBb
CrF6k1lMVDvR4QxTbb1I80hybcuRuH8frri2LzRh7RU5C4jr+cSvT8hZ7+Z35su1
W/rIdjPEzXhNERZyL0vrRm09FyI+dtk2PqXaNlI+Fm41MWaLgQtOBLSiguHrtwi3
1fVyy0EsaSJTQRD1wa1v2jTTwS9EAVeJj2EVEXCzs1vlCwhOeLSv8591t5GHgpSP
UF2mrp4a3W4zpFBAOClEKrxtmeLEjOA4DmHvg98LRi6h+G16oPsEYvih3xjlmCAF
oA8lCBhbhZBmzunyn9q8cWi04FF/6BD9NY0BV0ksGOPZhxv9ixiaFpT/zjQD5O2N
QHkmohEekTZqJpu1UO9T5Wm+zOVyjqRx9D1o8LzGeeqiBVRDfT6nXLORShYbEj3+
tILzYlPbedCazsl8ATpHfhC8zRelTlP4DYUnAdId/zb1LJ9EMKEWZmVu1n8HdxE+
Ufx5/wuwdcj15U8I0ElbQmzeWEQVnoa1z5K7Zp2MVXTDo0gZLi1nBnR9Im/RIbuA
IbVvZhDYTpnAszJWB3oy6MfPhCoWORx/Q2FdT3U6ypZp3jVNkFODMMV4OTrXNYjb
2291xHv2qvoFIb7hVlDOyg/vH1iw3JbYDrmfLasX0MAEU/M/kMe7Ktla6x+JjWHI
AwiypqI8oQiZ5v5Y1P4+jIaWMh0YU5Sg85Ksnd6VRFjZY/7LbU2wffyN9gygKRDv
2hRQywBXKGeDhsOLmJvETahcEnR2oy2YG4r/yS5q5EdFHyjcvguSlC4MSeqTJjjB
l/V96mXFK+rgQFdZwH+368aEfqDlguDmzcPI1exMzjv/e2RIkTZ60KQoewznGD59
DDvH4jeLB6KQPPj8rO7xfWX4gWBTqXJ9K2AQtuECQMShUu+jeLKeXNxI48+s7b0V
j1jP+ZfUx7VD5r1khpNKJU6x76MI3Y1MJ/xh7hyf5auqc6I1FwXAJ2J6pHJlXOKG
0o0sdzUzw5eQVjTiVU8spgc+zFDyLrdy0MI8aPbX3Wivu9637v5cNL6pmlatclGB
Ovugiulh4UCvNUaTi6dbZ/XY7S5qAT8Y+E1OWazvnArE0O0q84DmyvUC/0asZnGH
2SIMQMn0I9BRaKYiL/UPEOXV707AG3jVtjRSEhR0i1TL81qMnTU5z6uvbVOtwaJQ
gElVSI1+MYc3kxOqo4kiGw9Q5A5mMfNkyG7i4j7eSZC2NxOXdAB2vHg07qrkru6o
scthRMun7mkdX9qdm5Pupi1bnwrvrhDCd1xbHW9CYDT81RKbp56qDaWRd+YmQMXq
eM4ViLglEmfVZNL9usguBID23e+cKV52Z6vTMySlUgjreFB1mTCDz+7DESDo6vMe
Mwl/65MySqJc5txIcl5lXUrCg2whqF18yRAOSu7v3EUHdeAk7xi0mvbAk9Pf6KWU
1n5BnS1tKoQfXnIrxeLAMC9iQDOuupvTdIwHa9ccw3bf3Kku0oYvPlL0Tp5yivjU
fAZ4cFM3OlEznkAhVu6gxTmfadL+IYtBD+lYg/mU6IzDShP5wfcaI3htybDD/3IZ
PxQJXeSh6CQWCYfxfZP51vHi5umKiTyTQCh/Jb9sv1W1PPUG8ozS+vCzGWQGJ6VS
z87NC4+Yip15pog7zvj2BWOH5ScjddaSXqdm0Vv8436/G6vLy7TQ8FVTAcv9NLjM
Exl6dTw24pBpsgWL1LwL8ZL46XCC/DgN6vzLcDR3vbxMQRuc78a5Qx7d686thuZz
00VGu48K7KYH4yIsTtmcCD+3igO8Rzo7addHaT4f3KhqwElxG+9/cc2PpMHZK4Fg
R7qLVhKVHTJuQHnJRcfpif5Nm5K7Zc9njoRHJdnZvi6egkf5w/G3XbrZijEJpx2D
JHQIogZNRCQFUP+o7JxTAbm0a7P515FIZbApFTHtc/M4ubCdSWHZqUbTLoPvRfxC
3maO72y6qsFR4xwqf9RMWy+DqDFtzkMUMu8ELYhkqqif3K03mAalwiUUvxOkpg7P
kZL4LqTJ1L0MNCDgllkhRMV5nhihxeRGlt7Ir75KIXMgDGEPBGyxp6XlzSoBYy/r
t0/RFATU0dJwtvfh6ncTdt67xmauG6Tnw0dH/P3AbPcISi5j8+rn3vCSIrFRjBoM
y04r1kHQHnmiC3ZRosH3Yh4H8FgbcNVmRDs9XoKKns7XEbTmx5dSX9dIDUq/A0xN
tUr2uLIUB0/1o9iSgFnJ6zEd1RQFEW8AFSQ5jmOGRPLbwa6zUQ66uyQkVWxozpUv
MY1z1aHSdQu7scwRbSpVAMAFMb+T/rwbNRRp2ankuYypPQrzEm9V2vvUEyT8lWYQ
zGn6h3lDMWZki36ahWcUWFKeIYjI/qVKAASXFtfvx/ewjOSsyPG7010mihZV9tNO
0M+dvEiRxQCk/g7IJLgU1muYtHL1lGK3/uaeHY2L125csJHmu0JTZgfqG82SNCBt
Kw59SjeYTtuaVY0acdmdLr+hADmyV13NKdKP5TWO5aVV3mTP2q37LjyGP2ed/CGc
RwEGdEyyqLaiPn+GJu9T08WSVC44BpaG68QkUp7/2n/VKew+TnHs+8JqXoYfptbA
laR5auJS6ciGCLBKxXYqBcpyT+Onyrgx6t6yaW7yR5yeO8QGhFqB6C/uuZ4DHV2s
dLIofRZn7zL6iJLbduYdrXdQmDQcbGGfVr8rZcSjIUlVa+ErCo7AsWceMeaNMndJ
aWQfUjLLD4p0AffM8SEAI8IgBk5ZP3en2iXztM6qJtq0iAbzeYrbg2h3CF4dfJNQ
VIW1K6GdBuV0TRJ5pMGjhzGJWALEe69x+ktp9UPPhdhQMLq+SPywFyRYHwNjGwSN
XenJXZNb13Ui/RT8UffwVUS5XDwMk9ujiSXsYxkCI+FpGlm6BSdGbeN10O67+e7m
btk4m852zcniy72bYepQsw/wZVS1u7lOpXqIi8vqj/iFuRzkna4xqClKKmqaOYQB
M7P4fJiiX8OpPf4fdatXSEr3iQW3tSg4fChzNIWxZ/foO0LauKoOQk8i6xEIUSju
rSpSsFW3gHG2TFSFXodSQ6E1LEbP4Kx+p9xCbgUSPECDMDvx6F5hmsvtrVuHoSQh
qkkf9kP0lFtKgBgO35eV1LuW89TA5hJM5oaZ53R1nhWitJAoGoDSodryMwnCCOat
YfZKKjd1QcMnYL2dVycX6anzBkD3oZLYh5KxAvIDGt2uJKCpqol0GtdG/Ny/5Iwl
Ijgh1vHQ68UgdLdgiAptdWYuwfphmXMPmyt1qEjRE2wCTvCzvEoObArHoTch2FX+
CzJH8uMGvXihVeM4h/kNrGwSpqvDvfVXUnbVHyn0BCDKMhMnSlIvsWdfPL1GoDW5
PLzamASErLp7SPpux2G+rrEzvokU8/EK3yJVO8yxLNljkH0s4bokLM9fiPvbkXvh
R07i64ynyzuW9k9coWgUacQRY1SwmsPbRiFLo34lRXriFLkMSAQbAONv1VcBx1cS
xdavko8+US4X89cgJGL8EHFqFmNvgBeaUtPmXcYKG5Ew/UXp2zgEhO04kJiYerMC
5iq86oZLK6Vz85Xh9NvuP5uiszPaEo+VRU2UZl9QgAJnJzaG3F8VdaOF1G8EB93B
ntgPW6h/hfyXfBpdgEKsFFJjF4noHBJUZC8obDaB80lQRw7u0UpsrAIqhsQR+vLf
liP2TSotK8CUPoM0FTGf5cMGHPn2K1VFVL2HQZuPvXScoKYo7MKrfIzQqXybvxez
wExNKLRSPnqmwGTl8oYU4S3aapfzYu0pZpPlkg3K8CbfXSTCXf6kxLTmyjAp5oEA
IwkL++nNlQR+C0WPgjOVa/altzYubpXFYPykYP2hiVKJSQgqOodGrQe8xuHgggnT
ivE3xuDSF7nkXALoLUJeymfHVt97UFcHhlvUuLvlP3o8se/vqkGhH24EPou1+9hC
96rmhCc9MyQNaNZGRBpFJxvWU/ELbKZvyqNqNOKEJdWSDDy4fM5Yl1pP13DeD8Pl
KjdfYePqRwliz+HLVLAHBykBxTwZWnnvP7PQYSbq6ij8hz76h4sKqHw8/UqgYcV+
NtU1LMQXnrgCSYOu/LsJAYocuEbGbZKNcDSkXj6NL5KCXDanGeaZkGsT5353k22u
uvkg1WdJdZSOGmbUMHx70+XPhAiWqGN5W5WpK/JSFc/0Kn0pkFI2gb3XjTknVsOd
z3m2A44ZEONILJz0RAY7hTFvtrD2UOUFG0h5oFeSYlh2P+PodoLYmWCqmZ4m1fhJ
c23/ErEfmaZgN4csxf8C2pjmcAtFZFUhgrpnRp7d8SEp+DRNevmD6bJhNLw0ajc7
hOEK2rBfHZZHMTDaaWc43kciUsNELjZ7+u0FR5KRuXXc1NSbppR7qGdZvsZnCrA8
bXErJgtB+VZQLY17ofSutoobhD7HL/Ddslc2Z3HSCdwu0ooxHs0Omf/+8Teuf23H
ELefZNdLRfMKA92sI3hjCDRcqgRRGp1gL5KtgbRZMaItEx3xNKado40lTdCLVPor
rr0v9Euw7Di3/Wp1bz8iNIbFcqcA1bKowI22QigEAOWJJ4/l4grZcAnstcGfJpSE
F8emHsTiTnCJ8hWOibj48Ogbm/1nGw27fT00560bcm0FFSI33qLcmnA8ebYpqsmK
FX8IMGJPPInuYN2J/56MWoiPYwbkbqaOGnm0gJY2BV2vKjhlyfyndzOaeXpeF9aV
YEK8RQNSz776sMcYA6BiulO3zcm4oxzuRUGsHke/U9UF3L6kimFpBosho5TZIJk9
35WLUv3ufNKFYXRKsmJyvlZvEhzfMvLgO0s/tUnn+VHCrQX1F99rNzlo+nCTgQK5
lziwdQt80RK9cjXYm2cElIRMaozQ3cW3Pzn5pgkUpGXrVgZ+NvLK+jhfgs/isfut
3DNV0zW1rr4GJfKZibllfzxlIxOt7Rx2YVbyNkyyklNWy3amS2BbB1+z7DSUWdYZ
28RYye9Ej85xc8hA9Uo/uQcuc/DKWcg9ev+iOah4CFD74VHwQdpie6jw5Be+lT4+
GksX40XhGuQ2K/JbyQJ1SLNleRnHS+HhG6Eeqgrd6q3h4E+Ob+F6iX3zRW+bkEDs
UHRi+7Yt9z95NSabtMwdm/Fa9Uh4kNQzNmUjkXavFNC/MJJ/H3Q5u/RghP8cTbhi
O61a5Wubz61+T9LuFdpPytjCEhEtG0IFvA5IdZS6sS+HQYRG9LJThO54WW4ndfya
qPUquLN7aAy9tEw+VOHqVAWJZwt8HkGc0qGJ83mhJkYRjeDVoqAPHqCnrFTDPd+x
D8K3nkrNzdmWSuiw04X5soPZMZtO4mqOcFJN2h7oalvcW/LY/5lRKinFRD8hckoT
71z5kv4P/yLXRP5H8ibdNu3IwIoCAjOpHo63U6ZZI75qiIo1p8SytssiTLBWdmRb
apSwSFvxFYTntrQDeI925bmB8oLf+7fenUd9WWAi3IcQDZBe/FABfX4WOgzQ1rtq
ZjGTx0sq7wRJ5C8qUQVoL66xnl4hU3FNgGOsyzRqPi21q7Iu20FikWlJkHL8zrz3
DG5huufjA58H5x5P/RaB6XhTjGx8/uvTiYwd55XBa0IQubT2swetmBrUSEHv8TyY
chNP8ZCEjBrDX0HJ5IIHIYflDYY4QhGahVnF/gBpt97wW5YokqDsl13iDvydD4Iq
Os3RanPlrwIq95rK8/5KFxu65dq9rB9+ZY6OHKruK4/DVLN2raujuvIQobAie+EP
lGrLbQNV9npiaf2Qvm2eIopTeLpPipr7SC/75S33bLVa5bWxoTrgSM7lj1ifJA05
zgpKsMY55LBmT4SPvyrKdZUrPBmW3pPQ1N4gHtd9Od1jQKGiiw2EG7Exj8gU6+FX
T7TP8JaXYDXK3Z+VSkpZWPEoPa08k+gVyon764c42TSooBd11P94Bq49mra4VX5O
8dyve3Bn2PB2GOd2+si5o7dp1yGEwaiyCzIKaeIiQeb//Yv8y/rcYZmiZzeFVbCK
Bw+8WzC2mTosEnUSiZ5NZYSEr0qFyk55/KhsDLjvAbtdB7SkXFmFOWM/Y4Jb3Ojb
gw/4tHIJkKDsl/jHFdfeoXCEn21Z7WTZjeq4sO7zCatmDe2NPSx9nvzTuTooLaiL
8g1dYUofqb7+i9ts8ZnME4YZMpPF+HPNeVMLPObP/PK4tIYt2mA+ENz1Eozp66kJ
YWDvh+g5JGZtxiAWRjvZjGJZ4dTErgh7PVDKyhMu2wRMX6EROIgyc+8n0oTQ7IyJ
B3ZeVETmNxfe1y5rlCJjzbCIELY3SvvjlE41kZmQhUY1lG2CyIu6fyaL2Ia7b0mj
/TdMVbXzTg0rFHJqNDRtO2B/My7oeicr2EoFujCiPrmvyNBl5MSYtsmKQ85br7+w
2X7KtcyX5+xsMvqbTEfbKGbnmls3oFvfKA0r+WoHDg6wDSMuCFikWr6nR3aGiS1J
VhGaxAaUi51WvKHWb8pniXEsWTPx4nLComDJePQCoBHR/K0s2qxqZ2UVYF2wgRJh
BgoF3104L6Oa2IT2oeuoxwDO0/33Z5NrMLk6Iz3Vc8MH8JX20xSEVlZ0l+CK15s8
p+IsWaxLaYY+muV8KGez1Z951YT1Q60BsFl1PFwRgLp7spVlOoBiuE/FUJ7PBGFC
SWiWB7PlqJXJJr6Xn7ycD79jD1K5v1tmXankGDUMQb+kCr2jBezC06QATX34Aew3
UScHnJ/p1acAZw+BeUlZkM3EJtOLrYH4kSdjFv73MzAbe5s33h7p1kKeJDrTLyOT
U/JRry+UTUMkwnpCsRKSFdFC/GM1ZStFLqLYOerKd8Xz1XcpU6FV9CsXiwlrAipi
28K8xgQNuGMZjw+y13uh4lZzY3IpQxKanO02MwjCh7v5PRfY4WnMFZU9sn/sC4mm
F1736IfFHWCqQ1iJev9D/HX4FatjsUBDAho3yE4FTZFfdsk+sRKF4ND0D4w7WgYI
uQSfkHwhSVo6TeJ0PKbhkQYF7EhZQ8qXIjmQTIMU8tJOxTeyZ7u6VnmqytAHl2hy
8QKozgEl+KobXPxlUzL02v0oGWBto6YN9W0tG9omvdOLCLgmlYk1isNCUCQXbHAk
NVAULR74sQDBmkTp42oeKWG9+1zmMdQxRZEt/cKqaAnXOz825zBrqTw9XpEBkuok
fw8AJZIzttBD9s9izJ3cmEkSY24z7MuXpO+aGrP8zXqdRUoBrKhc0TRr5FOBmy/Z
v4VwkY+sFP0w9/q36b4qnkzyliUb5kJUQfsMNjE6S+cchni+dSr68xU/Zy96ztgB
XHT4CoTZBZaMp1I22mI53V0K3mJlH+Iyuy2ybGSJVILPl72A8MrBRF4qFVo+ooJp
2R24ooPVNYqOkFEfumy4FV15hZUPu44Qt1wlOchupnWu03ROSz5lRxnlSBPqUSsZ
PaZ2KV11xpbqdJw0Of01OIeA87PkhYhQ1CBzfQlu0bv0qVtwUJujxjXO5tWa1nDD
VLPcNk8dK4AEyfootUQjESN56kEJoOBqK7aelMkClEREII+CDEr6aKASWU0J43s9
zysx9R3CGol4q2seyCazq9fwJc40ib3EnBjImujPkAjIQgnjrJeszR6j0lUGxl5Y
G+mrX+Xw70CmTLqg8Ee4Loa1o4mgJ3yw/Uu6Lh7Kn0U6bdcWK8TU4oAb1XSJmhdO
lAAqJGTCHzi3H7uuX9+weRTpc/uCw1AuZQDsXLwQgSXXxDVA7ls9HRPRNcguZrlf
8UjkFI1XORwud2LZKBN4A/iv6hDJ26cAo5rsoRUYvctst2+E06yqboUGI/OtWpxs
QEYdzKKUriKH5FeOJuE8paJob13v5ihECtiE0skG4ybIvLgeXqIB8e4j9mU9syLO
Ud+EiEQoOV63qkZr2+nK7r+/yearHuTwKthxnfPrvyuzJLdp9gFf/svJfHaSDznl
P0jQDCBGay3v+SQ/wqDuXk+SjLuOlzleOdi1jqd2YeYXlFwAMZFbUvP1RzjL2Vmq
bBmjaT3U7FzdnYlbpabADOrJjxzs3/uUAT5WfMFfFs6JUnJ8aJFZT8QFRwq42nCz
J4LBmxNWJP/EHvIEQmPebADP1BmqRzL5xHSHSDCBPE2zcYhKfGP9UEtZAx1BsWn1
a3QMzQmrGcxm0K7LhD+dtwoEx/0QFxB9+kCXZsWSgcFwvYWy8H9mYqM0C7T2y08e
TbQqMOMJ12Z7jsf5dahM1ctc1U2V8msZInRn024D/ZoTNwcI5MFK+zWZWVaWVTfS
VDo2e+ku3GqTAk8/oDm14n8L3RS8wPXz0ao6hQCCc7O8KKQml/UTRgKQ8kbsLz0t
VizWnu//NONcXKQXpdjafeDY8H6gnDbHBwKoT/y8PtPiq9oVkHOOuMCsv8YJwI5M
WBNra6bxAmGc8sAxNh9mJvofDGfySyHEKMSi2+WfHsLvFHAprMKtNckdKWEUOsP/
PrZXIWr/BgaUZsO48xCBWqYHx8/+qm1ulS/JcicDtyWmVP4KJCTjW9kyKXreBxxK
dBfeZTJZ+DrBbDuLfOiJXvjHChwW+ewkRTsvyyPK69l1biVplHpqHM/97zL9Pulk
EI0XAXREVIsGiLuOQytsXt/FtlQKcviX09HsJlC8e2OKJ/NybWW1CWre1GEGKmOY
8xLoQj6dUJtu8B7i5LszOiZtiXG1welPrp1ATbRE0f5l3hLWZ+ZsxoD87eR3uwOY
69geqrQvfWaK9aqx2w6MbMMvZs1wrXtknG8iGR2QTuLrwrXfM+cudJKXNXbuohg3
3z2AUkdO9Lsx0RJAtKZLVHSZpdZHk7EdBhR5qYA0kVRqju5Gyqzr5wNB5gVM0k/0
3FeCiQqS/dSMw1RhrLs2G1Cg6q0OqI0kJO/7A0912M2L/N6HWxkMgap/Cc1K61qn
lQbmpD30op5Q5SvpG5kI//bxrgANjpR6f4zWDETNmNDKSYjCdG/RmTP3Ob4lUvPA
7SyzuqJn4WS74xdOIbYAsLMVMgDqvojffF+06QRS1epToEJhuA91FiqTvVDEQCLZ
oDx4EPvrgm6T7rBWNC/WQ3LDXZUsZ+SAlMZX7s7YC7eggrxhC5IVp+sug3HBqb+y
TM4PsRpxrf3Jr7UFQFEoKlBbbcLfOQ6cSyQwainuNRNmVEvHwkP/ilEClShI3RE9
cJsfCL3/WmS3HRZDIttNzdcjkLv/o2RhtrMfIDr3N4oMN8Ji6m630KYj0cK44DPg
SmSE8Go20pdPs3e7f936vUM0GNqFZFjL0nn5GjMBNdcjWDmi8iM07Dj+piQ5NHMR
fcZ5M79iHSY/+eLZwzzGm2FsmJKoPOzblHskWwZITkHKXeCe6OQ7NRxGIz7NIfU4
M3vgdcaBOPfLDa/tJcJI3VZhp0X53pGkb4HgxbOapEs99a7PnUF8SSB8hiVizhlJ
dlKt2IRx9toBU/yOOBNDE/5KxqHoUOUhI4fxGRap6npLPxbP/4A4tFYhKOxdDXM5
fjfKlI7FyCKPWQXG7iy3Dmky1/nX2eveGKxrefmhej6OnVkAavFxaWS0stDBomdb
5ix1uVpxAra9fHRQOZ7EhD5+Y0LHVsuncWcg4w+35hOVtZPzEw8Vdadxmb9pDu1F
O/jHHa8eLwX1BYS5as56kH7MJX3N0rdBfUv1xVijiir/MYNxZHHbQfQBQnqwaFMa
XKmbK4Zl2M5MU9FqklrLQGP58ym2h60fmrnqdHv4ncY2uEGMTD7vLRqUkkumrH0l
387eFaZ79xlgzGKnxlb3y/WpPuB7otVN9gMYVQjmtsjC3W/xJd+jN1FtTb/Qa9Uk
BWOzvdHbFDyZTnpoOiF8xk3ft7LgKkuhRrt1zd3bVcK5IAfk95hnHRPM4hMufGOS
6Ls48p3Gqw9jXpAVZmZXtk5uKmHr/cYUICJIo3KbL8ox7GpWwsdM+OooSH57xqid
oOFHONFx0W8uGJ3tNpV4dBUB32g8egZAhGllHBwKuc3rpTh7mJNnSDxv34/e109s
utd3kvT6zOuespbeg83XI3DlYBqh2EpJsEjjhi0rqAcW89nYnhP0OOW+8hMLqPtN
VmK0qIl7cuoQ/e8EFod4PdTFQT5hPZQiooomAJFTcrOYXFif5Fbg1NopSNr7CWPc
pWP4NkM2A7DHqvjvf0HhT6F3sIq4Ji/GWasnYWVcqPHeUuw+kMLHTzXmck7rl6Pd
jtYR4RMkRExPeNj74jco5feMRJNYMgrpw3XqmbSRWmP2u+jTDLCHpk7DRb4bFbOn
dI/joq9pPdGLzME6iWbDsEabPUs+sc+halyVLW94gC1wRghNQsS3Opune/ELuoPi
li7beyZ5B2ZW+XCYajkVHTBLQEbZL5bfbQEgQd+n7HKGCvLiYRYiiw+BoHQ0Vd/e
qMgMVMds+flpKA2lj2P6LvzxYIhkE74xkJTD16Ga4ty6xVGroWfP5jO6fqM3DOFw
n3HfBiFrL6TihrRsE1lOeF45BiDZOWcuOXTrLo2uLMRk1KcVtJ7d37M16+OFbRqf
ovS9JTdQYE9GRhD07az+iZAk8b47tns+Dj/UDea0BiRpcMr3i0VwtOCAzWxwgJvU
y4E4+gpzhx8t/2nxhmvszZdPRJ+UC7x6KPu7sDdNpVGeMWi1TQw56VzbzJ5rXN2L
SvWFP0LJcc4sSLGiMnpzX3JB9Lt/c75KnuTPgKCzlfQZKw0H3lFgAuOLl21Vwxy3
x8YzqUJ3HVo1C23Ujix6NlwzDCv/F0q8rr0IVOIYFzFzQ96Xs3yMoBhEDbSx3P3O
vnzpQhGGggjreLsfdPBtJV9tiMrqr7djG2DiTfrs2kX7fzRqHNUwDby7C1VFpl/T
1+ZGVH2LDyd80RwSsR53ecDjSV52Id56S83ZTEDxJ9ofQgpSxNICDWLuf3b7apva
eYK/36cPRMj6ZkkYZdVGYelWVzXZpzQ5BZIlEiitj9rCfoBvYqeaa3TfELnpT3YS
x4f71tfxg+A8eUfKijQRnKlkVvMoR97XCAyXKUkntumvakZem1qcpJYdbX8qQCv9
he2R95e9EYFeuQGHqZR8OCVLhcQXTdGpsh7StlGoy4+2yWyXaJU+uW/SB2f95z31
N0rBlk0fGrJrU+zboMb1wX+xJA1ldrBDBYUNC1M5I7IkfuekY9Z8MMFA3N18OtCu
BzkKz9MSg1l5dxiCbeq9AtI72u4boq5t39K5Ch3u9fjAo7IFElNOv+PuII7mt/0R
fbxc0jt+bOfkF8UI4XlzAOUq800S8HkH4ZDti6RWn37wA4Pr5+JJvvfUUbaXvyvc
7LhMvFqcWtSaHFgE/XVd+QUAqwzxUD7zQqyMwPcf5mEXB4cyBnD7lpvwaF5uFuvS
5f3HhDYqlqxui6aQjbB5z1Qd3voGbBZkqNCP/gR1nt7AQ/sCOQwLAw0gZqz8C0qJ
FO/7xgvx8VFvlSeBnZMrl70ovESA8lZBH/5TYEmsE4HUgCmUXbqHSvl0lYtvGT3G
3DcnekErm0+bKxtmWudDE0xjkoLDaGHJ/z4E2eLqIvOVkb3hlRQ2QTNz+iP08ma8
iONdD1iW281eubAurQBk8qgB1ERTn0rsHH0lGZv8SHghAiuO9ohMpBPj0McyRNJI
DRreBofu7gogPwTeCoPM4/9XFoBkJt9QvfYdrU+g+S28V3pOuzmPTOpOc7VN2okk
eGy+yW52xcMsExCs6fKLNWU2EbDnSE5rGIKvnzSc8/hU4hAymVfs2VxKaIS1BDeA
Tcm65c4xkQgz7hr3cJFfbnRWud7Gj1CUMZmHoe+WOoZ42wSOHY7TI4tW8gxHbq4V
Lbt1vsK/E4wF0OJk4fBAZ6NXNgMDYA41zTnV5Nq6rcsRN3kyMIiqVjktpeMbFb41
LFlMGuaJG88IbjTKbiwHey20d2bGNRL5JXWHkSP1eKc21/UXwZFPfLchJIFN9ffX
xaBlCs6ewzGhGW7pNfErFDusxncO3PCobYlHEPCsbFhgxxDFhp/wsyYqY1ZIRSO7
gT747/Kv8iSnICOl2FM5FZHZ+vLRApAkCuQVEqROg4vfDehziaUxr6hXSgIVAixW
X1BSM0RbXTzI7qxvdxwlw9+PKblqMQxF4AF6iFdQCtYtikD+k7zGkCcEeBGV4QQA
dt5csQOzHbPtJWnKpXLSjHtORyPEN4YIHtWCrMOk7SCoJJahbv2hQw3i3yr7Ff3z
2mEIyZmFxXQJqVrtO9ByZT1bNy8E1zU9U6qOXOVYmiZgevhhiEg9MLW+34Lu+pEb
ZbNBXCy7TOSUhZrd1DV6wZ+ryRr1jK7tDOs4hLMS8vKeVRhuzNqBDU0wXeTanatq
3nMm+eZt/xr6NM4ZPofzVz3l/u2zPEh85umTMh7qRF6KNV0X6ViiefbZ60RupUto
NDQW96lUCzK8eaaSYxTg6gZvT97u51/tGam7gbrb7GzgpRYikzrzmnAiH6+x6hBc
n/zlJ/mo5DYZpYwRvVpZ/mnBKXpq+pbV1ZAqXRQFXRE1gJRm9KnUfmYORfRYsrsn
srk1O/DJ5xKURE8+i2U8UxafEbXoE1doGFVH85liBmzaA+sE5P9qkcYxMkn3kL1p
quJp2Cy1mJXwT9g+gjY9zkXRti4QwoaZGSMpDy0aDDCwnXoTzh/VaErNPenOK+sO
P7dP7vBIXmmr1aE44Uwe/cpIWd9tbvGI039MmDu+zLr2g2tBvwfn+IIP1FEEhaB2
fP207s/rPa4Urx4P6XjjGkY8KntHRfT42nTQnSAWD5RFaw9Z+QXvTBGJHrr5teXc
akghdp32wchbCZgZgz3KvAkC+mMrBFcO/VyhJT3auDtu4ApWIjRfH41v5ucqSy3S
qp25kUy4BEFragSb6o0hS9C/QeZ5Y7+PtPaigqzq0oMVgR0NsXiSwL3ZZg+Pa/q2
qH4aPLcUFxFGc6JmYL4nm6aNl+d3b5Qxq+YRuJVPmk8OnWNLCHFdKMN1LQbKlot1
pAAxoerz17gRw6MXJh+RdG3xJjP/YuYFXZevnIFLfz1Owqs2i8Nl5ELSODm2OWg3
daGbm73VaKTlq2dQUv678pPwbc6YJsj954yJNzYFrJNbQvEXKg0POVr7o8I9l/Ox
lOe+TvHYKkLjUJjLYDYCvavN/r4ywhkrH567k2xIVKBMNWvH6xbsZDIdHb2etoDp
eMVvSDSFAXobiLR7IgzH0TbXKdhEtVI2kZT7aAEcVI2ya2QuLZK7vgFCho7B4s7j
UqA76rPdK8HJmqJsfzPqGtyD/YpCNfiMmRWa/4E7FpLnMnajyf92QE4dc84Et+go
Wvl4HKjv3RxikJVW7b9W7B9Ajjyl7tiRZHd1GgGEl89GNpWjBeySuW3xPUuOwFtr
Th2Ts4/YTzBbZDQX3oGyGYtJFF/mgCXpo9CXBtnKaN8AGa5Wx2lqwqF89UhHWrds
cDqMVIdLytG92LMvYmNFqZmxOWEGA4Yx7L2AvqOOFIsVZkY9lyaSrL2fxTcuKhpO
1kCqVEeanU+90L7v48pfDYiUn2yhhZvvZ+9w8UeNDnARdLAI7efJyBuMKiwwxHNI
KSD/EETh2RW3NWLC40mSjeihm39jTpBPx1KIOVN52JMoyteyncQBgFhU7BpfjRYB
4dKc6aW1U86F6QQ9xBH6j6YefYaQE4RX4EhO9nMrng0kBi9oK0gXyism1j4YuI9N
fQZ98pCLIk/SJ6b7HA5cEf5GhQgckZh0gVLOxuEabRlCOyCEZyxHvJPUHReT/QB4
c/5WNO/ETxz90tXGd3axmLnKhHph+y0UXTQGzspML8rBjMTotvIRq9LnC1vpOYqz
Zckwe1e2QSiHVQuQtlpcSVFU86w1LrnSblLHNz+qJPmdslkylHb+sHdqSgmt5wkM
lFhnOG2+cF+n8/Aya09XScIsKXLr1+31s5iiz7CwhFVNVJXfRfLZtvwHIXU/w1ef
B1kjvDUEyCoj6woABHMVljG28tFVo2PtsKWNPyTgs8hlqU1hj81yiHTYBGRH/bHM
lCe8Mc5eZV6giJPeE95iNokYw+p7VCzpMYUa6yg8L8e6EpXJIgPCR6zpJORtv8CB
59sdhrTuzOEUg0qXNV90a4TaiVhIHXIvIuu6UtnGr6sDIfxtmI4PBMkRG9s42OQe
8fuZq1t0+DuL5EdJTwiBP4cG33IJzoorU4aAmXVeUhQOq0H697g5MBkM1fkuetNi
0onVPYdBp2/k3iSImLTez3DTGADhIkUqGMiV0PyjwI6yIgcmN6in7M2t2thQYoTn
X9QoPsnfMsbsnAtKPgeR5x293UvxcxOrk4EttfRXmsbse4TyPCsJQCNg6V6oYWBg
228B155UC3210en8IMqNNeVrR33xBDA6bUj2Ueww/NsnLmqenL0BQ87XsJeGZYBL
d+Nmuwy7ahPD5OgZhMSgWygk5A6/6kz7Xg2kFCE1ZNxTvrZlps6Iy36rTaKw7Aiz
iv2mCKLSU1BwyyU8BIxCsr2Umoo/SrEXmeRfHn/A3f8pBSjOyjI8y8O5JTnSMNiT
//k4HFI03QF7VeB+T7IvNMMBehp5gZVs08uqlaKX11bu+Tgjp7ltSV2QE8OyKXIJ
xy7Hxnosb61RifAnpQ07VEtLzuW4Ti8TUMSF0ol1+i4eVm68Bst4v0434LUBLZc8
dl3JuwfODTELae76nJgt4Jx4DKXZcN2mLhA4xiOAM70mRmDwZWogvrWY8QFT5pIK
7pNkS+++LeTZDyBVqTCR9aNFX2cif1kDwlMJQj8Ub4E5wnOEKfJKz1DVsT2SdUFa
PWkHOkPSUjF4XCPDooqkQyTPXg8H4te4tQO2V4DbnDUguYMlKwi+Q0SzcV3K6AXH
lvybp7pul6czXFuvxf7c+mPp29i6CUixzYDCFLeuc+5/fIT6iLN4SR20Gs6VK/LB
/gr2tVQVdKpFE2u7F++VZX90gA0FQ2umjruksN1pmcy6qAFoIKcnrXQzBvmsD9Wf
hhoDh8o3mrXxSXQOYlBnaTG5hwDVubrAUTtx/rx3rp2nkJtfieACk43Y6NIGNYc0
kHjf2bZ6xRJXqDADFlHTTrKoL/rEN8hgyzZyrHZjfPyVsN+QkvgJhFY6w+5qZs6+
QX6cOaRx0ZWV9A8ZJIlyfi21fRhqt1CWmRzT1u2Mcj827dAgpxsp+era5oeN5xrf
dMDo+GeAiWILVU7mx12YkT3yeiMmNcQKvRO8iHQ8RiJIHtpbtJtBCWumnbT0xtp9
k51UHymp6+fPbsPcqKoIwfDi0EcY5e2ydlLReQwszvnuRxWE0E2T921SVHeuA2cl
qpagyAXVBPYcbKktjvT3wXtIveAx2tup6lKK06QD5se325EMcN+L/Th1tus5GLs9
FmNGNnvO4NTB1OeumWoJp8BGMFgBF1uHaKA2MiPG2SkwG2Y7cjC98P5retn3Bvae
vzHnA8/lCmAVjBadXhzYME4zG++bRKF2QaJQzjpHbYS3WbHU7mY7rc4h2EYCV0oO
UCYT8HSU20OfVU8PZRmWJM/FX7P9/pgZ8K77kLcNryFLccaq2n+hKKGpUObxW/GE
vyOc03NqLdV9991CmiOwsR6SMOBX2fXXKUYgsuoSuElWP+0nPLQ4uKWzqThaIL0V
Ezq0kCe3qPMFNe2A4FfSrxdGMqNpJsF8fZe3+EYXm8pgMW66tvORpmz3XAqVlFKe
tUhOc9TzVBlKsfkdSb9qcpYXooBU1Z5/h7wL6RzebhU6xPKiswgWONydNpk+67Vc
gDQ09qUxAH5o96c1GUyHfzBya9wQ2UJ55MH7RT1HL+wrS8yNYXWBhv6UQuusRpAj
chMpelFC89gnspyhLXL+znhWZkr/sQeWzV+YiHTe4TJTuOZga1kbFlKuenLm7Lds
tYzSAwgUphRJGtQ/AaKgBHEMOZXnH2d59M7DNrTkiRzgXd8IpKTBNwM2nsk0sL/+
PrVzSBNqck31mCxevbjL+HJda7SLAsBdpJ/cSyBwCwUzBLNXXEmAgdFR3Ifm3MjM
6X9r1xGyjvLPfTzBqXnSt0ROXkyN7YAY/29E8aQ327T698n+Xcz9+N27XE29M5IN
AJA62Z/wx4ybOPtFk3Nvt0gM8BRObmVWCEynfMliomcPOsy4ON4M9uI+ZTLCUk9i
lts9+YOTwpbltsEQ1bPMwSZYWMpJAFyOIeaw63LpBN2EhIbHPy8J3fBXWOp/AiPj
l5jGoV+3ut1szdoG3eMmfBXd0tz9WfLHR1Om0EHkJCMLln43Hcanpmz/ETFv397L
LojFHfPX4M4rVKFZc9StO+DMSGlFjTPfsxtRS97iqrgDPtjP7EujSQkU1aC971pq
2HrC60rmhby40WsIak1xiyFQsAy9nE2Vc77/e5UoD8CDtmX7agI9QHczCZpc3JCc
ViGJWoFjYCZoTDJe22eIx4jWiSZtIC1URH0uP9Wfc0a50GgI0xWLbNSmptZOpfwI
Q+btkoNLxWXFdVdIvTmGa0MULdXM+0gzuFMmFb31w0objNyqjhlQekEqkfKO9Z4k
X1mIpD2k6mroPNAb8RuyTW18pcrM2EItcL6k4NwSP1Nn2IJq2Hp1zKYD0ul6+oPC
YPy5X9oOxJ1OBfTKVyAymcDhFKSQt9vOOpjAx95eHaSpUsSV24YjCCqA3Xkvngbi
Zgwk84EP4HLAs1T6PgaxCkq9O8TvQqbN3yC/wPRzPPQG0iZI5VbXgn8TrfyQP4Ti
c3hDYwJMP+UvCxiGVqK7rhl7orn/6b3i6FnN5mBWiqt3tWtw/FvI9ZsNwAhZi+Rk
0tPet8fVUi1wNGAJd8T375S7ht1f064TGy0roYUmRD6pZJQaE/iNiVhTCWEoq+ek
1AgorQwZHqYEy+45HM3+QlyqcRqKtcyQPtgEAEghiZtd5Kx6ErpbWD4rVXyeUC/c
mtu6A/PfH6CYOnGVYK0OypPk7Jmne3sxLntbHgJ0pwUE4k3LD9DNQ2kJDxaaMdpT
JoBso5OPI0hrJBp8pEACciQqGjj/JKDrgnQy5TjXHr878d4LZNREfUulQxR9e69Z
DbTEU0U/oPFDpdCcg3qYyfpnI1PZA0CMh8pOTWmWs2ko9TQF/rI5vLgQAPD9CHyc
0X/RFd5eG2YWvmUfoNlo6WRMTIxk8GeQUABkeCLaYMkvM0Fmkqz+0oOns/DJvGBX
8Q9k1Qrc+bf/p7zl/3YCiD8aUW15O8nT6awscfrMgW1HLtr3x+tFqzqnMbGWVxRv
DWNqjVYxpZR1VcNq5YlZPIQ+dwaQrWGUO4trpZzuEhbZ05SYoZL5sliLUJV8QrBR
jPlcAZl94Cn+Fs1xb2nclmz0lfaMyrzDYkQ0rHmzV5OQzlvVWhtX0AeCaXEwuTrG
pIIdbS/bCQ2UqvJgfjjEpaNMTTwB4VQ84hNpCjK1cnSfHjXsewjhIuDQuQUz231g
faWTwdVp8J2dIbNfzsoL4xKFh8VboBCMfBFmCgMeTZj+PJvQAVRbT5JwF9hGW84k
mMEqZzv6fevCIp4+G8QD95Fy1AvUv4APXgXSrIYuXn3Gun1uKLoDvo23y8BVwe6f
+SZdR69z57vNXbroo4VDu8H7BfRWHpSHAzyjZiADBCfKwagVB42UB7f+pbM/BnI3
yBg7L0jvOwcRuym9FlWDoAgKRvi8Iys66PRNgn02485u2/e2ODdFABeacVVfsyPZ
ToBsplV08LDJWTo680Cl+kg1Tm1yz6+aSEYt9JtSXj8Bu4RNR1y/OT64Vf10Zzki
H+tBleOv6wDoMNTJhDZIsJM0GugEkfw78J5b6BAd1Q8EYLTSj8CDRku+UDp6djoM
aQ3riqj4lolVLTVMi8xzhphw4Cs7TtcaRVA5gPn5s4oDPQsdL6DCayoRGUrs0EFO
eZvH4GpBk5jww5CIkJmgLfwROJJT3RM1elSDEBZt1rYlttUi5mpOs9Xx7CajVB9q
To//9oJ97VET3wtcSFgaTxKPh2QSXnE9kXXJrob8H244SUYW5GsgmaRrx6aBgDB7
gitmIPVyYsmzCtJS+e0GjiVlIgRFFUUry9U2nGkbCqtwcNdYAcq7TzyWDs536pBY
RtJ9cgmHzscXhza1ctZH5ljWwEl7z/24L7nMdneXB+6fjKHQ+tV1+Lsdb2aRQVQH
RbaGj1dz3YTNxTTXQ1TZ7wmzsAaU1xR+JZCTvq/PbqN8z2XwQV77iIKhWxBZaV86
FwgYLyEve6LnPU9N7aTJLSkW0xwkNzatYcLbwvCfu3bBvxn0mTlEN0P6bcF2K3l0
iAevSUp/7scXlBy8DEs6XybvJjeHfBp76W8swNurISdMv8ff8drgfyG8HA1hICuD
55exgrt2xbIVDLtkLT/Ls8STxg5It8DAGvZ8VuSAgsDjgy5E9anDTIf7pZA+53r2
dZ899B24ZCdl4xwRBKSmxcX4cO3MUE/Erw2zUyU22ZumVTKne9xbKBmzsEQ+mVyW
b1auie3RA2H6z03VLbRHpOTu3KUt2M8MAAYPcvKmKgR3JxUfKJS678E0jL+07nya
b5d3c8jo4ZXa3BAqnl+UPL+rtSCpF4Xr9AvnPq8Eb6zOx9fPUtV/oDwjRvOZyBOC
+tzMAK95eH8i/CL7F+Xjx0bGEle0SC0kMUemZX/QJtYkIp5PCZ0SMOVWxr2x+Ovf
LNKCukACacwrPlAMFIIRM8H/VhWtfQgaLLciQx3UfOgRoF6TEqIERcyXO7YDu5E3
6V1HWVg/BVAW6yeQHJmqkEiWbD7KvA+TCuVQ/jWjJX7aV0+g+Nbi+t/GaYtPSfjG
L8xK6jikqOce7RVUnneYAWNOuGR449ZtWNj+b37od6QfDZjfwV3krmHFCg2uDAra
e0FDz5Tj5CXpTbR8/UsmOokcixlPhU4hckv3+SuAOvu/h0dczcLF+Hd9j2KRG6Jt
P6G76cL7XzbKy4Yaj4LncfAA/zeeFje4PsZlsp734KuOA3sQ0YNdtWPB0rSFqZ0S
MGBPyTEtn3Q61w89MhQtsxtQCXRnBEXntdr04N9gccK/a7a3frIfJnGIM7hZjp9V
Ki+WxFlUtHNVLDxLHXDIBROQIf05zFRlk+PfWhGd0Igkd2q0kTOdMpUak3VonWJW
RP+V+/uKmib0EoLy/eLtoVsITGrQhPYKFGB9C451AMD7UejAPcfd53T1yFVrBGag
IJeLpdtL6NuX7zX4Q+v+/JiZgPrpsEzA8ta9htPy3khhTnm6/kpPKXVgjfiU7I9E
wCH2Vb02D8qfP1d7HAVorZjDoLAH5sJD/OUADVq0Xel7HxH7DEo65Hb2sdH9FxZ5
jUOaB8ZrtlEmkOy3kFP40k1JQvHml0j5Q0btRQyGDGe9WaCXgrsvf0sq65yDcS8n
exB1cA3gKtW5/KY07oPzCHOdb6r2i9nXodzV3V9mSrOkd83DcVmP8L3+1VMJaYYN
Ry3cXK05mq84JMMKy6aNyQgBI+ySQc21kh/XdII/JJbMY1ZtKD/CfypS3KatkCRN
kqdwsQYT9t5kd0BPlj8Kvs39l2D8g0cvNnczld/YywwE+CZMmzvrKj/BF1NdxXV3
or+aqxw0mmIbje3HRbXRFwHwczEJF3fUPbNuLDnCOEFwiZnbMpXTncK5esomqJXI
/aL4Ldhr6j+4+ajhyWAh4u2JZtcmamlK/O+j73mio72P+pfUMD9haSm1mfIat7lJ
EgiSjQ48aRyAmhSVHrE92V6cpS6kVYJIvpEWjJbr/8nPp0dblc7UdkHKVnb9MXJq
tVW8Q9dFaD9wpaqHesNyzG/MUJR21XgokrArH3be+gvEqVuG0Gncj/TUHYw0rkV5
u4riUpm6apjloDYMiUN02cJ+9xd8J6NxavFlt0BpiQTxVIqNvDgA4RpSIDNC4+za
pCTbZpY6qcfWi9AEPT53iau9134AbawnMXiLd+Vv4qK/MtkVXWSlhIlFKI7GzM1c
3XsX/9MXsI31990g4jdHT9tb86b6icv7UsshIOGLil98Z2TRNnyqPBt7EMRcjweP
JN2oeElgU43+1FTpJWYXCY5YHc8fJ2pSrBjEx2AUVK5lVBtn/PIt0CTMNLhNSn9m
vKG5270ZKXqK2Smzr1HzeHMHselqKi5peVRqIK3Qepnda03HsXJP1P4yFSiBBunQ
OrXXPh3SoVxDoCGkDNd2d5KWrVJN5+VOxAMzjV5I7z9Uoel27WosAnbpwpDL/Ai4
mWu7soimRn1Dh81UArnztgiHZJ49g53tgk0bpqEMw3ehe8q3mJwUKdgzV/IMZ9Va
63Uy+B5Ff2kjtOfx4obwWI1l1mrhRFRJjWzNGRB4YP0GAClgxCt13+Nbj7C6bR4I
boFsqIkyG24sEz2kSLVoc29ZoZ++7UYZueJBERi+WIInkDLRhTo5E4mtcQixrTME
T7+yvMhKOLw2YbEx9rk3MJFyQWqknFeD6a8nX65DV9ykkz+Cnns6KRmNDI8QzqKM
JhUftw2JJu6TVNXkud4kHmNcDru9CMXSq6YKJW1T2K95Nydd5e2/A+BmlU60maEd
46l7qxjyl1HhMI5qn8ofk7xNhDxHreKXsN6ZOernnNp+enHfjSKTBJ3dRqPVpjAI
/SScxC2FSL1bUEa1tdcJWhgsVMSZOEwUWIVeMdwlBhFQ1b+j//PGBR2EiSzTsxV7
HbJ8t6ssbC/71R35xWRRpcNNnZtsxvAaUnbSgkMEBqeAgXZrhrnt368LYWZBcVWQ
rrNHE0kg15B46Ugbioc/2l6446mdjcMHZhxmPCGK5pjjQH9rYbvfBE7ytOY2duBo
KX7swmB6JRrsVuLavIyud+FKWS4bkQOvnTgdlQ4t2OH7bhYGy0QZgmxUYbPcTJyN
8nkWL+NDpU7QE5JElwwry4pDNpAUCD6A10t1Crq3ZGt2YaFWOT+qjXBxMFq7G5sW
zI0FLRBsqst0Ar2kNV/9+et+vwfynh4uD/RzT/zO9ZMaNSyJds7HgZEOjKbzQIOB
5EmKY8PVTwBqvL8lA/o+A9k9o1MGB3IDoEZZiQh6i4jT9VJNKOITNGTd5ldGt8vi
ChHVVm4ThuWUpRc38CouB0g1WVMi7lApbCekqxEKWFGzfs7x9J5sLAVuOyrK5JNs
y8f6CZAWMxwFobFy+Cd8HVsSjtGemdmfagF4/sHMITZOuYe2qLW+qbphrU+SgWA+
0s/wimuqoBmlJVGDhxaNE1CEvWcMINOV/vnB2s9AvROIAdlSy1y0hTOoX0BClREX
vsavaFSX5V5QQOfnDBZlotfRHXnNw/wnuSAlITwu9oDEpAa38TPOGQMqZdrsnNuD
OfDP6TNsLmmSH8kewVDyqmVI5gmPXMhsVMHUT6+zaXNqO2U4wikCc5llZ4LZItoH
RB5y7+j5uLVrL9FfvCJ1hQZK7T1nzEI5kcAn88S+hZAuHwcth5c/RnAb5WJP5uLQ
KwPfmkrS1Cz/oig3ZGf4zSW+s5Q+wkvnHIpZl2z/cl57BO1vu7fba0LSVfe55FZ/
dQsReyBK85hfHWMBslAw1Pr5D+CbD1rQgfuJROfBzKhw8PIdhX8ticpLqrUNrXAs
kvvEBpZklozTE2FWH0d/ijYDbxncCAWrtxOwxp9iz53dOiaRN/1o/TfDPDiUjweq
6Jjaxh1EfWwAfnmpoEA2ijNyPQpOoA+/eQMv4kdTMy4GX+mId0876y0FEjghfeB6
5YPZLryXRm41CoHRo5xnFDUZStbtYoXmicy+sDKJmpCfGWHMlNNkpSASchV9HQPV
tmPbKsDbtAiXN8M3vtSIPnKPe+PDer5yw5O8BB5mshzNbOt012YfsfchyXqC7+Ts
Jj+VOqyr7oR4B0eHDRplZltfIHbwCJI1gzVvcHrz1XNNEDwvgt6upur+kitvovXB
252odSeYdi//RrdrEwy1KSXBk+t0jA2aE3upjEcgE/Z/vWpFw3cL8VfkUqn7HM3F
Psxy+OepF10v5ofyPgiBP0G8qM9WoIJ6MVTyasWHjbOGcUQB8Wae9drewbiXTlMR
DprE+ZIkH4DTzVlZXi0LOWybHBPtsiJHzYOyLNEO+QCTyE3BFGpslWs0lNoHmZsE
7b8CPrv+4bKczpPsagJtT8/G0HTqlX6WIl6ssek6/pN6m3FkUtBokjWJ7V+4icLk
G7SPniFdss5JsiSYy0aOakN8W0cJmdokBnR9glyl5pOfXdnhoFqv75W5kwnJqXUt
n95rl1txv4msCYHeJr1cwd7uu2c3lMsRKHRU217cC/IPf+NhMAvoG+mpqMGW4hqW
6y8x5+MMCCIG5MGwFxFs/V0gv8ese3Ti9+dwfyZ+pk9qs9XYLfprhmwv4ZtJqCOj
stqLLPl9/rQm9AMCY8mct61UWLx4KHfAOTOb0O3vCOzOEjATZhEZvIS5RpNDfCz+
8Q/M2F0p4S+ddKOVUsiabu9q3DjHFVz8YbmWdfp+FXHHlNLpdU+AhjM9bltLhnEN
1xgOz0or5VeFGSerlpc8grznaZo7gdvwyS33uNm/27GrQXszO11AN+/aDc+EItGA
AFmxCcmWYwAWLmjCQLS47YTnqInzi2f0al2bht2JhyQQugEPy3DR6v0hQDJpLxam
v5O0YdubEOYXOgNsoSNANzTGkbW7NINT7mVePa759NkjkIKkSKT8aU9vWD81LouP
17+nma7ZYMeD6k3g+hO9GBFTR6AcD5uCtq2d60t/9PEEc6Wyvi8r++kZEv1KiRF5
/58ZU0lTJkI9f8yJtjqzjlgTGfPu+3vftgle2b2gAq4NjDFCRiMZ+x5v99DdJRJV
cqHmDJo7Z6c1gxQ//4EmPqHIiFTYjPXVDd9XtqygnVAAFcYuccBs5OvEulO7B1Io
qLtODoByQgv2ZOikwQzoR/uGcK1bYrihgG+m6lu1aqLVk7q+kv0CDbl1krG1IH3N
C1tw78aSFMpkl1AkrmAprwgZo0TJPjuZlvzL84nKLAGbRH8E6OJt8eBKR4xbhG+0
GHhrC/7ABd8fDVOCNhaDeMwZ/JH7we+Z3pNqb0tpc0q5k9sR8fsHzF7xkXAqe/1G
r1mBlmYRmfU+V35fQT1Zmsc+5RFuyPJhZ/JSOTMunNPQB4U9d5eg3FkF+JuN6uaX
NE5/LDFah3737fl0zyAoIoqghg7jblLE00VPdCnvFMaehaeRgtoPVBR1uMhcTPZ1
Etl3eOWIpK8/gpQIrpjYhgtM/qmV8tzI7H9NvBgp7hZGZ+3EVfBvn2SHipYVo89T
rvahw2Jj99h/HLchLUcavwo+Wj7xDYbSoQQZjPXkHfUOGGHcP+tY2vqZg9tnLsIy
MXc7WFDPKijOwp+2S/1j1yGohvp0W9WMlEwSphfxP/8XSF1eYazuSEoKnZ9A1Pmc
2nQbV/pnrbdxM1PuKUHsVbAsc2RnGHtTKCe90Tt7AuiaqkKa9wmvD3N2/7jBMDbh
PC3Io0DQGvQqTH0L4aV0brJCqW1+CCF4qRhHhPwqETOo8pfCEa+R/WUMylcD42j+
TJKdgjF6tklCZuoS0zwcpHsikS5q/7309TMzi+TWo95ZsQuRgAADn9S+XR7iYDSd
SCUn1vxy5Ivn+xQHrEaaKaRtJkm7He9DFIl/sQDPcULo924jSgeVlgMC/EdcGrfa
cGls24LquSuBOjOjLXA2uZTWKkFqqw8z5lZOm3vyEdGihR9JF5+Ikyp4w0tGRu4B
xK9xxXsYW1p0YHDGMrYU0lprUb15yhJeh0WQD7jBqDFE2PXpIGiBC4cyxnCn0ni0
6asBdOVfZ/UM0KkFRwQ52JmUmU0ZNdHE7no5aBUVdpfrQEb1MKZ2EBwFXY9EaxAP
6dBaFPXVevgF44DgUQr9grxAEPZJb+RqP08Evht/NaC0Gd3d+JyzvyfvQCTILbDC
fR9Jwp4Fywavwns2wifgQaCq563Gs6oUqfdMPt0euOAG85BiuJQQPXb824/qhO9U
EL5C3i2/mN0TNliVAoEvuEY3cK/edngFqpewBjux6toDEXL3+08aIz8L6uyi0CdB
tTzaaPThhO8miCqPNDB2iOQJIWb8RHcsfaj0oWc0TsPyZlEIhEA4ZdoASV6Ma5MN
Z+2WPUebD3asQkXG32GvzeqbGCrJuORTPKwjucjsDBvl+D8cAGWrva+NjdzSh5br
jimPCnNy4WrsaQn4Sm9DXp46HdKCpUfY52S25KBYOpjbp2oBQ+3IK79patvC4n2j
SvyVMldPR4YB+ZDwr39dL8hdJyJ1LiEXamenSH0XbjQ1YqJnh+VqTnsW3UFrRM0X
ukywHIu0WAzmX0N6vN0hYyzS5Pvex1DavW+TvqhPtuJu5iNI9ZBo+Oa/6Jr2Qy1A
BFk92+eVX+KqPaLuBIJd5e3TknrqYma1sfDanwWvQpqEmcRkU3B+xyY537sCHlQc
H9j0jt3vjojVprXJR4XPN1BQoVXKt/1JeYtKG6LU2+oDqe0UbukDRlgT6Emedev4
z3/C6X4oLTkJOSDInEUtrEPBXQJXy71YIhLSsbZIaGhy6DsgEIiN5VWQCS4fwaXg
GkEzF9ioG0honi9pXNTOJZ5ZqcRewVJx/WkxxqrYhxkyQUDbAo6Uo86WU7I79FcC
YJMLNlq6FXtuUuLhWZR4c0blEPW7r7jSmVjlBYG3duF6+Vb01kjOeIdbQjJkZlvW
CvlyISwouBgEnoY8/gYpveREkOF74hVzY5z028F3NBxrOPlsrbmRLe3rBLF7XpvY
Wz7VLYCxHqFHdpyguHd+VUDVSrA9vyNbED9nAEIkZjqci525IT9mL7apj8zxavG+
nxDkbMv4vLx4eimoKvh2cEFgex98uVItgmsuB+AX2q0WEQmn9rUv1T561dfiJnL2
4Vw2+sYnHWu1CNa22QolejLVKQEbJVJF8z0FnJaFe51vRHGlmt8i6+UjfKU+WRRX
8OD7L2kWefzWBD/+wmjcMdKUIX8WrJBdO1YtKj05DdBz45ypNHfd6SGTgHiJRrYR
oHDkXDFgkQ/zdcMeO3I77axVPmPZIug7bZm+LtnIMIuqJXA7JCAAtTbZ5ptB0ZtQ
1E6EdFE0cPkWPdP3ECwLjv2qdsow/ryNojToudYOJT4q/6DvJq2rN42fSqST+VFv
aqzXZMboR2iwZybPNUXVtyXTg7/D10Z3ENOpoLyELqnCqhJbR4WShtuSwY6QyFSV
FriiSykKk3jv5B2qnPiT12Vzk72CDZvWx+Zo5MmOshwQG7hVkz7ZSKIOC2VVHLY3
pq3yYIiPBVzd3cIKtaJPna0iWvFBmpJjt3bUPxLopnhLLQgNU5keiiYkOACa8Xzf
MNuIYxuSPifgmTJcfzY20OMNOMyuoKAZGj9fU34ZdlG+ovLvP7cWXxTlb1na8F0x
3EhnTfGZLOKAiZV28v1oEdpYgpYtXhcfGq2T3i3X9b5wFGvSji3VbZBpAA21qNHF
WSCz4FS24fBFMrqGodR/VpKaaKcSQ+izhlSzhDF6ZlBTDu7PYmjsopiliY3iamU3
9m42/FHIhBrLKnmmWGP6YNKoM9OJGdiPV3dvauGuK8v/7gxk7YV+x+QnVixwq5ou
wd/1oXWkrDpSOm/GkHjFpSQSicCZ3ZHHJzhDfqq89ANp6OSg39FSx9GxwNpESYK/
TfkgbWfcDbd/6ZpLk+kb38uPV1NrRbNWiA9D/xwmJJDyrzgt94b76VH4LXlXOp2W
Yz2aEtQNlx6/mULjTDMz11TXdC9qFgsk4FqfzBc1PzTywpsrSsMzjEk/LivQJeWl
OJYYoyxs0WGP3Qd7LTiTl9m2IlcTDygzFkL4MW6p2jjJFhOtjL/DuUE1XZCtmQ9g
3OM3TVDTixmNcHvm7wGBUJxF2ySmQzTMueTdEVX4Ajz1iTi2hlw19AzrnXqQ2XWP
Q0vCYufvX2VzE5s7Ck0EdqgW72sxqdPvNy/pu4f5arIE1WTZ2eX2EUscka7jW2Oy
xo/wRvWAyiAT+G9Q782wSEd7G0GNRfDDHUz/pehMDNwrTAtQYnmLrv6HG/rkGegL
nUXRfQcXv9HAu6BnmCpzJKKlgLZBd5EWahqRYBv0qCuO5we0WBeqIlyT9YRHuH/w
t14ppXp9+ez4r0yZW1C3s7cb0Pq+cJzb2LqUFBGjwG96BWQFp18IfQEBfuBEkas7
klSHj2kXpX/mESvexgqCqScwYPGhFeDhzFKW9ZorQccJqNrItc6UM1c8aiDf2b/4
93ppyimMRCfnJMFnIf/AB/4DjvDEJd2U7YwnTng/3AG+Jj2o7ucXDRYEiXSr3oj8
pcM77LzVESRrCBu71V+I9twcKLipUPkspTsVGOXMX5fcA6tiA7lgiLz062ScJCCO
ZJ2zXFKQDOTSSBsLsW/kWMv3ALp1VXFqrldGZIluMW6jqCh94EvSTsFMWw6fr+Mq
9xoavULztl9E/AOxFN/4bjbVIXSsEJvkjiEipAvpOBcAX4gnbCHcX2OzC8Dzwwal
AxAJMQtk9+P9X2RpsSC/kEaD0XgwWbU9vLjj91NmkWwuRXJa2zjFeFXkeRZc7/tT
J0qt7IpbOId2vlQiMbDo3zdRm1HFBjZMEN3M0rnLc4jyDgvKsMLqjklLVD7Q3SvR
SYy9gCpR4SyK4G3V+q5gl+9UU/Dg41OWfWXh0Da1MFpS0sbyGNWcgrteEi52jfvV
BB1CZPhWwGh9mx54PNaT/bXAjYRcfLxI/3Jx0SYZy+uLex9aVWKLUMYHUO6iFnJy
wWprf/YFZ98a9ilNDTcFPrVo3uYlwcFjhbexKVdSQn6iRz4Uc2QwT4vh/j2tPdSo
RGtKE3EPRk4TGHdyqcuaGn0DxpcGvlABycQHQLL52QSk6eWRBOor2zRYc4ePMpwW
jdk6ZxDSvloySpmamUDhsnuNe5MtAPx4sqCPSQMyL4kEQ6gProIA25m/T/fyH7CF
zpNOZxDGXiN49ekyMvWpIPZPdkIu9tLBA3mQ6Tfl3kdzck4B/HB3ViVNgyfE5YYE
0kTYU+gztZrZAYCq70YQFY9CZNUVgEz9hSi0mIH70uTpGAyzmLE9tTcyFEUvqkHM
/3gs2aHnjtM3f6TbHKMHB5AW0SHmKTCwbWNuvEBfeHaQ5UhXhBjHSc4W94jklm22
/D73tZC97QWpItmJWqEy3DZffhFuMnqF4cTN4OtcNxJmHcVPWgezX+PedHPZ3RFH
ZSDx2HTqTyuntbvGw9DXiaKkEvSJ/cHBufOzEDhJ+ggtytKtWwowVIefE7on0yWU
p9TM9U60REwAbo3PscPscDicHoO9pVpV2YnBUpr1txhvZPdiu6qB/EI4rget3t9Z
aS6KVKd84sHO5EJLgmKBt1vDyj5+4HpCpxeR3pkhwMwWy8XXplJpZkTTSh/TVAyr
pLN9iO6lJJNjJs22N3nKkucZVzVEuHYla3nMAR0Pvorhf3OU98RL1V7Bw8lzfzMZ
zOWF3o7tmy8ehhzon3xeyZg5n8CaIlBKkDAEo0TLTaXPuJARvnlnPM9pM7izg4SQ
PL5TOwMgFvH1KWcHOOjYx6CXdidPmgmHMD1KRX8pxYe7TlbR0wL7OD3OUfNQunHx
dsFVjXu17yrBo5Aus8zHoyK+cJa1hJWxVkdJTdC+wMf3TK2iFr3crUrsU17hNxGK
WVNpRaBpOwcegL8Db3H/FJWeQWO3VM5EU0XtlpnyqF2enzb1uBNI3Pdscn/SczBu
oma22bSEyn/C7yAg2Hubxk6IxxOShnIsJHaTUDvamMDhXHmmgRPRX7KciRSv8Hxk
Oo4251tUDd+h4qcjQbBvi3NmmlWA0+/qRKX2D0HcBp87EsvNGHV9c9IjlaDgzq1k
rJCbssmYrlY3ZmdqJQ3Pku7GT2a6K1jpJ8tc8H8r1jzu2E7kJYu0CrLlnRLXVrUR
aGYeeWeExrlXwTAGEpI64YV78lUuNQaKuu3L3VeRYi+fZtgHV8dxA10P81h2CDUn
liTWgFfhbuwlduw+jqBGORzNioYzWP6Urx3l6ZmcG6JIYMUObW2H+MercFb0SMwa
RaAVjgUPSydvy8SynxsZKME4Px1x9gSaNWuKMKNR907Ynk+vMxWvb0d4dXNXfRh9
C4Zw0qiGH/qrFBbKflFIBEzYoBUvtUsQbbYI9gdQ0hmCueBhAEZ/6ooB/RBC9lWm
4rV681kKJ3pFQI788HsNoZ/ktgV7acd05LGVfkMalOOCWRQHzbSX5nFngPqp17gp
2nocQwI1eGShUOdeVhHlOmPGVo7Tj6Oqpbb5tqd+uDBhaS78RhmC8Ji9ShWUKlNL
McSZRLVyVRJuEMZJPS6Oqct4DmOnYrqrul1KRmDqNMevnScx+811QiKeugrek1HP
rFYWpL2PIq+cZFtxf/tV9tQCqzW0Atnj/4OoTyBg64Vgx101Lhs9kBBATbReWpu3
QhWi4t+DwPq5HO2hZ953InV1rJ8/Du+0nlkBMAV0c9XkLv54g090fdLFUyjaMyiU
ZyiC9bhO3r35WJVbyMzMW5aKiqTImCDvbVbu0CKl/05QcZDWNGBXnVOD8eoQ3jf4
6YOJ7gFxsrYetPx7NfwAtZRwCuG3v6v4NcCg7bK6fqqqBX5UJRUrd9D4q1FSIm9U
5psxxdtUCjaPTse48NndTTseVxyeCWMIIpAwp/etIm/j7piaeWjyE8feVQnT5yzw
sScQQaCW3He3qf342OHX0l8vHyIy+BSrBljHOptm9MwP1Uxlr/47iLovoz99bM/4
o3IRgT//SA3jUb6wxDheBzwb+dQD0VUegQZ3Rhym8hcwD3muHcXF7gVCJ++6S/ui
X7wRP0wfOck59R9orf9/rbyMtAHtZidZTGDvyaEDd3242wPdlCmmvJuXYT5FyspG
ywiIcqS0jFB1n2omPgrDQyDW+0eIuyjenCqtDwrPfk8rC7O/gpHj7qgU4PmZQeOc
nSUdmoTj0bGFlJWAgJDMYjBvPmMNSn7T5zJ8ahMXLZlCrqvVjskT/8kyTCk+tz6K
b1ezupKvxR3NSiZc43vvC/5W0u8bE452NGrle2aOlb/ZTI7SaqWkQmOt1rbr4E+b
XfTw4KA4VPSoWqXe6GaNdaw/1KtS3d7W/FWahhtO16yEdlMb+IAKRk0QuVfhPFCg
gCucsVgodODWJ3186YyyYmEwfG+MI70pUndWBRaS5tfl+WCx/oaw6sdTw1WOUQQP
vyjcdJJH4gWJSoOsBFL35tSobBUtkH/1jBTpZbtunq0lG5MEpTY0o6gq7ROdlD4C
FsfCcFzvCo7ornxHDsjK9Qz690nuaPEmGmyVdb74OJiigBkKm08h27MeFjv/RMy1
XkfJz6YldYfdd4fWGPL5pRPYForeYthCVvGapgCc6Wa4Y8A1EDlc2BwJ/N4ljEuU
yJq/EX6pr8C3QwMPTcM79BksXaqkSqOuSpojNKl8wLe+Vt1AnfHvQRDxSFwuNoMJ
gMIXa/jRVOyQcTVwrshe8W9Fb6J8Y4xFvCFF7hewnduiVsakCEOaHYJfCC9/O1OS
HHI+eWRWGp2DraymrAVeUBY3F74Zfw3by95p8EKKm6JrEdg80TF0ZAiC+Xilrq+p
F4Ptmujwj5vmuOPMqjss1Oyk9hxR8GZP3gIcVO1Mw+CMU0VH4pHWYjrwni8P13lU
TnPch7NYh16mjcwnlgvSsHOf/H+haZs/vNHGNGkv3oOliGGhlE6SAvKOZDCLbcrg
jnO1ePhvx/8G9eWg04rKdYDbgy3FC0ZU5TDLmsX0X/x+Xry8afnZd43wChwmoUCd
G+s66nO3f+LDJJBe0PPgcEoFyS859nLGsDcrrjqa3SWxMAa9n+7ZCNQYXVyiwZot
C6t5X4EfWjv5Q2xKlRAg/HioVSfY1ZP3FdtqN0IN3XlbGkQoKw3g5D5oVQGD5cFd
e8R4v1mAt2+BrggeRoutLymDxoCM1eixMdcyJXlom/wJePhBd+AgzNaC5fDHvaXK
hpKt5SQNwBQqUIVR6SDEBMALDhO9xwxHJfIxU/mw3TxiBYlECVxr9E8FAGXv2S1I
ghSzgvu4f49CECcKgIY9Jjsn07ghD7FKE0GMTHAsfLJ1AKhYvy89Z+df3QjDnntA
jFe4/U6gg2FdVr2NoxVbesmHxSlRqhcErNO8CByV40gwY4eM2kkIItgZmcsLt1dV
hhx55I5PmltyWXuLfPoSrCX6WsX0bs1Jn/c63XJoxIp2jhzWomvmM3y7lyAVD609
+52CH+H2jtDGjoBeKppuo22w3MQVCCQnl1wlZGPeR2VI15s9cUVM17HZl1QtlzfA
wnHeybXem1Kv3YhSef0WctYlr4PgDQ7xLpjaKO7WJLFF2BOGgn0sM2x4kk5DpXqs
5/Z9NTOQ05R9YXVzGbI3l1l9A5bwt9FyBLay1dWU0hmJi8GhDgbrcmJJuqml1kSK
cm4GDHW7lBXepG2auljILpfjPevd38g8f0j+hkWyy645H5NL+vmBeDPSqcH2MhLv
0x9Lwpu+isNX4qH0KR69sExQjIBPC/ADlN/zR+1BOTNwbSFDbHA358Qvxp5PLt08
Tz7XUNTXVcKdycp8J96GPK9+xmL7Pk4qZuvdE7w7aMWjpWEO6+r+gsFHOIpb1YqK
HK3K1wSG23DfaYocqN3qyhfT7C0txNnjnQ2LxovgOP0hsQE31+nJVtA5MQY7kykH
OATu2ZkXPiFtQBK63kt3qf+Ndddy2AB92TemK7EQbZ9qUz7tZKOUDsN2rUPSD3wx
PHj9SFAJGefuh+rZrzK8Gpehq8EvNNjXtdjumSQMC1TEDGB0swM3fsqFl/O1siLr
G5LTvYGJgBQk+9FF/Oy+mQ==
//pragma protect end_data_block
//pragma protect digest_block
aZHFXReo0kzzVTViexaiuiEAhoA=
//pragma protect end_digest_block
//pragma protect end_protected
