// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p9CCY8u6/7zkRPfaIZFeCwJSjqXq0vV995qqofy/pvNFcfE3rXbMeW5Y+n3v
bBJhCCiy/UW2fz0L5aipFl9+eB+fbW8Ela0L6ltVdGSHKx34qBHC7UcYLGmA
kmLMU6sUBctKU6m+Ix1cFafTzY5T7r1HXv2CqCCa5C1jlQ5rJgxrx8MFdQSR
hY7Giz2YkwwlWJQAimwNaNHqXb6rTYGTmNoPlCu4O10J53/rKDjnJZYWB3ne
6gUepGd/t8uu8YbU125BmkfhFEyr4er6lnsx/WKoTuhdm/wRU9Y+DbLpNaC/
y3nVQMwVY/tiAkB/zIZ5GiQgRNOl5prZYrHgFauRlg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DTYEHEEm9OSwXIZqxXSH31BYNg2mwDmf2V98tuLB0NkWZS5PNtVpxsVaZQ5o
s9nD6L0lYK/dqOOjCU7KQzr/aN/c01tJK4UrK20k4KrcMWLoaIAC1gMMVA0w
EF6ELcCUlHuFuakKxz86aMMXS3UuiHAteobh3t33LBLAl2F6elYNXWzRzkMD
ljrKMZhIs+I+/v5UXX3XMR4GaBaKXWLZocVFHoYd6+YFbvcziO7UfUFxA5Sf
C8nuZCASTDCkurrP1u5HHSDgdQfYNx0DVsHA2oH/ITQM0YkrRcAGo4uOqimY
iSOBY+rr7YKUchbI7WA+zmKjGIKdx3NilGDh8w/pEA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gQssxUMRSCghIZyeDtuM7pqmcc6W1vSoXhyTPgjWQqFSU1tzIFMxKfU4z+4+
dBq+pF4zpovrvZ0CHHeufF28cuICYFPfLG87hYLZfuDMJWlkW2YcwaUtJOS+
OHTbIqU7OAEIxUgyG7fccWVZ+idTcwSt49WTxg2XiGf+YPZedahI20sVsSAa
S3cJwT9Wq4Vm/42R0m+UE/fycJPoVkTVI0ytofZGD9hc8kWt1Xzj7dFNgKOo
PxdUuTcLCtWNjUn4a5CLsN/KQzRHEIvt0xVhJEVmnnw5lTYr75C6naagIrht
PK28h1iyGgdIJrngHPKkye6xZoEeYSkyu2egShyFig==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mqTWZ4Cs7fUp45bdrIqX5eX2UsuIj5Yw6YPeZfxIZxtP50TufW265guiNU3P
WZ7/65uCR0/g0NDBO0A7BYz7fillsvsM8zGpjhD91ojMEHxDCGJC2IbSW3Hi
lylD32AMsyYFKpZkBYHS2icCzY0MXYwz/NnGtPw8UDb4ejCpbvY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WrnNliUxE7JHFEBAabn5vEq9NuYKv6E/KovgCRvxG5S4uHvokR2BGX1uSlEv
kJrVV3/C9d6ulVCsnkbsBXjY8k5XyGkA5+aQkobUf0i/A5HI7dScUGDvti3t
RmJx8/qq5SL2DK2a27EGcL7B2f8+96Lief3XUJmpzpCT91RUn5+gLD9B9BtS
au6ilnjnMzXzeYHVRW4/vBCwtdPeypDhFiWxAIrwSxgmhgjJIKYM3Badp5Az
0YI6AIhyNKllGDseVxYcT8Ac7Ts/tADZa95YVl8FRmN5+a8+Mcn1H1tNgv0w
RB+I8RllkduK1MCCG5x8/8XVH0SS5jLj10AklARud+5WDSgKodeLKZ6TcWlH
yIzxoUvRBfx2ZZLSZ2YGLOxE+fhQV47V5XxADqXXFcwZE/n339A5mUA7EyDp
HHQEwsZltJEyehVZIlZZN1oy+hCby2Xo2WdnuVyM/8ae+dsfs7y2L6dO12yZ
lvNNHvvNA1NgRPmVwtnPeIu4+LffMeEc


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eVlogNDg/Pu6Pcru83fO9hl18jV2VxBHR6Z1ds3oGLmLqa1MyR7feDEzMvzt
OU6cFbOTNo6HQH6hAPKHSZx8Yw48t/1FaiJN6R7bqNhcorTxFjxRZb1YCuPP
OTyLKmfFPZDTpBb375laiz0wsujFqUxhetP7t+YRyYyqGestiyg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RoCLib9hMKO9ZviqS622WPeMoFVzo5SQMo4jxUM4bWVHMPonhXGCkc/PAQEM
zLwkJl2sOe4aoVDQ6vR3mLQUm82Y5lKgF169FyOJM1nWW1RnMod+TrcFvjen
wptTgYXkl3OuKyNMSWTut2eV03oo6eMxlJxt3qx9yqPMP7KFKfY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21856)
`pragma protect data_block
GJBBzvFYuhXVx6Gl+0XCv42shkPGKUdPo0rrdVcetIqxxidKkt53Bzl1WsGf
R+wk1QE3Mtb7+WBAfZ1xvzoo/MtaZLmpH/1H4wjLPc59zKnCzoX7UvowlEq+
fYllkUh5EYz6iGjAMgonW63vifDXP68mkBp5Ca4ssMhW70GLNnHOcXRRG5pp
QAl2SJiYW3nejUdL4kDvPCyWSIKCQgvqC8+tJavLGT7Jq5emx7fBaRYDS2LT
DvAT0mAw2bhMjYIFZKYhanf1DXBMtCci4UICmf50i7yNAcMGEQSADW5llxG0
5mdml4M4bojqjB8M0UfyFOwDiCYHTkzLvGuxNMdsm8y9I+9cVZnAW9FTvt4i
UTF++R4KhmRxdOuLyZfZgsSW5M8VY6ldZ/owqMJ1PjAoyOWca/mMhY7+80ZP
XxK9MTTKp7O6fVepDrGheJM4qemmNDV2tlft3Uc4d/EerGa3cCnqB6fmTt+i
uQmDkcSId0biDoLCQnSG7PAVaQmFvtKR2/mceWrh7sODdMC7yOG37qceCaFF
lS8VA/NdN9GzeKSTvlzHewJh8nPJPpsjHUJCwMCxH/pLoLj3R/55kZf12Znm
pd3fe/ubOXDli2vOtb42jDsa7ebRpqHuYQnK1rJjnaP+t6JoDT24zSGqS6pr
fNPJb1IstzmoH2buNXQ6k2RHp/kF7KR7PigEWmq+b0eJo4us9UMa2IAmg4dE
TLtK0au7UWUEyN/py533+6zIxs+K8qqrScZkXLPPArQkBcy+SlK/mR/RyOak
S5atFk62DizqFpLveK6sgh2sMqz8ZrRJDqP3mR5FHqBiduNhH3oEBQqoOidJ
wZo4Fm3oJAyQyfTC8kHyz4C+1PhKMUKqVwsUsWUXiMz+92ZpSjo8H1Y8o3K3
rMgg1z/6dGIAw46/C2Q06jRQcaggjzaGr8Jg6mjTh3x5/cTuzWH5NzPOn+Bd
DFo7YdYvmFKcNkHlE+CNCysCZ5ktY4UhUyT/3c38PWI/PfWhDczTR+Sp9a2C
xemcRncLWnRTwxfAzA570gCIPMk53yG9PN8MdF9B716DvijD+Dn+Cz0M8XOv
mw6ZtOFyAjLgq93zT8E4dDtAz4/G+iqtcFhn2aYspwHErGnHiusKle926yaG
gousR2zX3GxpJyRu0DWnVNmbTyyQy/3xqwM77pHrOIHovbzINYjDljDvRhAK
qqTdVmPqn3GuhBeDcNqbW+uZJaRQz7RVY1ceQjdRRoumEpu7kLvUOrKYufE6
E2q8qeYzOk11vTACMVKxFdT/x4GUW9TjYZFUrTmd6oEhPjYefBa8v4J+BcF0
A7x+iT8E3w9i10mUM85WU9QJpT+THQBx/2jBXp1UVj2V1tyuRAlsX6lNZpJQ
MgjL0B6RH+i5wtIEjn1yYMcDVcDOd2mKkyDKGe79fVht8rU/hQs04f5L4gmN
N210zJVtk+8jYZ/q6ET6QyYS7Gwxd4bj+7eUgYfY/XHKAGJXf9GTNnRzr7p/
mZj4f3meZDKn1Ejxw+2GLTjOFnKR01CRFQqwROBUET18ME65ISICJOv8R5FH
c68h0jOXrDjiEugE3t2WWTK315gW/gOkJcKumr+VixzCQTbltXRECs9QDSYw
EvowHUcwajPUJvsy+tuGXYvEzYLp+unM1ldSnujeMik63D7+Ra6LG7ph70XH
dhAumLOBkAlTTq++R+F9sR6Y7ja91KRKTVpFwQeAUtfUjKpMbmouRw2x49i1
V+TCpHfJLpt0cYsN/oziptfP/is97mOx9Uq5L3pSj9F6wK6j4T577tqoYXxk
QsmTIQJcD2NAWnYqrRXftD3BoXw6vkZcP5UnyVHQJgmxnMXbb2ZjWTyJ0YML
IHw9DdjpSTGJv0vL5OU+8UCebQkpEe7XFy6CHm6gSx5ho5g2ehNa6DbpkvqU
+VxYm+avn4/sc5OzS4W8Hef8EKv2bnqWdpzCJ6H3gQHaups8upZvOvIwM9PT
X9pARymM0esPlhEqotoxFPmrD4eiKafLuAVMs+hdaPC/G/0cYIPwouePbR3H
/OQntH7YnYeAsIKwFdsmdwXXYvCUcijLQnlHHAyni4P310vI4vgdUNJK4eeI
VuMyEs3KtVi3RFGOW+TfeN7DPxxA5haSjYy0oPtIHtgEWLYQgU02Cx3PJ8mr
A96QOZcm5uPpJdd7qCPatEYvBJ7fTYidTIF2qs8HJmlwS1JOKQKnj42ikzKY
DNJfDrDQCbPnaV+Mb4+M/IriV1eF5Q9aeIQEguAvZHHd1V291wHVm7PoguAc
ElVLdppkYefPw1/SyWxizXO7pfEp26qTg82jN4GQZGQkegioEmRr/kHyvMT6
sNqSKhyZQVUJIg+G5RmASQ14kLIX1g+Vcx7D0Pliazpa2T+wY3Ceqiz0hDOD
PTXb9R9XB9YXaVVmjVvms7bxj6+LztdhG98u8XLn53x3DL+3ttcuCVLG6qxF
zvCCHN4LdWA0SovjjlNj+euiE9+7DD5q0kIIi5Aav25EkBYTIIzIej0pny5/
oChiNhxli8L4uPXgFrkwU3QjJqXhfIfkKA51JKE19wmzw1HwJM+1pQbvzTXU
e9Wq2rqoZon2ORAl6JbL8lIaq/wvXYZItXBxh9wpCTA0uoL/HnhZAES8S4H7
SZgsYGuWsvAZi7B607nf92twxBbTI7Nl6lQDZbil1rtnu3NYst0Mc1A6pj1H
j2alZJvqZO4KAl1alZ4RshHRlg+Y72r7NOGG18sT3mh/fmIW1Eqa5Y21+P2Q
JQgQlVA+qwhPAtLo8qVm0PK4PEI/Oo7esZE+J1dBupxRosLRumDem7PxVvea
8usLc5HQEBi2QeCRGJLT4BjQn+GLvBYLnb/AUcI7dudSNLZeHqIUE4vv8EBv
9QZfsfjftEkhAM8tk4nA1J0OE3kQph+oc+J/L/mnhFDqW2FYGCve1PrMn4RY
r8eKI6DRl8DTl0Fjsw6e8cGJd1mB7c1xil+ZHJAdRiM+kjGjYocYZTtevWBP
wNFFhiaVCFSp0K4RzjAAZ0NAp54RqgGSripf2BoURn4vJefFLtoHYrtrPz0Y
MbyHoOtPCbARu9phuse1BQCZICcFKv8E1HRJ2ZPUnhLIyGqRDXTWKyyihqFE
52NaS0V9gc2aZRYkZ9z2XmVbw9CYy4CnnKn7YTKv6RkvcVjts46hxTJss7Z/
dIUzSr3P3EnmUDVti6Hk52x59WA8qCGBRwxx6mvG96mYNFUI2kpMT46TXdej
vjGek1FzabD9kq94mlPOAkuZBdu10Zt5Py+2ypIsGBUY66DlYNqmTmTlo4ri
jgrWdZlJPL5JHWqt4YOLNI86Z8Ln3oCpRlXsbHIH5K1aNnoTdjzoddtWZvT1
g9Pp+EJKyCprtz31PJuBhD6XHZpVcZtBuKAwXSLbqHEX732a9omG49bZdO2c
j+q196YpyRk+ZKfjVopq7I8INjV//CDhsSGw/h8RR2kUsrxHQGiC/qk24X+N
XqUMidKIJRrpupPLHJbk/rD9rtj5u1A+iKajmWY/sVoz5dUV9yN0QC+FFrbT
DCoYHCNMh+vbPH2MFgn1FMHSc0hcVVGDRTBtU7XTkmtYjcvM1hcD4MLsWR4t
ncYSUcR2bxcmNAl+hQWNK6RtafMpFWGQwqvn0HnEtg3PApq4+oCnikeMsBZQ
tI6DJ3lTFEy4SUbSSyoVgKPtVWbRmbWoIclqZhsBkhF8oH4Mdysjd73TGlq7
yzYIPPJbsajOtLP39x3WHKwGOqAYlPze/N868WpZ528C1asJ1XJA3yRB7b7d
6yc/0UZsGrTnGTz8qRrcdyphilGUa/qiATttSIigWe6ZJeGv4093zjkvxmBq
jjOG4H9kPq2nNhZqx+ss8eKlgYF+iiF9qBag8FyhXIvFV+gPr+chs2ld329K
q1LxMbYNZbIgzc6Biwhl+8h7mQ5fA/LVped4muMKeY8dzMzsdX0TevOWADjr
Z5ndWe7fpfD8bw9HA/5ZFgFNpQ+53cXX3qwMKZBcQJSeIlYaFPqgMEhDm0kE
JerTJPX/OhUOBQFM+iAn1YODgmmi0/kcPtoA4yb8zLR7W/SKdcHGxA3fi39F
9YPtAmaDPsK/mGJwTPRp4Ki6TibwFn+w9reXA/Q0GJmfwR35n/YcQZGjQfPX
YKvNyrKyVYd31uWAWoJLa1O+ScaKjcMbzA+6S5dVC7n0rsbu114plP5tiU1c
88Ywv1is0rJ9qX2kBWlxy/KXtSK5zj2Fh/1h/QMe2CG3rw+rOExLlrc3xmOn
2Zlhw3hJBsnS37aey/v7THlqct8be+jwcUiyc4va6962ZP0sQOhhDR3b1bdq
cox6fdB54Kyo7gq7dLIZE08uJFCtufCBsnGg0fCCIZRP4hGO8SYf9+pRbWI5
EVcHgQhiDQvqYYjut2Gd9oH/HR2IpfIhJltrckQUwku7O3c5c2vPNMt4MEAB
wfvPB1R21pjjW2ygd2btaESba870giD6ty0Fz8JvuTZRSDYfWip8SiCDfE7k
X61FTb3jIEa7O0ArO3DEYnrfpxzH6sAch7ghnJ7yLH5M8UpV01Iph6iRKK+u
mZLVi7clRSW0MylKLYgTNPFsdF3Qt6MxJCP59FbEPOCWPxDxor84uwb/nx+0
LEycfMY/axB1/T7s19NLJJXe5svvd2MEz8sWye/Dujkv58xySOiD+AQSJAVs
7VhtSN3pTtmx4R+vRy5htN2u2k3hGRilaDzqeORHjVd/0dMsvRUppX1ez85t
wkbRX2YCBZKVxLHKm0sKbij8oY8RoYOKmmob2dynhFeGOmXpvNT6xRIIstQ4
MNniMbv5xXhom05Qs3nE1fETn6WePD7UBCyIMshYCHdkpcOoppluDJ8B8Kne
6as9c2Lgr5prU5Jn7e27JkenC/Vf8ujfS4J+q5sBcjrduMk0WlFR4kyys4Ds
lWBhzelGZ5+iEpDKHSol6K4eBOn/S2AUnbQIA1VICJPRtIC2JOE3wyMKbhtv
yDUhfi+Kit9uCft9IlF6wbTwQ1i6gHumayAWDGutTzoNSRHsCN1zWZ39CT3I
0oxpR32IE3H6bDV4GTvL0+O4WRSn5ZWFr772iTpfMMEpx/gHBAZxGLB4cu55
PIIZaD7lktD+3hMbh+5FwNjFrtKQF5D8Cqy6rrTpDhCqtNjVQLHhW4RJZaU0
A07LemaPC8Db1ghjhkKiaqP3lUnNngyxm/Dmp8+Tyd/7YGoq3+zptw/N7Crn
B0ZHKnhGC6lkrCDxu23iDGbUNe0yxyJeHuDI73OsorI242F+c+HBC2H24X3p
TTPNT+4HAwpT+YMo26ZVJAWkoZY8ZgD2xIS8yO1+0jWZMjrp3Yf7sKmU7Vbf
1aOj2pxu0TMtDSbubjnbYxeJUWmhivB8q5Gmg731uqXecnv+JPADoEFL1RGP
Lh7YeGykRt3aQaW6mERqsxlSJwTSjA5lFfwdwLHD4XCGGkyNSYRiQjIhbfSJ
Y1B7rp9Qsb4X4bk2nmJvv7aTiS0lKt2Qb7Xdj3bEbZDmC+TAf81A/VpLepuM
gnJOGZf7Ntr5328RPbD1YI99oNpwQhFZzlo+xynnInuqTn/RM2ir2By7LvqR
T8GOf/KnptYOOLpR0FrFwunX+cgNYolZhYCdj3gsp/HKRYbVaB1heoNpm/4Q
uoH6X+TykZ29fwlJsp9BZ2JnISdPh20aKbLKNxIOh++Dm1yl/7cH3+LZMJsq
vzzxDpc2ZNHKsMjVylg8O5vwXVs4lWCewXROq5cmgind1+vlvK6z99m2YYe4
H2SfBmYg8zMJi6vBrCGlUyEz3RgS6/LH4nyae2uEhhRsGe5buLtVGK32L9dG
/cZb7T2lJ9BxtIzyHS7hIgjAXJiof5m1JMlOOFrxe0/aym1N4FIbK/KWeik7
k+YtufFSuT+hkEUEESEXpTicHxupEdhTYZa1AQmdWyQDPCxf+f7OqtCuqf+w
OkIQCFnf6z6t3Tsyvjsn76rnrNMsJ3TRypfLj9QmvHTKzg+WtN3+nmB7JxUD
ISdHxCnrvww+GscV7oD92p4vmVcKG2WfnlQ++6tYAE/mGGSSOrtqkE2t7Bge
Mt3SLzgC3GSD4h6/J+aE/CuGC/0pQkwcsCSgENBjDv8ryKgJqDxb7VHgPSSS
8j/v5uPWG53hl4WDEV16uAgYpDS0KSR88GMQ7O/brdT4EXAI9XYm+gEBBG72
AMzJAFKOElIbUy9B3smDMrWGLCowVyzur+ymra9CRiZL6VcVlj5Ty7uofSXw
eqVFHl9veHr8Yb2gl5gPuFuUE3HF6P5zZW1SjK+Sd2gosp+/pJj3ZVRvNBiu
6WxpQRUiP02ckR5LsMY6L1oX4WC44HuQqfSUdJfA7gK+UM9rBDuCP9B7E18a
uYPngh0iUNYRIOXYqMMFcrH0v+1VaJBSatxHXEEB7Ha5LY9Y0g+EZSdYF/KU
vEq/TmEmjYIKu7AVN//QmnoYvD1C77KoGVxpjKHfnTlsob1bO21yrAiVcEDF
iF8Ql4UvbWj554lZTAaaji504SJj0Ofh9TtNaSGstE9giPnGB8xd+lxfumXr
Z87/bwrwr3L/FQomzdSZ17Ooa8DQWfCfNd56EUteWA52oxI60H+9R/xSVxbc
DbrJZeVuoGqNkennnn9rGTqx1nZ0xxJo5kuprnEzgSEqasqd7/UMW8rFRSCz
IQjRH7XSwcjktY0sd0uCQBPD76QU3A0eXzmnnaVqjL9T9NnYh2a6yPDvkQxJ
x2v+2pF0/aD9raw1cLWzhi1qbNb6uOEj9pOs2fhDwzgFKPRXyaze3ep6sCMS
T4KYsVXKMRveonhCgqYVZ9ZLvrOtbUBtDniMSxnCURGQ7mKd1x5BHcCVYH/7
a9jdefIpmLiyZjA5odTsya143iSTKlfWknNNABqtpucd90RBhZTDeTfo/AYI
foqLEIPN6JOwqK9FsF0OtoNYl4P7PKIvz+KrmR7aRK/gVT0dqJuEhTvcx8Vq
P22j1KMmKXKBhFIWUVrRKZdeAqPDHibTTKF86HRIcRRhkEB1wUhSct10NyS8
0++rhQCW8WHcNTdv4joDrvkreIiS5IXTCzIarfSjfOQxVFJHXOY8zPXh7/oI
J4jZEFlJKINMiqnGdwVZ3FFnsn8aOKAlM3P6jB+JkeIRKGpbWh2sxcXoGDlf
SVaQdjfBIFTUevGhvCK5ljq8vANTu1+mlL/NCSB0r5J33k4hNorGvzV2sq9X
7BCOTOFiqB2VnnfmXhumECBmQGOz0vzdxjXyPwC8Z5geR+3nRmMxwjo+nIEc
S3qJwMKLEYiJUuGyCUHlJDnmqqFKtpIwBXOcsVBByv1gKSnm9GBHhA7Z1vF+
9d9NOx15qFYk/PdkxqYvrBU7Axi3SuYRMLkgVNFXhim9mOH6/ZTgye3yjehB
AHVg+jINkf5xBQqyzY5rrxASLGV6ooFYIY04HVtvl6rBywPwiNcL0CD30H0C
2E43lpYEWGQi6LCYR17jDzmrwNT+9wteIP3wT5nN12ODNJc4yno6o0ae8ZbR
RSUyhW26MNaE0LT9tB8I8xyw2PuPklcAdnmgO/crkNH7PP//Dzm4V7LBWXFi
tqaEj9mBru8RIWGkc+n/gbv1PUlYuRXfXWXcjI0/a5Zaf+gBraYKhiH+Mwiz
UgRvjzpC/mla6iiMxqMRZZ3pFFlKewEOCovsFa4g6CuY6uZ52OiQsGf/fdmC
rEC4lbLZOoHgxcsclnD0dTabylGInk0h0dHbhBYq8iE1dYcKuZ03S6gw65Sz
AwUPVdu/qmLM4MQx/yP8eYkqwJV+Ymyt9Fz7AJov8ws1Lh1aS1zKexoYKDQd
EHE4b9L0m885MOlllgWLRtCQBhfsdcupt71Ropt1sOq1sH+zBiwClQHm+WrU
0cKbSQVMk8uiZguNIz6dTCmQuuG2lBFswm6J/WrUCu6/NdX5Dz1R7rRMyD7R
eRDygfkMgJmSeeBMf5bQeqjv1T76Jk3DkBfulcC4Fw+5pNgITvHHAazVJAbH
/oUk46ZN+QTxv3UvfwQCbiyFXAGTyQkwSkVkzpYvwbEVVGEU1VV2wRESz3AV
d7dUAGmjgCNgGWVpJy2zC+v5IVjA4FARGd5dYYzzvlzElzWd4K2pSc4eITlj
6n+LoHkt63TZ4hb4SyD7O6B3o/421VHyjB8R4SjXQUFX49xgDxXgsrZonM+5
FSIEBS/p3EHQAyNiJs8w/puiveFLacIrj2Am/u+Pe7f8i/6lB/YuvtGTAdtt
wKweOBcSPpnpkfpa+Zu21vUNBQ8xRoRYn4gvBH4qCP9wZiFoatElg92d5MvH
ywdLCpMhPUUSkebmnV0b0Autatl+NN85eZ3mtU4q40AlRDdX53phPfzxExA7
guWbuQ8XLrFCckrZ59JNmcGMgJHdVi1j15bRWVGiFc0Vgz24ytOmVIuC66qJ
E86n9AjQrB9/JZTbdO5nGfNAsLeDWZHqJ95LeOvCzwn7rTlQswk7IhrmX8eo
AFZv0I+thiw6r/LJFtv2SbNtH3DGdLjIOh6FsSdhp/BWqugwuDDi/y8JvJKy
CNj99TzZkPh0ARbPCxAWI3KCCxfry9qso8AiPtqmI3WraIoHX+Dk5GijNq1m
rEBT5y4Sav3yLysbYTG5lISL1STdhu5onDIbHOvg7QhVKNEWjqUb6ORjTDbG
o4inBV11Q9SoHxYguCoatMDOJZT0UWSDZPQ3Pli82pY58bjxFlyOBVKN4tTp
wYZ2opqqUktorAkQOjxlW8Z1hQdfesrUURecWrLMg5OFcAzdWt059NsaGc2q
QaH9H1YFua4JkFd5cAj4iSwe0joWQnpQM90Y8V//mNbrS9+5yunaGHeDcHJv
om361eEuMRbCvpzOPJIVWZlt4HeAFpOCJEb+MDD6kPqXSacY9j1VwXW9Dt/S
CTzHwyrkjbNF6z9Tn5T+rervyVtKB2AEInd5QHm6pta5l07a96mxTfxUMRVj
esofIxuTM67Gyazcus4aa74nSLrmGwXV2q0eMfv5myOuyZVRrnCbUn3gP7Qj
ra5qqN7QsjfUTwUBzcbUQAh1cqf9/PFC6/KcAp49GlJFTd8pD42Gd8dkXZD/
pXfeSZGfd3tJRGpqCUW8J/SBzlYUrqUXPg7qncEdk784JikVqLSs92xqfla3
/mtBU6ONLUh2NcVjX3/q0XpT/qwbCq7Xxybk7k97W+gHb+Labv4UyQT31yLO
iuM7SdsPBM3JRTo+MEWvEDCChqN+DL2RUUtx4gOtWAhJkoKW4FMpRd2SjoKU
lK1FDiuw2lDxY5KnN5cYVDPPtTftBR+3MI3xpupgPXTQBtmlluHX1+FeqVbh
jQ9VCGmSKt2Jp3Ly4Q4/mLeFTbGsl9cgiSLQpI1W00ig4cLsgEGzL33OnA0a
ZHLGXRVTH641cKtPoeF1LAmUq4tDZFv7/xBnZWqMAqPl3u7rKYTfPtWeQ1gH
Kd+fUczvCQtv0vJvshHawm6zOTH4RnP1e1kd5kfxnS4dq03vQaDFyK41OIj3
PNhIBBjIb7hoWpAZWU/FSz6oSIFg6IVSGuqXcLkEQOixzDDwkazedAKaDzrV
oSSHFSC8DWmMcbuHfP4VtrpyOMs5JxxzlSUJAKdsyBjwJ1X6NKbBkUzdo3gf
tdJjQID9ERJX39tnggql5FSZ9CX8EnuRBAE4BMi/9mgBtEJLkKL3Og9YT4Aj
gG5UQPCJlEQwD8YwGelRyzHRAIflfhpmDY+GQHnruSCns6xwg76UjuX8YzWg
qX8cuAydCdHDHlHyCDd5/FZ/mjp0OICEmwuQNXv8x6xcL8J0DBEEobiXiUH2
unbLTJ3XYYpCxJB4eCSblpxksLTsKYGJQUcl8elcS+qsEpJuNGT9K/6yJE2r
WjKp+LLbIE/TUeNf6Cbf4C+ktsGIsl7EbiOc4QQ7EfF2IR56dmDSFtB18qBr
geN8vgQBkPEBRPilr+uvmMClVQpK0UAUDT+1gn+0dKdkMzjeCnp+RuXMadrr
iJT9MgXX0xkKooOzsCK5+a8HhkvLrvXdfAZjJrkQIlNq3iDy2Soo6Bz7rCop
qBa5CAHZi4Qga5J8tEgjWrlcW2U8LJVZRTi5a9depCU389oCw6M8SloTRo5M
focNJJ2pg6L9eRHAh87GSrIZ12L/0bh1fWfxzJCVKv1In3lPjwI88Rp1C0z1
L/Bl9+FYKSnWt03VA4YYow5ZVzaBQgWGC950ioCLp1jlPW/hJFJefz3uHuIA
n/Lm1HsksqI7lxfMspZklBeAcxhTheibc4W227rXQjA2yNNW6iVgRCTwPbgS
kp5iC4wT4Jweqllmn1t6Oke7rTGJUAfnzQFF0QcQn85QfM1j6isSdS4D9ANS
EEJq0qIqItCrWnq/EgsLOhNwNEWRq9y8BhoewNVqZL8laJCM91fgTVCsLEFd
zkFYO++b/ejn2kp7/PS2xNrrM2LBMcSL/UPfuWR819I7ivpW5cUYOB/dCstU
ys2zl3viuiyft8gpC6h5NIbvZ3kt1yuTxXuGNYuszVaV47KvL9XE99LMgLVT
oEksKxzr8KqHMCTQilremDuhZn/H5VmwvoIPiCBz5x/L8zPnXM7EvBF9kuXQ
QzwRFj4E/cESlsqdK0C1/1ilbXpGvUvWyLzX7mIMX07p+EXCTZav2ermapyK
v1PYbbh35GVQ37gJRRpu8n+cXq1wZCCOQXKT0oqqJ3ZbVaQmTmrAwacBnNGW
JFRfeTAUW1IXw3sxOlU/uSXoj0L+AGTGeXRrklHUz7LVF0fCHTZ4VNYo24ET
nwks1jZ+RazVAbvPUiKoIjK1c9cxW7e12XSCJqPrh5lOpIfbdNQi3vqFV2mC
8sLp/efVx12c2kV6IjUidZShTmTr5rsC6JxtsaIOSn7vOJecDqbyL8S3euEQ
1uKyt0T3p1aquKOw4/SCuuvG5vp/PVznBlWRAazdpqWNM1oQNStxgrf9n/Og
0GbzgDhfDrm7lwuQ95OpYNZRqvQBC9DLO4p6Zj3OsGgypil/bTJFs/Wh4Iry
YPutvSyvyZbsxANn130s0i/pMI6L22jIQM1GLnIIeFoleC+aNHKTXliRQ8c4
AVfkxG+Vf05do92NyL/JnPCJwDetwf5t54A4fywQaPOXCIRGiw996GIdheBa
llw4jm1a3JYiOk/29zerq09wHk4ky9QUVV55r0zCF3ddMQrrVq+hsQq0hw+Y
YJbN+m/Sc/1BCTCcebyoD/F3EDbj7MVYrLisla1KvaVw9lr5eYcdHOJHCN1x
mNC9Y5paIvk+DPQU0gUnAtnsZVqrsH9CcNJvO2NM1Qtgn4P2oAlw5Kic926u
D7tcbCaPlAxShiXasm6eyGJCQC3Ay4VSfx7Wiv38WA5ihQleKtf++Ez/oruJ
tcYLkm98Mm/reb2FSanfN+AQjhBZL/zmqD7Rf9Ws4VZ/fWbVKgbfvIxs65Ty
DqDZtfmnwIZ/6u3KRtkyIHUYwwCB5n6eEHvGwicJMNbofuAt4i38oRrt113Y
gozeRkNh2vOmoypK3QIuC/RdrY03KuWdaKaMh6KLi52Jp3tJ1b67/q9p2Q8+
E9F5P0h0tnLLfeKWaDNWs+juXCoT5v+6Fi8WzRPP3Ic59lFRxAJq5q37tZMe
x7XA1tyzXdK5r4ZBMtIUiK0lehH98654JY90+bElBgtwfIhONoC+Z1TLCbX9
VVkgci2Yfnxhe8aF5J6jxYNDW8nPTe415S1fjb2BpBXYk6TYo5+Q2HwtmBG1
4p2vI3+5kRPnOZu6OaG4DQMPV/LWkkRfVYqOVATl3UGo6tb7xOqehbYKSV6c
wgA3hNfGVLepaOgA6HfL4Xe3vBsb/+lBdhWqzvXkNdwwc7DbP0zbyc6lwk39
hj63UKHuztSc37E6gDEtALqLkcJG13VhImLIMr8dAVsm5vZMCND6nhR+C3D2
t4BWA82N1JK3ik6ZE8D32W15cQBnCfhi8J668uw7pRp8pew5hfriJOfhmjip
FJnalbDFnHf9NGI3ZstYv+f5pS/O9Cg7+dJeXikY/O+BQfI70m/dDq5Nm5sL
eLHgwhwgkSLfInxp2vLjStFecFar/MeQNCvp2sqwx71IGBkIwQ+FU4JBZgKw
VCV6oZkeFgxPacwsOseZliClfm2cZQK62bnNR1zxb+eLn5mQ/Nth0XtrBe11
uNkbHFUk6ZJnsHeXwtW2i7aie4vr1c7kU0aPYA1YySKXDgsyqc1CGuppGa1c
loalM/38wWa+jf7LCOhOvduBseSTVBrj/XyZESzq9NV1l9XFXfNHPvP3GUFV
KTsnl6JBi654vPzU/uacBJz8ww7wNTelwV+WhtLDLGCM8iOI5PIZR+c17yQQ
SueGtHMvDNXvGI44b97eXpKIcazTQ/rf5dSGCEpl+QciX4rOHMJBityi87b9
5oKOmR5RcnS3/OEpfeUJ21pGth+kBeJTxxaTxopD5ZYf0oGv93MPWXOBJV1q
L2tGkrQvu31dIwEIb9NIRGSCTOkdrH2HMYBaFGLkrxe5YE2mFqFyxX9F40r1
KdXUe+3yNvSaJ1AsvkbR83UGBbrLK11LThmzKzTTd4MZFlxLNojK+h/fcLn/
42Zue+COvMdGorHBggu8q5k0jq44FoLks8vpdX0Afp7rNvyNlEa9eyhaP8TQ
i0VpB0sW9AgKVXKcxW+tYNclfPqy8t1m12lXuz1jm0XLTNJTpCFABrx4cCGe
SbEJzKbqoBwxZDmCzzrUEb47qcP1a1nTH/b/7XJJBvj/TK2xhZ+ICBp1VVXo
LPp0rByFHbp0+o+SlHK5fzLa3A3dim2uThCiPxar7qzU4B9ev3VOnqHCEqgn
I5B/A4dGyjvrGF2qGZcMc9Zz4K0NVaRK73RGe9Ww40S9Cj/XdviPPS0Kyh4i
YfYXb0h9njo6icyNIHqMKpTAVVjzvKBAOE67UOUuHq40J9ENUjorn5LIhdP1
egO5rRC6af1gYLzV7YDo5Bs+YNj9OCDYASK5PrhPqb+mxRR0sf8P8WpFMCww
moQao4ht0dERPsz998ed9gatjpoVKY/qFtiIOU4x8JOiQ1O9m5Piy3bH3Hu1
wiJNixaCw77tIx8Sur80BqVwf63eTch3kDp08J7R2Kr5abPAEmKO8Q6/HigU
nQ52YY76spnleLE2/wo2dLrScrCmXtqaRXnboApcNsbCmTAkYOQlzT7/Drfl
p0Xd7Y9FaI8tDSL7Rx5IJCyR2TWQwCAP7JaLmNAdrKsPMdNRdGbGgQiEaCRT
miji2eTLZRO7SgUBQz8Pz33axw+1cqpBIdZAS3HsfWTwXDAa8wZtyY4iHxte
6V1PKgHnuTN6pPu0bCRGp5Lg4qW6OR8AQnZStY9G8+OMZGJz3e3m4I3WgPVR
AAezc1U/rjzae9TVNf7bvgAEfmF3rgGvnp3+cuNoBOJT3DfI9ozQPuG5VKqL
sIpwXCiXKkwq4WaCOeB4RyDs3AyXxpYYYO4ubPrH5xYRTmksWIbUeHacExVm
z4vWRnVtmbGDnh7OdJ26lsu30gKuwVbPs9gcCrDfCSyB22pWr/jXgGGrCY2W
wyzKj3sH8eDohRSCbOqnicFc+EqjCed8SfW+YSS1JvmKg94SHQv/gWdeekea
h//s6P8KsqWKKTPG4jMTMhDnWommWwAZpE5ubJRStNo/G2U4MIheUASInIkE
DO4oo3PHWDhyMww4qnsOeaJjUoi+dLGcQGrsYHwa0DVBF4Zx+JsH98LqgPH9
E2dv2zI6Kl0U/RdvAEDw5X/ag+Ikn6uVnBBPZAXxhgPiX5SDnracM1XqV9/J
rLKja1zM7qtmITG8Yxd1ioEkCB1tMHy/n3CXbn2YAvHD5chNghLmu/031Qp+
v2p66xIM4+5KNznE4QEeKnN4ZErpAb5/pvUp0mToc49Z13FJjJXVXQcmWMJ9
bedYeJOH8dIuOq0NlhLAjo+F9fFvszGzCIL4i5VuhW3uX+7VNwr9het7NtHI
zGWe4Qo148TtrJSUzvtlNH/YcqMW860lr6TzG+0YA75XzoE1Aht/B/x/Ty4t
s4+l+YZGFK00rY5robXnVuQ1CpHhx5eroJBxZpBFM71Uo5Q847+PHVXnRVlC
I/78eNmrUw82fAdj8xlzYQtVxrgarUoBGr1ynY7p8nitp9VocjPO96X9wgXz
qXJ+dgbCMtndBeAe21/88XSRXVog9u+t28iAJpTnBY/DTQNl+ad/iV8yHXMy
HnUUXc02Gd6slL8mWSqsykor29fUjbJjucPsibrkbxaG/7WZGiy4FqjfclAy
N3vmXSLQYxc4eFLeHyzoODEYwYKdwDXzZPZ91A2Jry/IaPbIgfQXW7NZVeMo
qA7Msf9QsJe50ErH840JPljt6hqbDJlyymZr9Ow6MwiPUJxaIx8fonF9QxKl
dG5yrR93GipbgJ7ex2g4p/OkJqMYZkRCIVlRohS3f+jqg+X99kWWvBlO/vnX
0uFV7NPCUgmgC3/tOwThjPuyNQSC9lDggtpCGkk8+9WzfL/ZdAOi5s29RKFi
+FvUQynmz8npLWEN0kzUsHMdp9uWnLbooXzZDKMV6XXEFNMh3/Fl3DmJVmef
q93AG8F7V7y3zEaYFEHASClHE38+4vuKkCYI7tQJRRbLOQqiUeXOY8S5XKOO
maGnaliRD6l9XhgvzyTvcW7XUslIAgH+rVi2vKjIgRIT2zjsExvw7DEgP5eK
QjmpRHJOK5ZQvAyBMTTEOcWFguuf0bDnNIOG/W31eHWHHQv1kGIrCqIXvs41
0DoeaK61/nMMcO4Ak32lIrnx79yNzQtUFsj+ggg+twdMTdMMM37rWQTpZCUK
zlHRa9uYR+ekOfM6zlUO/oylcQFIArE5aSQlbxKuJKoQPqDIqlUY84R+33R/
/y+GTRxeqADTUr9wcY5j+dHTWZCa5H0eK9w+NJYtAteGz+czeIBsIj+A6QZs
Eu1QdfExugPd28czpACXg4Qjppqa0CMzlfMBPB+O7S/2JSUPzBxp8iv3dmcV
RVrGluQzlxDJUtcqt+TrQOTytrAUW5mzJDfhemWHLlCKI1q6pvS/6Uqi3MWf
ajCbMTSD4x1poU9PiFNtbw5ipQHM+qjuq2r8oVj1r/PptYMUAm3aIdS5rUNB
6EnLS+UdKqOxyqpgLnIIG1Dv5XLP8Guhh45XbUvKmbJ6n2P+1XGEIzcjdj9P
kQ5OKSeduyU0bvh+UcIErdHAgYBxWjWcg1xRtVat6oMAnpMCGDoHrFSCmDtM
3x1MB1ehSJu2KqHesZR026/7//2I+ghrJ+EJeTml5pX1Wa1KnMx+hKCzrsgh
VgoU6pBgHLqJQYfpbSoiHpAZ9/ZyJHtMtHih850TKm1bdDlSSQzsKBS6t9SI
rHryoG7pmIbXRe5FmVUVS1MuzUAqxhEPllvqeGcRVBY3kEKiIW4V8cMUILgd
aR7R3apB0UjE4Zwu+jg/cxADd0u9ho5c8SS8rl00KjBJ4WojYp9Lw2YD3ACI
Vg4VFHt4ODPnX+Aa6aWRBaMFjDhC/sQuOAESspyrXYIVCYi3vIZwyKGs/UmE
NhKBkbFP8bh3+eduNEsAhcpqZ39TizxtB5jZfgJm70ciuI6vIsIFiNPgjFFP
Cak5+QgaFyQr0ZoGEXxBC8msd4OIX8N89YP+lgqmbp3eF+IT6XojVxsvPcbp
kFMMc/nEaiTAOBg40YmRsWf2T5tFA55NWH2OQnfz1jBiTU3PFM9svL+VIB8B
67g5bmRAaxcBaer+jBTK3AgmTrHcP5o/uN+C1wwitOp0Z8UzCkFdO1MBeXY2
gtzURZW3zs25oq88RF1/usYxt3IIzWclaDsD4IINR0iEbYHlGj+Qu2V11a/s
FKAGigwfvW1LF3zFMhXYQswGNdfthI58bwbw+2XPRUM5PdsM5OUEK4jr1LtV
bpgyqXJHAGcpSG4UJAuFnb/IgdL40bkD+vT/Ga4WpMFzPTe9J0aZsfht8LVs
OPKzOUGlriYqsxcGZCR7hPnDAYUJRUNu4UHTpjOaVVIPBsIVVNWS6GZLDfAP
6mYB2d1PmDC+J1OVws8td2IQJ67nzFKwF1kC3eUfS74m3AKt3GjGXIXIKasS
dlakAFu7Cvn8Gu8CLrRuDMz2UG1iHrxmrZGDkdPONQw8jbRa1YHtjsHIMXMn
VoZwWOQxHjEIxOAU3f4V189hiYTy7U4+75vMHHoupquC6d1o7+T+UmlFEKXc
KZ8CNpsCIGgFN/tT1lI4JppCqsucMIgstP7FyR2RxuwIdH3y0oni4U1Uv036
x/yHFLft1dO3sGktUpc/WKdak9o3qaeWT8pzoyRldDYc+gqYoujhu54XTgPE
1YmMu6BgBP/rWnbDPBSFAzKLwX65/HxpcAUUcdN+T8jvvdqgdTWiuES7P+L6
WqARignLcRQN1pJrflgwZ7vhiFEk5l+z18cLVd+n2o+rR5WF/jaI/aQAo0e0
u9WPRrAgmqC8Hq/dF5QtWWDFh8H2sBQtcue9N5ql1VfC1Q59QHVX/6VSKE+q
yD4bhxfqiHT/zfoc45mULgD7LHcBpIbJzkpExNcCsev6FvL4kZRhbNQAp8b8
ue+qdNIyT5/QJtQs9aCwym0SrP8flcFBu42Mj77CIyASqKkPCehy4oKRBfiy
JG3KBUXcY9kdKaHn4GrEQ84Dal/os9/s2flxDgP0Lhl2tFYkKUsWphqid/zo
W1esHgPo1EBg5SjiqJ2USNGU2vWJE2np1Gvg0YEUapzd1Q7ruYTbaLF2odi9
aHn3arPwDcuzLCbAB0DCm0YXmw09GyPcXtNlc5OL1jM700WDxn2X4GIZ2pqh
slgNQQbEGXc+0pHUJL0oiFcRIt97wTp6A1uwGUgJJ9qVftxSg2pBVPCK59z+
2FMVSsh1Jd+Hd1/Q5MUI7hjlkCD2LZ2ajOLlsG/jNhwIkVZGRqJlzglZWNl6
T8Hzl02i+65yTIeRVdDpfRp4/0O5imV2iW9oKv17AxIKINf8KUPmkK+vbxEj
2Npmiju/Gckeay7FR5UTyp/5UlCbn5UTMaiG9a8g8huZMwcBR2/YRCuJ9wKI
Jh6s/xUUM7V24uoTD/6ytz60dBkV94exR/irh/Tofgh9b+f0iiBImqKPAHaV
wq4+dXn6GdwydV8XLtoYGiTrHZ5+zr04q2pjVwwLU1UQH+CQ00K8eNKxqVwE
+ZF0wKNSswhukbfV2MIy5jMkY9WgVdgiiNjiryDnuH7E47D5nJdJSYLSfy2P
YvtRO+rc25fdnTIEBMbZ1vkir3yZS6GTuaUU2vQlSrSWc9PEZqG37LYtbIN6
uIeWeQxzIJruzd/WYfR1OCE7dek/ymgrqYbBb7tZSe1XHDyPlshPP9pMOtIJ
zAn1B0QWDesN/u357CX0EBERZbgADwjOkUvW4T68phJJmzR1/JL+hBe1hrX6
ojJtJTRN/dnY3KIYyfY5StZR5JpHEERK6lf79MZMx+j/7aBAK2X+vQTuKON5
jpSf6w7e6Y3F8S+EuqdLr2l2bPqXEgvpxTGX0/W86qlVt9iVQKQLNOfp3Y7p
8IoeXlPfZtr0wFgcidwlQQrPfhrmSX9xC3HoG66bp9MEZo4bBKuFX3hmDNv8
31tSfwvKCMlpRi/5mVh0i+/vf8isfkHFWH8JGTPr0vdCgXrJffRzcFbLM0Nn
ESNraXQX2r1B29EgCJ9w3sXIaOz2B/vCwjsNbxiXaWxC1BwIN9ys5mBtlDwT
GuZJXTnA1ZMa+C4ELANE9mU+JQD/pXXW/wl/J5GDw3n/hEl/3eBx9K07x6pc
j/nI2Q4cbMSL0H9+H9nldSL467N0X8DEZUpetmioyR2pWl4g4+nMRRsOc457
eeGVsphvR/4t3PZ8t2vgT5GJsNTGYmmcMsFCHeQ3TER1Ke5/tKVIrfBLOhXl
bNl6KN7fPyxEBBtnoljW7WPHsXLyRVJA+QEVqkHlTD0HHHHNQ35AyjiLTytS
axfIPASVIftXJLxJ9e1BTJyonQBhJArl6IUhTFujKt39jfY/J4lGFuJ7zxc+
/+xnlUb8xc0c1IEJ73EoLUCpA8EpPIsBcdeHMtzDFiWBLv969mb5M2QiK/ZU
Nk9k5sU3ZeY/lkfbgFJF6EL638rMSXt098x756ARbe1zUJ/Hwl+jFwtsRFHZ
xhAQbRTRpTSRC0t78tcipQub2bFt9xP/AnprQsffyuZI52YBFAjJK3pAjWkG
ZZV9VRz2htOQU/D6mrKS9zDNjh1U0F111+k/iqN8bHXXQ/Rf+KWqTNO1cFUo
FFFORcYw9OT00Gw1658ZyGQTYJACwbG4TN/KuSlIccLSAVDm/US8pOdi5tqt
F6+9rZd+wJ8HCjw9CxStzQSJ5VwY33KbStMbgehrBXv6aoykWmPLvzgxtc4U
vftiQTtUeKxrmbxNZkhc8wuU7TQmlsRQsTFAcu6uoThhJkysoTOyJDw29Set
6tGveAzXizn+YJ5ukhFcw9bBjPdt+STOOyILB4YEFVI1SZjwZ7O3J4T/mDGH
e9ABgbyY50SP9Q17v07fP6+wYMiZQdZkwTV9Hm7f0A1nbLr6rkFm3SM/HSCJ
X0zFdOGGzV3v/sBHBfpehv50wa7ZJQW4F6op9BrburhayR3Lg/2es5m5l/XO
GOpqrbZODxhjILbzSKrvskrOjXvAoIcFWtk4CBQi5McYPEInINoWMOgzPTgL
LUzrgkz6KZMhjdb6jvHsxtmk82K5dKOaUGd4GJIiMFN3o7CZ+A6Il+bZC6Ye
24bJqJ8OqXf6H3Mve/ltgj49eYaXHckh/d3rjAWXbeyyxTILdxXqSca2RIqF
yyPNPDTFgNUSHZGH9+l284lBFZOLd4DuQYY3aMR9oO3GW+3DH0Rs2XTHdPtE
71QVi3fFo6gBtfQb8A6PC/8MjeeBDdHJnCKFE4vfihp9/SVTOvT+ooqQXk2S
9pKv4kvKkvoT+tYKu1zUrjm1b66rrEsPH5aPgytau36LT7hJv+uTkb/HnlE+
zxU8xh+8K0TgNF7RMoryRtEKCwFtHzc3ae/KH2cG+xD9iPMQj4SYNnw9nxVp
ecOrJ+JN4NpNYu+SmQ4nWRnjdvFBp37CKDB62iHxmA2M1aXbRsqIzcyHujYf
VeS2e5/2votAeoe8h9b093IY6FuuwH54OMJtT2Ld31CmKpLjdmo+n3g5JSTx
CZDmnY113IBV5O1DFV7tdv8K6EvA0dgk1IFt/6u7MaSPAHBRE9FrEkcLN62Y
idrU2njOH51ga/RnZ9sTWGev1EYor4YJG9zzx64Q8tjmvnhGSU98lY/zm+AK
SLQVJE9GkouHrHrXj3xE0OUQqLAJyRS+7pE+ULyFprwK3ZFs81qV+p5bukUD
6SPS1usCQoE783uZc3G3H/TNrDd7jlcx60bSsbP5cYc06v4kF4FayW5hgFZh
bDBvzfqB2rL0/m2sQO2NhgSTA4acXCKLdYSHO1ooZiW+NzFJP7q/K2yj4/RR
K5ttBG4NPqduaXj2FLCtqx0TbWyvzkECmg/o14/oBLb3s0JhUhHnt1yeudfd
+EUinviZSJo1iTMzI5UCuSzWyI/xdlMHie2V4fPrOiNVyMBUs6j3J0NErQAk
K0yqtKbr8dH53pKuJKS9ATDpPXuxWyOOZvHRmopGWwFaygg0iwU0KqeYKDU4
FW4hvHzp0ARIopzm4FnDFd14hoMbzCqF9+6VI5zCVlrnFCyzgcyVNr7LL6pA
/LVOZG/X7tyeP0v/O2QiAnFNpltPBIhd8YaaXXx5prKzcG+pDWqoTCT82T3d
kncvJamgu6lpwJoZuscatWww4RqNaj5Q3pD2Tkyve3lQfJG6cGtisukzQNOp
L/6DIwD4ZEalJZAtU1DVGPCUsmQu8YJLXX8XK/LhXfRIovYdbZ6kKqmSVyv8
BuPToHMF6dKu/xH2Venze+A0202n7E9sMRX8Ibb7uLVcjT+KVsWckusx3HUu
Z+szqzRswHe6S9nZi0Opkid6HsyKyM6x623JROefNjBDz606Ykb1yAj37FIw
o8vgy9I8AaRlCn6S9dgFQQ7CtNRAtNoYHl7cF0Ox5/awbV1wsDTI8MVNB5CI
0zlZNymODinQ/KxP1OHuaV/4DLXOQcqdFVCE3pQTc2FF5OJel2dn+GIImzMF
F1xYIzPnZKeOtN5bFwEYnp2Z+pjN09o+JW8BlUo197nt6jRfb9vAHMB14dxw
39o+JHpbt+QhAR8ThymSdNDEFzP3rt7xMfuRQUAUVO36mnzDaCTMbFCEmD9p
x8h1OB6+YlCRtNV1b8uCHmfr7kCilsvJa3TjW0UBpKGlOPnjK4Q0fkwWLVKz
JUjP/nAvr9XSL4avKdAHuhbilRmvEgbCiXVFNt/96z9f6xPsL3vqAe4FzudU
SOAlPiGhddTaCxa+gmIVnx8U6Ist9NjIavoqMZWrsGptKj5l+KnXm9ppUt1K
pOwLlbksRfpJb+gShCXGPYMLVQiT9v5m4F6g0TtDtwSwZ0+rmQU3ViIccKse
4jdS3fSgbPHrjQN1yikYvivb5f4uswnJSKPVsNZRsJP9+y752M0eIX1ga4Y2
wVaf9Hz+vn2JxuwhgNcUhrY34TEdJITt4e6SVrYfwuPIRgmQit5VzW46JZbS
XdUWQ99UvbZnxBhtnDyK8oCTuZ3o0xMAh16o+jsd7xnpEU8q9Gb5W/gRQME1
5bzQOWVnDVIZlUTL4ofHMa2egAoftmu31A3QcgfwvYzONgBnU3EAo2xnfBuB
va6AU9FQh6EhQqyyzbKmbleqzSA395MD5FMP0unzEidPv83GGjllBJX86lvt
VzLJoUXZgUWcQAP7JO6h5zt4Df2Emg8j4J8zSnVgebNr7sTAy4wWrNaGOIXs
uiAsG6tPLcVlQ3/+UU0cd8awgWHtXIcX+5QW7G88gA2iGZL122i1+WVR0fse
keIN1qkTB6GPwinYHght5jAQjl0UsMX6tRhRZHpfEz+dgkr2p7j7W4VxHs6Z
dYCLfoHl43zDzkYqS+0Lo6vmOVJg1J80XhhXVvxRVRf7AkISYCeOELH5OGL9
/JWgbdD2SQwQVRahTBupufvnst3rHGosmyzGaFlQ69NEuy17/nxN+hABe6J2
16malCITltVoxhcfbAaGD1OgX90Hew/Dabx52pof2cIW6xJHJYEPPZEQHeDZ
ewHb3R0cd/BC8BF8Wls1YyTTyRPu1bQ1BAYr8JsubyZ+08mvLK27dsCeSjAD
SfE5SyplixB2uYC+8TrfJv21YtKSraARunUY7K1F+rBpEfWpHLgRX8YJQoYw
n7rgyw8CPxC5eBxZaj3dntw+p2aRtNPGjbBnGr7aV1XqEGwYyTVjIXoTRWBy
m0Kj88Byo4LMUfr+cycNwLDxvAAJuaeT/YKOopQ8Uwzq+imbQCT+tqXpcDUS
RUMqCAy8rcf6hYBtQOH3iF8JB+VzzIs9K+VHijlRoBzfeit78G7CiZ4HHcXZ
kaaRd+7Eig71exXxC/gTGdEx/EXVGl6ORYWdhUdnX12s6ZfnpXL6l3HK22zE
utDdG77eyAr47R8nLmPwjyF1YPKuJ7J2xk5Ba7IaO43r3TRUB+uxbbVMVsVs
ZuQtBSXhrtq8ugOTCgkw7FqVx3A04MScrA1U3SRkd6OT+ikPxlJEAUdNdL4P
xBYY+qasMB849XCXj0vmKF/saprxL3FsGbYyryOq/HjB3nqZBlKbcpMCpqqY
HLnLO2DOBU/lMMemKyR1SdNCLIbWPQSS8D9GUZxbrepHXeEk/fK8O2wkVCV/
DXrkitVcMFE2eKtNz/ttPmGPoO1IDrHp3USKMPYuhVMUqlbtSoBffDz7BkqN
WaTBEm8HEGEaPpzd3JroEQoieUqnZ3tlygtKjCEDImKa0LWc2+3FB2N94HeO
hAWfZnfBYVJOtFhug+vwJsXGPWu8wesqS9oOncO9JJAL3785mEeYUQ5GGQ/C
La2C3y/kzHL0te5PomVtVp/EbaaxLYKvGXbsMTiDzT7wdyY6TZU1tvdaWOeN
jcKEbTdKfZVF4vdiRPXLBrxIgNhSLO7jPi8+p3G3YFAivZJZ2PNaEU0A4UeU
vK7zQoZc/ogD16JbdbOUspC7Ps72t9AkzIb7/wxWN7/kNLMAEoeuGUwjwE1w
xq5Gc+io9+mjYJMPx3qT6OJlY6Zk3Gl5s+YxyjROPVzUH4vq4oenmuL3F1FY
5zbZHqVzZnevbPu9JVwmvMACpuFWyhu314zKZQrYvaA5r2AWQV/DHWDgJCf7
GSKvX/7u4pK3UGRTJw08VpzhuVDb/V9rFLywcZ6mAAmx9J162UpIyCTluWYF
EcIsiaFUya+IAIsLLrkTgLIHj1JmqY/yb8BGiD9X62RZsktyhUAfPetximFb
TinmJVeapbrLKFLeqS3k/flqlH4mmDNkZhCf8jbPcufenn6AnxIWJwi87xU6
cHIEXSVR+KHeYbn/L4nBqjlbTsvFnOs0emz7XRIOVGYsd6+PA6LbgKVvXWQx
2KihB9NMQaMH7zZ5oZRSzwr7Ril+O5EmrBD0PsBY2NU7jj8aD9+eaRgm5R+q
zy5d4Ga6Ye61/X2YgS6kMgmrgJCVfDcGFGGV3bkxyWO9gVSE18Y8OaRFkpZu
7mHRyQ/41aYeJ0OCXgHynfZaiIKU06Xv1TkS2uZv5xX7jBxRlTi2REyz+9QL
qqNOfYCQWar0EjvvhltN8G0/aFE973bfo688/YX+grjlkOHNCU34ygO18Ro7
bkP8Sg5F112IfXLcfry3Tq3iKYi+CpB0xlIAtUE8xF999bG8et04y7U3H5VJ
lbI0MhAUf40Xkrr3v6Q5gw1IF0Fg0FN14oWnhVxUXlSRCHrhorlqJc3aJZWF
d+tE9rQvAizp3DNv0+WpZQB5tjO1hAkhaVQgcXPg8EHi8hCXZKr6HPtHhJJr
6gZdteONaO/HvcRGdw3ET4mQ+DpKaeDryI0h5C69zSLoZmCrHJJFzQwU7NAB
PjzOa1GfTSqbvmwyxWoprT6Hkk4ID0Enz/P34mR+qsELRKFWoKkLgotrrGoG
Vsa4L+bh/Eb6F9drFWTbkfPUa2jH8vTB7j1qwYu2rcI8Q2vXJebxSOG1VW3Q
U6fcO/jiKcMewl+8ESgYLTxnkLWx4Y/XCn7ebjZAgkWw4/7jIkoTBQNWn8W3
tnjOHLKLpFb449tqyYD+0SffWW+iBlvj26pnx94zGVM93voEZUNR7CH5p5KJ
Rl+jTLDQiSiexmAtb/b8Hrdv/mm5zatjEfwC0p6R2EpTHwheU4nKJMuhA/dC
sr+NclnLSvRHZIWzzV3M6lO/qT2n3eADUKKiCS+Zn5ZoPzkz8VpWkI0RDk6F
jmYUhTUB7K0bRG81RtM71OYU7KMMaT/mJtMKDiIcI3VdfMkeL2avgA/4BhnT
vKJUeyp2NNqrEyeUIM2ghkF8NfxhRJ/joliVlRu0syiH81th0oMaJTbzPjEh
kTYaSJwQeOyUzz1d7tfJ6Hrlw3vL5ImLwn2cETStaOiZCtqvoMb50Nb0Y5ww
KBpwdGPnh3tKBzs/SPpCPCw6BcnU4aEwwf2wWN8++Uztmxj/6Ha46vNaE0Z/
7e+0O4kHon4YJFuQ+PjxTJI1WkDPZ/0Lm0tatPBLSZ8lXRnyJCU4eTwranqG
QieEnRYQD6XanZAU7oQz0nwPXX6qNhWZTUugrlJOKqruPb68x50hQZvJnbuM
dhy6ToScnzWsM5QbOXlZjkdMoc2ARX/TwObv5aJV1ax7WP+v975evTx5/O0W
UveNVQhn9VI93c2ViRVDqJr4OCa/trdEIvDDGtzmjYU8WFqqbZ4YzpMBfVjV
XfYMxTWiZi6k0Aj5es8IW7j57c1g3SR2Jnk6LXlk44zhE7X7I/JDsfMZYCgl
Y/zIaYbbNEUUq1m8LecxQnZ1FTUhwAvj9wn+zyhlEnHgOcv5YbBDH6QquWN1
4C+YKSGlc78ko66wE884P0egZHgEt/82K0Pkf13DM/BSL4p3mO/VQXs3XfXZ
+tGtBOj0KkqwFhX9Bj+caaqwdBHriHutyvbomgfWOCIJSNzhzSojETSgUooO
LEygtI4yswE5w3jQ/ozX8MXnHfkRwUneEzl6jhp7batvuRFCSCoudquj9GR8
rx32JQPsB055KJN7gMIGhDn/Afi0fWwQmH+PH1bEOX0Fru3V5YkAGkoBBo6B
SXYyeSw77kWMZsIMjpvVp4bWvE39klYWE4bGwgddhjqcg5qpvbceK1FLz+qW
oc3FQ5u+tr3WO3Um6hLmshcmnc4VJ7rY0deJ8a9AODBpS8sufABgdGuQGoa8
guBdrYXgLadmmK4SnLok+bAm7VT7FybFDgD5egnlSC3iCiQofWI5O/3pJZV4
dE6As9vuqJdRgFgAe9i1l1lz0SGd9d07qCjHZpjd0CeBpbsL22HzMsKrbI9d
S+u3uVJ8ePwKDnLE/7syTLGG734sZ/zjQ8xVTH9XuzBUzLm3II22xIvzdRgh
di3JQN/Cn0U475W4eX5uTdb6s9jUr7aLSBi7KTqgHwE2yiji3SXPSOvwfzk1
vjZsSKlKm2dD+ImyeEdm+2Sv8fcafyERICjYHy4TxxZ0s+H4YKerkMA9D/eI
07Xrs7L1A7RbOpEMQ4hOyaGqiUr6fwuIjBGQK6P+qan4TCERbwU/R+Hl9msR
Z3JXf2WO4vFIvNWtiNjcUv5anIRet3+aRazpdqHdsJAD8sfLPizr96oKCcSZ
ADEEIwIPGlWgjVPMPb/mEYyTe27UmdigR9SqhXXsNa/Ec4cEs5DAKkN2xoMv
9gj14iSmsWX0OzAOwmlmLyI0JCa8A2Fe5P/QeBh0YVMVZDEm8TLal8bvtMvc
lAp/Pqt/c0k6JJNfKq1c8XEWsp+dLe89aNf8ZTVnZxVV83cPCaO6no8ejpr1
lXNr0FT6CQL4BwjA6/qHSO49tqHroEajFj36EnKRG+kJ7w48/Mq3HC+H73Dv
l1jGJAHDWx6ogVU0uOyHXLxbxF8vAIQncyaJX76Xq1aGW4+yYyjS4vC5A80Y
4yEF4cEbLyXfx0v3d0JMFnjyGaeBkBQ3+vGPREW4PHi8YSY4BFQs/J9SfZw4
dgvngRJUp1sM3ooK204wwv9WlWpzrY04S8aPfvxaiVSZwfGo2JTIVqSkAk+f
eHjRgCmDkwuV0PSLb6fYQXjX8p6kUn38vFFrt72FOIm8BBgBOEowtOXUe2hV
IBdVk6jBzAjZmaD9XeJ9H7o1cXi/rMyUWVaI9jBMEevEw12chN2JnJ3/em6l
s3josGknNqVDTgWcGRIN6fnXSzEpjw7V7o8FQ0pqvidh+V7RIna5794fpCeT
Tj7HEpTK7yJQCmlrBCYoeeDRUiSIEzfZuOEKxg4d5apNBNgYGAki34GBhS2o
rmCVz0oAv73TI33vpRMD3nCrjJC96+zWTQlPSfm06Lid/eIKw0EoCAhVHXhH
1SSJ7L3K+VtkZjx577pBC1lgNqcRljB+NV2j2EluVcvw63eTWIawc7+GpiJH
7URJ1AAg3faPuZtkpcq7u74THhtAO2fvXVu1oonx7C76l5Qb3hSoTym6hdA2
40quwvw2Wl9B2U6eRpuvqc9V+PY9+llzBYi5tP73gVEE+QkhfFvzwIP9eHtJ
u2+TjSWzLqI7U4dKTvdawzg6Qju8cEiezTX3Y22dgJ2iXLR0b/vGmUiGtlLH
HAZAbGBcOe/zhWptSlPDRe0QF8rs3WV7NwuwX9QzcHuXvSmUIG9LBeG5gZTa
GZ5l1zE0E48CHQd1uCs38GjepjhDjF1qE+ye1a9xb+HacbvVt3RIolBvM8g1
RL0W7zhSCtLhK1TZf7OXKMmKYEInflNLcMTFs+D6/BXm7Q05bZ3QWtaUQwqC
0ZE3NcvJmoGb3Z+VleyLwePWIt7+rFnB0VpAxJAuvoNjpldNj72UKb2lNcvP
ba9oyPvwdQOsmua+zB1GJX+18uLJdRPkzjLM6bLsPnV0/v/JF+nhGyzCO2SQ
chPHwB3l5xVVFLs3rml3rVyNSzLIEtN14VEUXEfqyPyDvH4b0OnMaEzOADeQ
RvTH6JxHtA9Fkol9DEZWJVDWX3IWlYdzEV4owNgVuJli7a18cAwoj3PqaW1G
6k05BcqAhu1w4hQSqTB2y6fxxIKmWTkzD34AimkbYRxSSwiZK8sSP+UgK+zB
ZLm+txpBeEFsrva/oApQVvP1chOOScXKujZNmob0vSdJmgsN12Xrnph4j+Jk
SZWQbiZqoqz65RoFAb2JCIfTNtqQLzv7vvLoI6Psz7660MQQadn1D6nNH+TL
3QG5LTemjPXavQnEmH5p6uFu7TVd4dLO3RPzqLIHYBEkyjV4Pwyb9OBpY5G4
DlslLXNEleGFh207YWeK8Oe9669MZ87wKXVDtfMVN0/umyF3cgjmYhIgJWl7
uePpgCCmIb3QgEzo6cjIIG0BmwjOqbi/EOjAUcakuci4raOoJ/g5MBzjWUO8
xSI/18HInlVb1J7Ok3I4CxYLhR0NOp7a5PE9OXm401DezdXkAuIuLjSRQqQK
8ONfirg/Qge8/YmO9uxZuWDLUAXCs46ud6smB5ddkq7iA09Vx1wO94Gin4TI
6MHsJiPXZrl7evCaXV9NxJ6nJLwarSRr2yVaZjaA9n76fnN8jDGbruCzfrky
Nvctx5rBFSQtKcRrva6sQzJ0E8BZu0ArkLSSrgzonTkd+i810uUybXo9T6jW
RFyCdd3bMjcOUj4+xCCur6Z8bXdyL2g+tD/wuu3APRab3dh6Q1O6eXL86/aX
YGmFcSabe+qszTWL2pq7v87DAYAA5lqpbu0F1upf/HCGPHd4k8s7ex2pj/ms
sIi6SC3goN0p3wX1XKenSg/Dl1xE9s3yRkapfk4Bb1gRvT1QRxMU5xj7+pDC
pZfLKQW3JaY4khfkcIaAnC5aka1NHfPjMS1Wb/LOtfSC/aldbr1Fv/D7D/Y2
/t5RTI8QH/nv94hb0N48rOKr/jDOaTQLlZSD2bQ0vbB2QfqzLA3apKT3UZdz
KAPCDhANJxQLyHRxv1HuGPcRSwsbpysY0Xf0pPEkxGLWT5kLrcgrfuhx2Gvi
gWucafxuekwnGIzcFUVchvfhWDu6hXrMg649/CGepMOGyShhho74+g7DYYwN
l692tdRrTtpZaporRdI8dpVromc6Orc6eqDHwoWKkPLcWbH7lCBhFV8xvxra
Qi3qHgSZi/Sj5JNsbqdCMjYBUHlP2SLisugWGGUMV9NMzdlUny8ZnEdFnQUg
7LoVKSqp0Cv7Qc12rT7Dpc76tgR/ou8t10RdNwJvnKQP+IyOkMGOE8ReUM8H
WdklXrKycZmOFhznTBIexlgJFwBumyvAnbBjAQfIByJfL00XKAX4zaeqR/bu
gGXwYmIJMvVlM16b77wWprzFwwItsmtM152Fi8Z/W0iU6NruTekez/tLu7G7
Bnc/O0toeQec8aYDLKMHYW3qA5sTXa+a2szepvg+l/gwr9qoeXToEA8JuJXu
FIbrT+K1/bbbcgzMlZcxbgCBDRmKuVjkIMA3ya9AB8pxHh5aft2wzGGHiFVj
9ZIlbRr9e70J4Bm9fbobqBUa+/0uvfX74H3fITOXMyHF6Xi0yfq+avm5uYu5
pXoiw19Nk8nMw0f3BnsCY4MJMYZTh3a9RhC+sVN1aEGJe62DtP3tV9gNODV8
EOUWlb70zz7DhRp0YZu6OGRncP0dX1XeGmU7XpiWimddpx4m7B6ktuckHvD0
c9sZwwYR4ejiYENUBo7YSzDiraZ7kOzHyoJI9I4MbNeUuY2WqcBK5UKsJE6N
edQ5gXmqDuXXYMYNQ/FZg/E6MbgVch7zlry6n9+ALFGIDecNjfwlUp7d0QY6
xxUH3oUl6tao26M/VZKhgvi88MlJGGjncZ4usPK2oxnuppDBLYUwegkr7nhB
9fZMLvSU461WDqZSdhpiMooKOt20hdLTXLQRYHdWOG/CS3m60PW10DuQB3in
oRirlmxgnnbcq77XzGDYJMbugy0OQ7RjePOf/0d0OuLYd6MwxOge9H3LqPtI
WKXV1oWPlZGGk9cqNcXvjpdjKT4x7yJHl9M7yRnnaBYQOkuFD/QxH5v9DS+i
W13SMKePgyIFYjeV5JhgADFibh5Z7aAfyeSMPmUFZtKTI6edilgwbGP1Wm9p
eY61LVXA3oiRhFVX7gYlIJMirTWuJpUmk/Z0SUtKYxvNGx7o6Bnaot5AYZdT
wL/4Mjeg5es6+H1ePKODd1qOkGLexlxCeNza6fYEJlNpDElfXxOBOcDWU6/i
ZYpIljGD5br2szNjcsQhxBQ74llpQWliyJmnZXgQUWTCCNrUM4EInpdnihl9
DIOEAwkiFx0KAczyKpbOURTJNqTVQHvhHwGRfnGK+odGQ2LwSaSzeZIQnEt2
9cdAMB5J2FX91AeaHFI2tkA+h6PVCpFscFpU/l9xco/s7DFWt+20hKS6uA4g
fe7Thh7HYmzf6KemUv9kG5YKPSWyVf+B6xnVFoDOvJbF52mCVM5s9FJahxqG
1GOG3qJtjrlkifEfcf+eVX/I9+3r9o15dKnOtvTLBxjqaw2UBKseGq2ENsq7
HVizd/MGABaDG1/wsowSrVT/f4pRBwYInhV5XKyv1uo3NQ+qqRaoNnk+Hfsk
Oabcx7URLB4lseiijsaWPQxtNL8A7z69pjM8v5Ioi/PzkHN9/Sy/RxOJgo7N
UdNsBuGrzoSsbfxWJzlwxGSCkMAstD0ZJ77tT5rsOAhOXiV2sogwy8HAInxU
chOu+jB+UEFgYNFZbOYlK9oCTsv1FYYjPAIj7lSuYufUIwVbew0D/cT8y7XT
fj1YTK4VtVR35kvXhvgdCpO3gBL62W6CnGdX+HXMwXZO/Xg9ke8jyyxoSBCk
xZoV+rLHt1DzjwfTwpDcXY3YCYEPEu/BxIYW5bfFUOTf8WEU3edUDrnYFTOY
au6qyqR0O/2hELhQNSwPZkFUEFUEHoFM88IcK0wiuZ1A9sBgBptNQj6OC3+G
KYBseI2+ElJzwmbPr/RAlPbBWm4V5rMKS51o4qY3XYvXwBylTnU9FreSSEyU
fuyO08dTCYjCbyHovpfrEZ3UbLWoT15pHMCGZGEmcMLLq1p9pxoLlSGkDfI6
pA/lD2s8Bn8OtoTPjCPvLLuLZ14KFUvwTZCUtgSLMREqNRBc5SCBNbac4oBd
fYiALo82aBVc+N1znjWxU0VvxfOefQmcY3yR3JwLtGmlfP8TGkTsgno+KT4I
CXEFP9jEd0Jqv52XNT79mQeE2VOBnrMF0ho9/v0cuQ==

`pragma protect end_protected
