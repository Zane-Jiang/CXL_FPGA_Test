// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
46uO9C/Mc1/sKuF+Tq4QzseJwhYTlv6vUv8748gCH3hS3ERBFO+lCYZ5OLK/oon2
zVb2akjDmSqHMKQSZfOxvITB/UkQUFYqmpufr4zP7HHKSKlgXZlyK4qpp0jOawHs
O8c2ytZXj4yOYgw7H8ReinM3VmsGu9gmn4LMXNzAStFMFg6e5sChRw==
//pragma protect end_key_block
//pragma protect digest_block
qXIG26bcr99XD722qv59BY614Rs=
//pragma protect end_digest_block
//pragma protect data_block
5wKAhkd9Idf3JR1P66ROP5VwLh/UxMTULyjZjXrxVuH7DkBRMIzn5xettzt+flcN
nDPKFPoNBvj/8t5wzVI2GrWlIjSkp8dkoYl/VkZ7JytWTqfW3r0x9ZmmGMX2E1FI
ZzMTm6wUbkTwdz54UbH33PZsXExY4NVJIU3RW4+5taGDnn7QTAOMKRtHnE48UlUH
SzKQ0Ot5ahnMYF6WAfo2gfrYiIP0Cg+Gepo5i5H5dmBvreYxEoYc0ka3O7vfsRVA
rGE9O1n8ejeHeEXIZ3cxeoXli9IQmKawtAEHB64q3oE/MLxwulcCl5dY/B+zefkl
qYHkZc4QSraYTEE7g37ftywuuWO/ScOiMClb5+iQwEpMTT8otmq85ope6ERYuWTp
iMTgHrufzoYUddt5LhfcwQXI+wwR50kyEg8OrffrWhe/yUJThV/d5JdP5ehY/VoN
H5Q5TUyffKnFYOoY/UPJi/K+uom0FbUJ/XQo5Qia9XJFTLI6v9KXoKEMheMK8Aae
2Vg89yVjPnrQLH2DEnLuHY2g3qctjJQm4yIIUnt/C13oHZiIsQs2NbfsArVT2ojO
h4198BfFAJtViTky17iTYUkxvFi/xnTglg6lGK0vlizbABFSFEIkBefai3nkDYJm
VeHjyvtAdOrzpPwkVYy/t/mSpUbpylxytD0Y39MQSh/sHhpFjWmBPXsPIXC9h5hl
WtU9KNJFiu2CMe5SnRFzM7f86MMpAxfypIvvrEcDmCEgPVF5RCUonYQHht35kXAk
sAf42rbQ8WwtbGdpStajPY/8nwoyz2cGi/9NBQ6mxDtRdgv70zYVBI+LiWwr/mcj
s6ojO3H79KBCnRcRHiQ/wiUwnlpUa9bQ48EC/nB7yriI7skvbyzLXh+mB/SRviJH
uRnOEazD5/3p5TnS24sJHN7IUkrkXpTeANgkl+OfxbDiYYbVYPKN54YhzrXAAmvt
pnFa+moD20COTIIighHLsDQb8FRSDnNft+49WqkmbcjeVSr2KeMF7TzNaUb6h0UT
PO2+g6MY2Il3rBjRBp1PYAY7KbkmJ/Uwv0W0kAthyZcLmSR0NEiYAzOkL/HmMFxV
61uc9kJVrS0d6T7ZRDVNr/ANTfu1rNQE5vjY6IxDkIqkg+rjP5Cr03XcDa+bvZKK
0iRmU2SkQlVSChhz3i+O37wgxi1B/Mx/xJVH1QvHG0FSuHNdkYDUbeGKE+WxlzEG
D9y0zRBHgHIPiybciE4j7JwjvNBoUT6Iq+oU1hXH9q+XA/GJ/C3k2XbWkKXC+btd
aVr+wkJ9dp8A+BMUw7oTX7VAPkhpkrjBjgmT+gwL18QlKRqKu2Nlx9o39syqfUJ4
3pfDzEB7yrkfvK2WSR5+htgmeYoHo6Guw/Ss7sxKrvbHiuCMl+4Pghz9L7FsWhHG
C+cwbRTvNMAMTbD7XQGwFSsjq7V4soKpFUMslVBsJVpARhbgAkiVRC5Y3HzXldSp
HjKMbZW2gAilcr+xaC29ZbVlIwG9yIH4uc4XC/bgA7jdwg7c3kxKW3pRcmZoHxfR
YdvPtnQJW+9pNJon1AuWrGnv6GOsdoR7HazWqGtZ7PguLnDWisoUZ3F7TynYCaLf
Uy9VPbxjqt8NB0FGHzx7cTCYNfnBl/rYIyOYmEJN8o82BbVR8W+bdpjnXrGZte3C
BR3CKhgomEuWR7rIWjqf6biuY8w/8o5IbR7n9R5JPB5Cu76hSP0fDi1kbVC/2597
Asq2SIFBMo+IfwvPZTAmcMbuH6UD5TCol77mL3Yh7Yf+kEjtAoSZ9BJooR7GSFA8
UoRozVjZB4OYPvL20TXu6dfq3IrCI/C9c6s9Gy7NEjGo/C9EMOhYkdkBevpkWsxb
adTMI8f8TMjL3fIiTZb7n8MjJe/CZxIUje+ntkCv87H6n7b8SCeKYcYpmVC+TnvK
dF42F26ACCN03nim+zjUhJcj5MhQ1md1exgHd18DJema1cbYca6cSuJYzv8cWYWk
Gjgvee53L/Te3X+JQTMSWs+yRWqBfdKcYwZ5GC4GVVcFaehLz02xU9OoKPYxHcGT
NGKkIUQS/B/HkRxoAg1TG+RqMn2nVaDpCpHzjqYBe3t6o5+rRXWGP6jZWGsE275t
P1TE/aGo0Efz7TrPqVzCx8kZo4ELBQBv6dzdKiTzIPli7flXBOaL7gdh1YG7skg2
+BkXVSvdqSDxkpfrQ/A8dJWc56SopUoMXg0lC3SxliCOPYEmnieWEPCrQGO1OHzN
+NSUlWuMvD1c+YbmLegLJZoFK3CAiF4WrviyboOGXNB+FZ1VG9dogDZ9753tzhGu
FIHUDm99hq148m/Pk1FDf61VsAbzR927b02+MjnbP07WRe0esOSXNcKf41jTv/XJ
A6P7sW0YQJNNxoXeA8lPeoA8C7ii/ewG+HRkKBtbeRgZbDcRApraHoT7EBpahz5s
8hzy1YcjFxvYvd93NjsexroRAXQxm1iIO3V68EbjsPMruQz39XePq5vVFp11ZxvS
Gipf39TLsKHFBdYiC6z3Wtd30wvmaoBP26hkYezo2NKCMmv9gBitYKbxtnw6YJ47
l5ZSa4LQZIibQQR2cZBqymUj+9ggMm6Bi2hHUQMnAoUMZbdaQohCsfNrDehHDxAP
ahWPeXA8jYs1QYHn+2jhdHzEdZ4Q9YqyFEF/AQlljFnW9/lCU5rvcBq+hPfPAxeh
bzqAHy8YH+rBIeMiSoWPv6fPvcNRBSqGYL8FpKA82NuvY6jfhDtRMSUHyafiS9D7
kPf0ie0zEFAkAeJzN/ld08cz+5vh/OE9QMACkWbBtxULqVVq71vJLPDxITHs3HDx
MoJYA7pejnprKEeidfuy6KVUlBW2LIRjrEtDURAvBAh1szCLx4x7hBJcSFae/eeb
m+xqM4dBCDZ8G0fICWvbl5OWqmysJkQ/eXPlOEsyZHc/a/OzCh5WJAmTbOX06ygj
92pCcnJCQN37ArPoM4P/jPljK/b+ZZQbEpK71wKJqk5NnqFLQILU/7Verl0w4VIq
HxcBqI4XbJJoCt+z0wYDVpf34+TsDljdl8gsyOiJdf9RPp6s864Fqr4k7GWhYpV/
rrKE8GOjxYF4Zz16U9Hd1fIt9lC3xNJ5esTofgt2HYxoNVKqO4s5sQdDeL/jm3ZS
pKlsZ2841fMh7DMQrlq6KiX2m4dhej4ziYoF3Rvb0sqkDJElN9h8GTalZa4vimC4
2khbDSsl2Q9QoTjPlkDwsRs2NaFYKbCFkSzSxYSYZ6MknUAoerDUGw891/v8L0ha
Z0Ud7Fbt7c6OewYqyeqiPM5zzX0deuyno7cBHnLKmqG5JtC8gpAT0VaQ/zmBjNTJ
lNRBMjDpX/21f0jNJnZ030HkR1zFUPc69oD6O/7W/o30SHRjL2/TDnq7AGMjkMny
Il6jCzBLGuvas+A6v+HaYi3ODV7NTcyl7REign33l7lIUhJ9NpA7n0/JSJo2lxqg
2Pznz1NtiRtbTzM/cOuV5EjN/+zQsPIqOuY6PiJuoTSlxNNouQiCAgmWMLCcV27k
JMmd1w8j4vpVohGTgmC0/iYq8SZXvV8OHiEyNoh5BDqtr9YRqjj1lc8MoSk4pa9w
7NC9AtkEnrTK2UqfN2odbpc3hx1aolRV4CxOew0danILTx0fwYcNtldYQ8R+pN0j
bwZ6ckn75z5Px6oViWSytIQoj53Uc662c/RgJONKkM5AbbfDPmxoUi9Vv6B8+TbT
jCIjGFFBXWHKZ7h64loqCulY05dibOQyuYoenPX1CY+YP/3aQXwcOXcxHxUDYMPK
N/TBrATh9ozlkPI8TcjuEVdb0qkR5fpmb7OIY4lROzQXqSEKktDHz1mCcQJuje4W
DSWNZBc+EgRmFP1KrbTE64TaG6bVC07BUcioKhcWQo+xSlQsYjlTiESA9akn4Sf4
kYcdTjm1Jg0kEviXlPLPWKsTnGameG84bxLqhWpTKoJOp9IDZM/5vOayg72U5yEN
LzkS7u/CVfsTPHOAezz9f3Sp826KmQYPmT6Zh0S10bsDeqyMtHQ/J3JOSH6BLYFy
XVH2GjFLSUcYIcC9gJnxEOn7X0VvDa7WmAb8KgQ+HDChmCLiHufoOW+3XcX0emVO
DPIv4+gTPQ2K7gqLaR0h5lvYjGp5ji7f/YJr1nWjXswhDMnZG0hkZGTdZSmWOc6H
NvOFYd70H1A/bF2xSzeWdmcxIThH5NgvZ9Dx+8XcINV5ZuSboM6Te97vnVuiu66Q
BzGPjDKV++AjPI3TCEkpWyDWGCv4z+3AF8J5gVt9jBgzMsCR++tocg1YpMQUb7yM
y1j8j/C7Hk45rM2jUKT6/FgaPn75v1BIXW/iK1zgzWTy0C1UlKXvj8cm3Z9chWEu
8nsz38HlYOxiGd0HgM0mcqXvrzPJ3O3aPGtLUJ3huZUqIBCQdXwlhhKSPjqCnrRS
HB+Qq3S5IIBgOybHtYia+xM94Kb86mIBsmclM7NZKUnxuoSH0bJoGBA2EyJx+21J
nENc4agpK6kUVd5fHOLgVXMcnNdZhyetUktg05b30teqfglbu/XKluHBNMYeN4wc
EGEcXSUjW/j5Yw2iy9JmL6eknqyiI+V3JiTXSfuGSJPV5Phs8z8nSbv1Ixb/hgNV
pJYbCKMMfaIyIRpsWD7/MqDHz+sy4V5pq6DU5BUNrRRtZA5r3Y5/BArHKvbGrBZo
GTy1nkUy5BYlJxmzVk6DmiqoEe2ABxJdWCPet2LSilwYO3KNvuhstp4S0qeLCbeD
F+OQZJH5Lelhi7l6+8zfSpMpzZDeztj+KP0vN4m56dle2miIVx1ZRKR0u2hb7pu5
23EYFP83/3Hh/W+BZ0z4SU5BYRG7F0vFDm3lcHkEoMa5JBwCA/jB4oyf0xwx6GKf
RhU2n3yCeoYRhwWFjQtU3f7hD/zWpTAEAnNPpjYek8+M/bRLPybDkT5Yf2R19wv6
FTgIoGOF0r0MGK40Xva1xVP0mG3Uyyvn4VAZIrPF/MJHbrBryj37d7xelrvnqHrA
jIGJxYYCrdMuFUGHFJROkxaZCxNmWgC6eBjyEVmbfYUKoEE/SjvJ3wAgfRG8AVUB
IFq3spsKcpFkhMlw6Ns+xzOt+iUNlIzTheIKZZKVS05hfkwT+l+R3tSobUK48Iov
JEPD85cGYWgo7hv9jM6gYw6HeUzWtZIDRbiByC0QGOQQrfRiiRKWCspjlBnAGExQ
iabaAbn3odto9YewBZ9ZAOTjuEfPuwA0CCPqWJZX5ZPHQq4EvmChFlKCy3MSuAOV
UcQwP0VfWIsAjl2UEQI67h0hqZTBOx9X4J2fmRvvI+iVWhLfL3mvE5nwIVUPz6KU
eJHbvw6jE1yi3ltGwOSQF4vXcK2qBWjNVtbjE8i8XbiQjYvMAsHhbKIeVHxm9BWt
KjzolM5Iu3et+NT7X9cMbVJ86YdRjV+ro0oouVH3vWPEH762Zy1VZMDa+lqdWU8m
qvaWZ/31f9WEbxCy8X9VmrBofk4E7COxftC7JZaS6tBNs9YjpKoAPRubOuNu7cbl
a0xXyniFc990KcCpXEJZN2EcaRiM+/OCqCy/Te8Hrh+cUwsa9D5W+HrX5IQQNPeR
GTJbp/+byNv1TEvn8MYB7Maf9lbQHVVWRV1P8inGdqj7EbdsocsogHSqLQzjLCtB
vgiX/T3kkImJZAykt6GAA/30/Ll83fzvbw8P+USt+YidSsoVYDLI7XUl/FDPEzH/
NgVjFMRy2kgQ/U6gl65fMeBN0Mp3K2Xc65xGJptKtGiX/M158vnSHPf+lKywQVAz
OxmS3xWuI71UiAZ46Ik4MrXO0SmG4p2HV+1rgLQNVTJ124wMxqMTXeJ8XhhuJaYx
CUP1rsQaIyMrbsvhPa81L7xG6vX1HphcB/fYIfG1B3VcjeX8Jk+9QvCqXgJknMWM
FtTzu9N0ywmRMCc0OgRJJeiEVMZLWsHRuqxXpTTH18dKUMga4rxr+8cjSiSXyUwr
hYjV9hgwI+0nTFi1YuG+6MS+egA7yQMNmC5Ungwf1QdqUGXBhhblWPxiaZgvv3YQ
+HN8sWyiQvmXpcHvesOcZE6VzikJ2YqZ6TX07gh5vOfO08ayp1xukqHP4E3y6ISk
MNy8VckUpAwKcfcDXmQz4OkO6dCKh+1cF8DysHUrwE+gukzLt4POPA6Kw1ieY52f
gp0vhzvXzceQEpre5mkUcF3QNUICwPAFUjKHa+k5QDZWaYz2CqwoO+mlTAmEgufz
ImtxUuedyPbc53XB3lqe2OwGfpSINsNJEpSNUQqxDwQlqeNc5r6skDliRLJi3IwP
4iyS5kE5gLLSuYedlNnNrWnUZeZsiCOfOp1ct8rX03TrnnvoHkkIn8KK/+K8k5kW
R4vRT0Q1z7bwOmC0X4jSHUCdtZxmmVYp0dO+TOC67RoqFwBrOY/m/2hJdd6lFPEx
QwSAfqX7aBC9bOkyz68NTL5Z1Gpcmf3tLUJn9yu7U1oKmB1pf5EQ+bAMt5aSac+1
9wm09EeXAhlgnD6h5IY/bvZws+qH/3tKoZdcV3bn/GmZKlkMHxc7zEJrgsSDeCfD
M4br0gCn3NhvkFH71PBj7rOOSqPeepKIM+xC/IHN9xqrbQqZUkQ3RaI++1QyT6eA
XXskWvT0XbzQBQhW9wptLwEC8DLpQkR3sd5KWY+XHipF426TsQp1z8dGIBTMrLbb
149eIkhLa6IXHP5CmP3UzUuZLTFZqjv+TjfWDGVPxs0cWwSFvWsq9Rn0W8AzwazG
6gDKrvS1tQ1hp5Rx0PLWRzbTNdivhoKjFR07ZQTF8UnDUbvTUwWXpVQZrl3BVJN2
qAzIGd1DOEUZOOGu3zQrwUh+Ed0vGJYddGiHmNYvG0ti7i8ZGPDgPJY2XqgL+h/e
dFfewwapHuF6Ah1l1g9l46u3O49aC4XytO5cqd2fZEUiWXqbQi8RG5CHW7B9uivb
j6bR/g0dH6MmsXJCvrM58W3XHm84LdzXXY5w6KJkUvLEpwCPDcjK6vgU2L3bjhJH
/tAzl0rAhblqgw/mEMbfhdX1XAlSslej6DK3hdFeCLdzHCrB/bgRFuCCsn/Ug+oX
Tk2leTt6PMhDOrBA8YNnnmd+zFVT+XOYxKq9zfdJySGeBQv8KD8QpWxON1nXu24j
AE2foWAQ/TRbpuGC1uTsbZacH0lNWJmnJmDVC8U3DLoKuGhoXDjMjPh2j/ncOvnl
39IaKH+dBj9z7rjmuXs5EiZYSUxmhSN9uLfmanWaM44NfueMmJcTx5ExuST8out2
uMDOnWXsFiAsfT98hGyHlSxVUh2cPSfV+A5OZacwKuzkrEwyGuJ3hyMizu8/qXx7
L/ZoFjHtx4LHGLsG6z4Bmms0fkV4e1efDKd5SnP+nw559qncm8+rDk4coXgYfxrx
KLMkiHDK2JiDZwX8Tx2bJoDtryUVZkUnsglSerJMK4XhYkhdHYJ1rShDWR1bI9GB
jG/sPIMd3+Pzs0hWTUY5gkmYn0KjuWJ7LYKL4p5sFQ6L4+B/59Z9zujq1ZGLdhfT
mKOIxUzjLKcIiuC6GMDieAaw7dvBf4gIZDwlIRiR5e2eRi+4vq7NHdnaV2cvA7xK
EujYMR7L1U0gz7pfzCREx+sjqEWcostk0BWeE0XFxdQ=
//pragma protect end_data_block
//pragma protect digest_block
3ZJiTKxiHGVsNj1iW4pDpDyCaOk=
//pragma protect end_digest_block
//pragma protect end_protected
