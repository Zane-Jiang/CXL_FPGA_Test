// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wLWVOO+dR3OB39jQhGZkwH7DLWqLr0T4yxL8BlU3b3MvbLTke2RqXVUa9pyp
TrC/1JYwOnkYrKtEh5Hd+JCFQmwmlyzUlmSy6eXIWDMvmhBnPLgnah5ENMd4
sZfgo7rW7jpCxfHBPNlFDKqn4kdD/b4ln4K7CmLlnlL/Jpg0dOEIhN+IP2hZ
XmFNFPV/rBwNlBSNYRxQldKYgodA2ggXKI+3emOl2DS3V1bUHaCjdc+UqWxY
YW4zeH9qY77xjJ5I33bj9sAjm/uplmZvtzTOU3UqGps1UUiJK52rPX9oAw2h
caf0dfWiqJO+EqMeOOcWTa9obSjO102/HrgPAFSwlA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KzEmX8wDDKhXwJFPL3EibF3eSpooEHlocAHN6DXHEcEJ5clCZwmAK1gWh7+t
B/+7++LshYx5u4MpTVTaBUWYkN3oaMOuguMSp//Bpzg4HfGN9TRGWzjGBOMi
t5U3308ssfF5Q470IKKKjPUtmh+VlnuZzPgUsj4wNKMiZXw4UAHMRNr1OCIx
R0Wr0Qn3VJ53KhOlTb26OY6yM+UuUCEPot9JZzi0+/E+3HUiY0syH6AjDX5s
ZU/Suhqg9YUNWGZnWI5FNNLzFTjbpj434za+H590A19EQ1JFYTH6GgySADSy
fZq5lMFntp1WT6bcvLwGF64b/4Fnl9FuyEZwqjLWyQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mSVQT63w8d4y/TvQdAkFLNFvSvQ4sGst0v3OhtY7c2JaR17JFYHiOGk/5N6x
aPhOFdUg4uof9a3SMvkdBeJZcp53MqId4AOYjZx2BJwyR4Azj0p+KXr77Mxs
o2mXY8WpzLl/mI/cnjpsSki+IRzNQm5jz1pIaoWDsJhdTBoEBLQzB8MQih1G
WL3bJPGnj1R0zyT8is8NvN5ftdkeabX1kr0i+VEVbf5RewrPDwix6u4ttUKW
syUxNaUTpRde8TGeqyMOmRAeymPFSf+hiCeDaUVqkv7MF0lPIEt9cRIxCb2t
f3N8yKvjAFhN7hzzxc9pjau14t7yNNx5bktABHlm9A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FdeC67H1kczdGSCON8rV98C2IdgzS8vNPnNByn6uAeEfExt7nCR80qR0uMWj
e27+i6SfLf2ufMVwp9tdoKFwwwOyx3Dk6HRyfac3g07RUH+o4h79OqFCl6nC
AUYTc+EY0NQ1TafILF/D6WB9FkJ8koD3qTj+PPS9B3LXwGtkeBE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VIFMKsfL7AIFezun74PLnFgopjH0jaRASB7YH6E2An4f4zlUtmUSH4PpbQE6
D+auwnj2TQhviiFjTj/IZxwxHlFyJ02ZvLUlHlS1Uh+kcFRPu3OhICbRA2fr
bEh9Ts3uN22H9cIxAuMi/MZ+ZIdOt7afSeWf/TVQGsbKY74qvEXrH6VGTMIU
K8M+5SY9gNA7fe6wSN40wwIlEx618i4g6f19zMqCRBF9iQsrVT8QLqxroiUX
Ty7QWtgYPJF0diSlSLPpp7lwAeXYMj4CqYD5ol63RieWzqWEwV0Y9B7Jb3a/
UgETeMTsq6olKP1Jwz8CjBOIQ4UHZTn56hrE9O5lPRmvaO5fNDMbsHcteLAL
aCJL6MxypV5G05wRb/Eg8yLNE6y9q9xCGieJmlpQnKXd5ReRngaVPENcSINc
GrqVkRo5mWhc9HLXVx3nm4srsf7o+XiYsxPvvqTbUkuJw8N7f8N+2uWWBJ7+
2A6Zv/4Alj7x3jKwczWCMPXZSUM2LGlM


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iXPYFyIy4yQf9cc/IUX0Oo89DFvW6iFazJSzOTc/oR01ctC41koQRiw6GC9M
BDBX5UhshfMccLMN+VSjLJuRN5Vaa2a3EWcpaQdsD5/99o8eLWpYZGreJdF7
AKloAKuS3+4xfdhkcVFhg6+xq2pl8jo4FSU5N3VEM7Jyc1vFRLE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
syzz1+j2d3opiw9HBYsdj5s45uh/St6SA9Kn81ZENyfPZjOhXJfUzJKxhWkr
gsiKlZoSeTLMllmSBFuQGagex6Kua3czcq86Sqj8zSfAY5nFCbseaoTLO1qS
ijKb9LfUBZ9OVqw9Hdc2dNmbO6y2g+cGWxrx+nNeBVN9JHogs/o=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 151984)
`pragma protect data_block
ogILdabfTa5Z7prtl6r7hd6jxmtwqkYGM09FC3LUMVncGx5ualxE7U/U/NAT
JY2HhFn4S300QYc75KbNqN0dKNRQ8kBT2+LcHFOFmwtrRhPKKSiiV4UxpTtD
P8w/GH4af3POsNPQ6nmcxcKLQyxMubgcNLd+xSLao4uVjZiGpa7mhmAp5tBZ
tKI8GswTpGhU5sKBgdBbJovl3f1RZJjepsZLLdq2LbiOAQ0icEnMDISrrHgC
G3wnytHCI07MDfEKDhK5r0mg0H/W8l2aHOBaiX/iWfse8gakVug6aiS0csje
V7PMOC0/FFSRs41xqaFypssSfSjEM/A4vhbVO3LKeoZIMm85v+v+Arb88t+Y
ZckNtQbng6GRtF5dPIpy6W0J5WgBUwSVUjEol+a5hg2wJg0GUi2/8eEsMmEp
BHiCMt8OrJBaEhDvaJicsd3yq/R7OCKWdMnzH07N3SZBut9Z+u3AdSZN2h3x
fhzJH6qqx/2pn2tXfsSkOQ25uIIKOTeqMVBeT9klPdbGpjWeAB5X8MOTTS/w
aU109uEsy1072WLE6qPSkvJbp4gjI2UJfnF2qy4B4CYcfLRAhxHsgVzzlzD1
EF7CZWXWyZ9eoARHj8fhqn6x+ME/WWRI0OvkpWwwiKYbpVxKHrA27cLDQz4U
X8Ma1ybNA3u/JZZVc3JDd+bQwL43AsdX6C/y68ZjCGVYyzIT+5kLLh74SMLa
nBf7C8ZPCypchjM5rZW1+0CUjfkk45HL7UaJDTrVfcR4WZC8GtdOFAMkth4P
He3FjgMMd+IB4Xkl1INb79q68fwDcrCulBkxvWLfd7xiR3tAQrRGCEuGAK8t
aXy1YXnzDaR3qXZ+68yLWv/mlSei9tNp0ll7RWC7/rBTe+l4SxBUWxEeVxWE
uW64vA+hAl8j5Gow0xR4Z6mkqpthgaicl25v3ITtD6ZkCjT+FsZHf+E/T7wE
zvTzTbFow9VzLU/FgUVRaEVSTikIrn3yrfUO3ceLgveocrshslzxn31KmVko
XEVMz02mcp3MyQ8Q9GrfBETuSIOB3JivADTvU3ouDMTCHPo4lacHOGhDWo/7
pHn/2j/PMrpbxB5+vU4l2F/9vIAM90rdCUgv73mhprCcLg2gCt/z81K0rmRT
GscZCEaVjbjnTBgas1YIGL5/Nv0dKevZehS1NMbeHIn9HRLMu0hIpWyMFmCU
lUrjKQiDghmg0txluRZbpz2k2hYZukGOtvvedfv7skTCkeCf26G0Txceyh1f
BbWMlEsLSxga8U4nE5BxjOcUelSatWCNYUlbO6gbxVKrA3imBN39w1xTtJ+k
Hh+Sc+CSGmDzgazyJwvL+eFw6rY5kzxrlXcvp7/l8+hI+2pKusrPaxYaMKjD
9CcOdbnGyvkzlRuMxJk4w8PKD7I+w+EJbC4xZU3y1G0JPz7EtVWhSlVSfF3R
LLtdlo8uqABK3Og15EidWlNDq+kjafN7SPh4u3qXngjlO8p2SKGOue7KfwdW
38KRX6voZviKtPpZri+hOY927PuNrIkElVl4E6RU8qW1slJR/VNxdE0wj6oK
FotoLMJ6dh2+srxKErLFUM+15Ve9aphO4/w7cR6A9vG4Jd0VAf/2q4+E7Nn+
sf0TLjvXd8lZkrTsu3iipCfc5ezr/V4w2Nb7XO87bc/P2ZVDAqoHxaI7YMWd
EoICXxFYxMh7kh0l0hJOTBab0l62ss84muYu5+SR6MVWy2R8aizuyIrPEFgm
ubVFWNXqmXN5tDtaAW/U855iDHCj6AeXok5SPQEjRFqWkFNSH027JT6LcKVi
yyTfGXR5y/eHTuW6ciHREAsuIY4fj43lw4U+aNEa1PFwNCNAVTH5OKEcgQTQ
oM2s1iNA+FD6QcFL4DAXGyV2pR68Hf8xpxa/ahoZQV4UltnsDcbXX5Cq8ezD
prJLLkg0QE6Qlsd36WuaLtIes1cst61ZUEFJF4skGqV/t/uPZKaNLbiQSp4F
0ea9hZjQoRthSgehGxURgqxjtPuC81iQDJcHFq/sDeSR/ifu6u4YK1kxBjXE
ibjEnd9WVsaBk+SBfK3hRsMYN+4QB67XNgB2gb8eibM3pomwRtW4d0JtFk4T
iwzvt+J7NNZsOVPhDxPCnD29+or+KrpCr+ZRQmoyeGvPGkZhdhOvBFbSDxcf
CG5eJnmul/IVBaXfoHCUc/wLIOIxG5jWx1l2hPo9H2WKq5j/z4g+951G6SvW
haJMx0hvU0jiQNed/wA9ecLXMIUp3GvSDSGQva2zz9h1dEyvvvQtXFLmehK5
uAUbMFJrPdOebDm5CXkaM/Id+CagsJVv39b52Ytoln12jpuWrZg96QibyCsP
iJyMbUveKSCIHTLl+YyH+jrrGeSYcRoFhRyNbibEpdHwxGLrpzU5EWOjQyQH
lTYYvnmUCzOJEPOBbOeJBaARac5tywtZoZ5CJm1PjfactvOOdQMUDYdsT3MN
e+T2XpVmaXaJAUSrpDRH6u3Re6D2oUaWbbQujFteQ4aLPnEGCQMJE+UlkCb1
sA3L5g5dsh7RjjU7hr0sGn/oR6KDb8sd0wk83jQlmtqQw6voHs3NWSBK9DNq
wxP0MGIu/71ZEeU6AmZ4qV9Son+CmoVsotQy3cTpZlDqo0BwGNjup9hdNJRS
ZSg7uDv5YpkV8RIRn93MAKmmwgM0rQFSK8oqj+SR0E24Bd2F6B9pzggU0OVS
ahkurahd5uYtTMQQ5cUt8aa6d7VxuOu+qIlIKXa5IZSiAhoL8jzdv00FE5Mk
21RRyaqAxKr+Njn/oVUdS1mzBCJ8AuNkR7Zk4Wqw96qQew/50D3O79j513xT
lIkRdAUw5vEnKYqTTOFrkqoeg9Ypr9JolmcIKGc2q2aIkfKGjuKEy89EUkzz
hRedmy80QrIhtgfkmDCEyEImI7DSiBrzxCncPMHXh53fDFtxVvpXW65+THnd
hzyEuvDyyg/TiaFP3v+9jpRahuXSLTEuGTmHj+JxliruFGULr+uxhb8teEhR
agalr61Lg13FI+edrYN6a4/vBiQqWX7NycZKvgLbSU9DHMlj/em1U8swtZ9R
t9SsLPqJoYRzofovBKm+qLLOKWzNpMu1E9NsqJA+LOqFbijkI8C2oZdd5chF
6AlzWVdREGIAa9+B3cNozgHzDZVjR2ENV9y4mXoizBiWAANiw7G2qvl5MX5N
IbWLpgH/jeg8zXNatH7cby7HvE5q7rfFgATOWGB9w5Dpr8n7E/69Td3LZ2jH
ukpEiKV4/VMYQslNwo0WTB6Kj2wSiSxyEasDaGsemV5rBuGcXBflICOU3rx9
tH4jKLx/aJiIIID5RktF/qtJNUjJ6pjfVb6bUR0JrQNPc49qwJmdXsfIL6bI
0zuZJMU4VYNtOQV5ZqlfNCJPHguR71k534UY1DOSf1a+AAlvReGHi8fO4CeB
suz+XBF5Cg1DuDfOgo88/XyNKTffn30/QEXqCrFifNJTOOm+ymxKcVQjM6kH
LI8BQFff/++37dSmJX3l4VytGV65yfj+W2pIKsoaMUJwADg4RFnZF24MY1KC
ipNQDNTEc7N1DcAUahwl0UZYHgS6XJtJ34dMdUUyzxQBTmH9n1htoC2uW5ND
Pspv3KjtYlOjIc/Nq//HHTDCuYykJntGJmrTRJHpvaIQ2e9fmcyXOiqhElrw
q+xDAOhLmAfEiePzF6kmt3olH2Gd/eIhb0EoSXxkmAPEJX0OtI+D4bbBhXOO
+ofEbuCe7NTcAuhN94HA8b1r2zGqbUQgg/bSqxPVN+eTFHf4XWi8MLfwU1iC
hMKSb7W3+M/P805ivyQcYvDx9lGxaYCDnAoIHf33/HomkFUWXp+KLwlkVuqI
HX+h2YrlypQbewuD+ZsgizzntLM5vDA8Fkg07a6qF1pxHtYxYcYhKerp3kRH
RQhxwtzwjQ5DpZ4zBvlZ/9BwqOgaMV7vHsFuvYxOZTAJpRD7aj5ekZRBdPOT
qcSY0KcUsk/Bv3VEWduV9MMHGfXLy6jBFqoe4xmqOJo8+Ca8xhyB2BW2KyJx
ZPJl1gZXvJ7x9g7I568nyZgq6J/OWXsyvJmwiP5ZL1BHyOA5vwsUo0sXS7al
uCwjrVR0MHsTN8VrFeMs7Sgw8E0cfpZlG7efCx25swDd7lCAu3CiFQLn0xyo
8gZl2L6NKfGSvXEE8WbedS3OTGwhUcSO9G1pgvl8u0ZS9bib2lcB5VV7L1Qt
IN32KcWxycnRFTjmIQy1Sci9xbcrSNDDlrpkFYD8nQFbr8cY8vOuhx6o66ck
uHmeErt7UgY0Wbz9pAoFK3+KcPVF8EO+HadJGSZ8zJAQ0F0XPaoN+5bdDxwg
i9Rrm+EkISRxv0iP9Jn10RKxfdyPo0JXDxiiGtB3NffrdsGtOy9zsN/pYYBv
CC4JglIW3Twk1auDJeLh+9EjiWWU/fMiK8+U+gREnbibRwmYktdN/CLlIbgD
LRYSqSurZMRQmChrx/WlP2InHeIBF9vMXanUNTO0bihUgkddPFDorTAO+rCE
Vged4Sl+cI8M4o2Sr2bl6Rr8mjR/Yq9xtDf67g8UopUw6+aMGy3+e42f2L57
fqWdnylAUho0nU50uxMeK2gxLjiKpgVTgjxJtn6jxCVS0Z22evYtewnkcjnt
iSO6Bh6WVDyCiJz5NCS+Fcch9gZkTgenS0VlASXg0FmKJknsg8g/ZaPZOd+X
Mj/HYfEuOkiQKoeUPfs9hOx41P+arz0fQ1T4eHzGz+aSPDfLKIxLsnKwX5aM
qWZzJ68g2OeZ3zXas8+j1Gf/srpiVf/gZEKm278TgtQh4cKsVAfiittWNf9u
u8M4AXPI/71DRlArr6SuSRuUriQkP7bMYvAqFIKP/Hi4H4vkQt1wQxEJK0Us
A7Eba5xbKgucqsGWxhcKY4fscAyQEplePqNoIZ4E2zHGSUMMz2Xu1l1vAD/V
vMJllKNqT5LNLTclArodnUVJS9X09JRIm1sF1FecW0Hxk8fDj+NplVWOeUMZ
fV6OqyfQ4lEB7vQTHdOxVQ99OHdJTOFw4TCZGiCiptfkyn644WZjKYJEhWbn
PRO/xWMyLLIsY0LWHhmBvTBwPxp8eEfyOA5TXoLXLuX35PgxExnmFVUclQxZ
dXqlqst6aeoX0t83mL1pGSkCFrOt+V86RwIrXMR3F7IfuUaoyHGSlqWTqeM/
C6axJCWr5vzxCt/BXUWnMMG9b6/cZ20LpyXKghOFHnCkySHedM8g3mDwOuV1
RTldOF+0hrfAo62tHHfBJQ5dzBsrUbbqiNRicXoVDNrPZZVujBWP1FpXPAFN
wLcs9vmZM6ZbXzrVApYoljcB99q3NWNELTt0rneUgY2Y3+66KdfdL7XU9ARz
T2XixuJiukcDsUVI7XqiZVn1ktpR8fv1gFWevN7yVDhkW8YuBt7TUX6hw+Ey
h7TxDYCpnWBW/qbLcNKhWGHUftMwJ2YJdWVSuhgNHmBpqFC+mF3/6FrhZiym
FAiy7R2x6VY8s6ldLL41IYt59RsSDAedi0sXwaRAsGJtGdCnqoQB3CbVgkJb
znIJ5K/902vJDauYq5/GWYzLVgLdYg/5CVrbItOHg5zNa4bGhLcND+VsZNhU
ko/4hUZZUcB/4IxG+uoL7ANdKqDBScyGtspvPeS+i1xmrxBf18ztbDbFv0Jl
uuP9Nxi466q5Uxzd7TZr9QCL1YoC75khNtBgyrwIfrlApAzsmr1X41DSwwdO
BSbCRMpF8T6bM6IcvQbgzokANZgEtWNCBAUU1/zxhtme37iLeW9b2jB9c52m
ifl6YBcH15HfOTegTmJNB0ylFhVKsujqCnkxM6ubGEUaCR3FUYyz5yPZWoho
gXTBDF9kUw/BnR3SxJYgPQg969ghaThNYrG8DlvnTvn4oXMsSfrzilKqETe1
rVbH5PnRsYmS8CmRrD4wo7oBSwX3RCH9SZB3w4S54ojG7BqoNDZG/9aq1oWf
CMhkS0ni5kbydSj+Oh5uAR4qP6PRA0djK1IwNtO2Lo+sGVquwji/rbJ5mQin
QQKLnYybAfMIkC0OS6veTjQ4a8oEvZByjgYGbcDHMFeqK83+tQFsFn7/XjLK
I/9stT/axWHsqn/9cvDtx9+eUS9pToHYeGabp2lYCEnCwej5WYe1VbS6/Awd
AQWlrNNXO2ahbOupt7x6ez8VVc/DcV0uokpmHNQdAwZGBZP9d/vFjrPO8T5m
xj+p9ButEY8CKaKe9TuKy+GXIMGGoqlgv73eDsXhH1LqYCl4LiDK354kfMkn
n3uHo2bDL7gdtXquXL//S7aZ9oqDUjIYjDij/jmDbl9xgimUNFjy5L5Zg6Fo
BK7V2VaWYSVb2OToJ/6txDMFIrGX/ljVTzavKMk/4wGTvwPukqAMv7w/pZIi
WgYcCfazNH3qLCLbi73ca5J58cNN4ZE9zgdxt57EdWS9jVA864Pta1pUHy8/
N+ybxef0cgRwutyH6ywH2NVik/eKjdcVzt9WDX8ZqzDS6WjwYT+ksXduhA2n
sSlYdjmW8DmQh9y5uS3K7+6yCvvD+uyKIcvMOmzESzX8kNvlqg4Z0XqjTHl2
wZf6dobfB0Pc+iXRBDHoIQCaGl133rJ8ljtipEPJkCRQaS/PgO7RjKAcBeQe
i4iLaG9jILrIRhIQW0VO1908srLU0VIHmLy4dpVu/+Eykra8+VdtBlBZeUg1
GavpUHejeRaHeUeJ5Wj0aKkK2L543m0OBSBOFE7zpPdk0WIN00s/0XIkW56c
1mXTPCRSjt0L5Sdk+5QDTGM9EUgliUtadd0NWW4YtPE/PFUxyzuI9oyk79DX
pJIp70g/AsPAoLOHzORaVpWCzCdpTO/KLeKKfZEOm97RF+nA3Kmk8Oej+SVt
3oLIT+uvNvc7DQqxY5kV2nURKhjr8CthjubmAAZOvFkq6tznJqAthJnDxDhV
ouxf3vXgrBIiDHokI8k/YfEndYZum/1YMqrfJB87AUms3emwAtbGxozb7Jku
zXTc2BBfdaaMSok0vVxPNDP5LLjJQkRin2GkFfqcjtwmvjgKzmO4T31H/8LL
yqlaepgwIK+phNYqtjXv6Ji7LUVGdsyPbtP4+svIUZXv3MVxhg9q2iptgWdQ
6EnBp73JXSJrqRSQGspSqUaNuWJfskJOExVbqiUxMgOAIiWIRdiPQFaWFzvi
ZYteFsz/NKYJ7kgaDosAP37QuuAkwH9g+t5Q+q9/p3r5S12oCU6lUW4TZsHz
lYVkXO/piR+1wINK/0BpGugFif7Fq2b9AY1NGjc7e9DmUBBm6o7zbEpPxWgL
bEONOwYHz2dNKj2ZtROoq4vYgJ6r+4vmJlUrgv/lO58TXhhyY7mETUif8RAk
cisGKLUCrN2SLJwor+sBfvkYKccVeoNL/ciUX6jPCez6JYehtxg/ENkZh6uY
ozkzHRY4d3+M4EA62aR5wbnO+5sntljXzBQAYKlNZMdnz/bJJTPNIaVrXVGB
X8pmb9BDA8TAAHMuJGsKZB3eXBbCg1gH+r4OVKZRIVCOqzvCEyyQDxJnbHNY
kF4/pssdvMZ8s78WNvI+eaaFVqDV1WX0GYuawQw9uKGqZejxUlDu03RADmom
jik7zDcBczNa986gLmrwmMy26VbICZt9HStqFYs5lfAZ9nD+BBPohVdu/Kj2
YMda9ATLUGbyWXtQ5iSHfEbt7WkOiiWVZLDS3jVfAKg3tCNR2p3xneUFOb1h
aadYU6m1TJ98cocA2FtrpOT/kpVfI6DZiq817CpY2Jb5lObQb9s8Wmaz9hgB
P6OWKqHUbpVGsCdenZRs8rSJXCfTDmDDBtg7VrXC+Z/E7VONtJc4CZH7+/aw
0/4O7hA/3Xn3X+6phkyJJ5bwKpk+JY9CEVboKawJlDwvmDHQjw47rJYHsEn1
9EC7ZfikmR6QeyPq6QjSFXOwbafoxdYrz4rg7qXFL87VbAjE86hUBzkwK6V3
0VnowrMVfrsjKY1QgghblSNgjmt0GxOW549I8Kyc/D2Zfh/vTx/Nsu881lYL
R4wypJox443cXYIDIvSxpiWRyDx5z6+UNy/AcEnAnv1hKMcH4l/DynxBQi3p
Wh61YZ5wSdsc3t58rCFTBtVcL8odCxNIIBZnmZW3lMQhNZpqXoY1vgda4ex3
obyV6R224T3FAv6E9i2mJudlq7hPvy3a0G3eot+RWv0T4B9F1LBtKrJqCcgD
4rdMnixc5lt/5akDmL5GdhmlCkWKhzvCM7NpY2cCUUBrFX23hMye7++z46eg
F8c3IUye7EhF5rzgbDOGZuCZsmKug07Ul/F+K2GbkD90V01McL/+ZX9XCTTS
8bURIs/FQ/XQMeUPgtOIT6PnuIWAYL3tZLtuSh9+0vgAQtpgq7UtwF7zG1Vo
fV8C7paTNtFyWtWV2N2h101T8nVD2NdPy1ycG42iVhbpBwKjK9ejUx6wWrj0
hpu3zFZYWNMTCNG2I1t5eJyxOzkyp7W6NaScCSZaTzvffLPM5D6N6gM1hpLv
lJFd/2l/H76ZVGBpWiodrWSY61rtr8LQkyJXoNPAC+VyoFnhcZgIHu2eI8Ne
3oROb8zpTZhe5PpRGoV78SktijU5fqLYT3JNbIoP/zlhB/+LuUOfMDhRosEX
ZJ93x+dlczS9Xq0sRjpwp52LgrlzlFteKX6pXqoZ4gIqFXdtjZNBHx7GLTiF
EW1G3c1lRuQuUEhuWTVq+sEtzD3nJAYA08n6lqmN3qRsrTYAkrc6jM/GZneh
Ofz1l4u2LgC6M11RscNXbOTofPP5tS5xRbWlcEEEiFA03+y55/4RQi3hfcwQ
nNlve26IY32UUVh1HS7RzYo/ZggBRFJWjn5ugEISQLePgz/lAxi/HrUQlnuk
OCfqgtjNPcPzAo99pSVdwscH6ap7jLT0uv6HGCOGKWleC/VmVfOOCB5UEnA0
XEBAUJmtLNDQl86v0TWLtUs9YOnIKx7tZZu1vHKXtna8CFqeFtaMdS3pTnue
TjiyWdzeaaQaqlXV9rDxnqtJJFbg0kFarunlzOttf/jgQaW1W7yTjhA0mkNE
/NhbYgybzNi/6o71cWOKJKCmPfRpwxubaIqGN3E2hCRFtre2w1fRqgKytweN
wnXWA4+Q2TnUuzUogTV25yWGd2ceWpmGG/I/pfAr+BPx9HOP2sa/zaQu8gji
j3OyP3kT2zqON80nDxjirsHmCi3kN5Jkt8JhjVGg5EWuwJfvkT8hPniwlg1O
DsEuauzY4mtcq4QLieHoiQXUifBRB3MP9gpfWCZP9ZAdY52G3NwQz3Wc+4Qi
DTqTsftl+PR4LozWNtO9V5VnHLrziALzaeshU2rtaf6KDRj6FUcFkn+ei4IQ
SWBh5qW2M8BdMd0tMaoOp7sIxql2Is+BkAzhFiYdEAGraRrK1qjAVgv7zXs8
MhRVRs2JE6dYBJjHSeainq3Er847O7ewFiGKAd/XVxh9LoK4qljIOiv/1ejn
bs/b9bSVzTFwfT54Z1m9VeD0LSJvo+eKHIZ4PEug10SjIKs5EE1p71lVPqhr
ls1jbytOu2xACZ9Gr0PJjzEeC8dyJb2fdemgyBgGxhzOnc11sq3kenmP938y
tWHUji/yr1VFXYneYhFd8SRRBL5FD/OY55TBpCCMrldSs4mAoU9jUxKXgvEB
wioGsFi0XP+nvRRx6slArA73+XB89SJVx3UuVXWkz2r4NJ1lek+T5f4cxGnT
wvzjyViIv0Q6nYxPxPKviPR1f4nPMqootqT5aeebruP0T0IEM1CdULF1MaTo
KUIjnhfih1XRfnqL2DGKhFt+eLuQ6ekZDXc8VXOk+5TVeSndfNUu4pImdEL9
Mhj6WSvQuDZeZHSJrh6mzZDt+anlU3gvRugDM4iUaLWhcuHuImn/Ma3RKnVn
m77KmL6Syc2YxDoXXV6Qn/9ZV7K5mBcPzIK5ztzqdHasJslJkI/dVnCBWESd
bNOr2qvK2SUGJVjZ0Xcll43hdseVgoDaW20LxguEdGw7UXTC4cTqrnZmV9nc
ZsMzUgQlR9maCbTXRyL2xG5qN9I6SK9cHX8PG7eGKxW67fap1VKVz6gexIAp
GdHzbpyoJsz3e+TD30BW8A/eaKlcYVUM64jDdYHbmvvlnf45kX3lvU50mjfe
5Sg6o8PiwsR926HKcADJq6thFpJzKZyQ8l75SnMM1ZftCybWZqTqw+pawORs
woxdMB67dw2a89MTm1a04RSQEDZZJnf6u523KQ7qXYoDvUX/y5EVxqMA4g0A
asiIIKNk+OM1m3KFhH69kDkgSEhUWX7XNpi9emssa6MRxtvx3AKJMztWQH6U
lTgk9YVLHm19khw02agU+4wRca/Jqm2LdCTZBX02tcK+DTJ6QLybWJLm8ap7
ojxXjIcGEBsA6swj1r3pVFztM7dIZ4uRinTV2+Bh2JnPm6yfhzgtk9ncdh0c
po/b/c4P0sji4o56duMR4DwXrOMGTNPQAKKZkUckNZalH5BLxIp8e2VCyltT
KuTlFDQi4HVVt1FTPywsm0jJ3fqZcnIQ7mj4+3vnJ8lWGr9wX8C96/ZEL+9L
NlVhKn1mCYK5ymZDcmVG48E/WGeLgbhPlGNHhW6JeYIlvsn9Pa3Ug265Zt3C
4TZWjKHsr17jZh3LuAVBZ8HLlQ6mvEBLybtF84+uSwBgc/Fb6yu9UpdTN7Hh
5vLsN5MKUOr6xQpBkOUUXaTeWLKNxXr+Q6TvKMMDYT26MTDt5ALgnpMNFUOL
oZLmc6x41GghISB6H8pcS2rbcTghDd6bmcqpn0oeAWr8y/DxCLGZuD9G4LhF
gnBVBVST2BOwLfZOIzgawwKjXydYY3IxKmRp1cV064De6H++SakcK+bfYof8
m4Dek63olwKqdllmcYfUk38l9GZ/yIH5E4SknNhkjCEoDuE2VY8hcZ533zfL
3pBJQccU+uYmLMiPyC9BM24lqJNNweIf9wjzJ5quNtCfmbwQKcBNg0r2LI6b
wH2KbtUXnODCKYlPpf773GrwwNZiGAwfxXNcusZRgv8YWtBXMFvE2J/AMreT
5FyAm8lDYVfdn971HrgroI2137SEoXulQRzlXBTwgSMy66SY7cSZ5D2jFMNe
Sd5XxBIiXz6GwAIJvdi00m45b5mzKaXhkjDNvdpRE+ZUNLo5Nvm2JHEeGyJB
RRQM2JpbM5Hdlm7RPfEN2PVbxzrO0EyvApEByNuTdHthDNQV4ZYR6BYs2PwA
j45F62QS4qZl16vqDfw2B4x1j37jj5FO075iNiwpTQghJnBXWZuubRjROwMb
+BCDK/BrgdLLn5SPVl6MQiH5CCLhJj/dJsTH6OtWrjc3Z4PYAvOxJUX0Pc2D
PnxaSM1DGZTwEjCN5yNlcq2ZkdyqGipKG1pE6QlJG4hS+IyJntm4IGoyfOAm
9MFkmnS5HdrwVj9gmiBOEQDgKmQEv5MRkUTqzre/mBXsfuM2e5guOE1SZxB1
JbFZptxt+95dDPmAa6a9scfBnV8cUUbH1W1fj0m3iw9evo0CrlDs3Hh8nAbJ
LKdsUejOGDNuMI7F8tquMkLBlRWrZINtmkXFnxCdSGjudn3InOCmu4gTplFu
f/FfsMF/55MenqkwC7aC03kFAcs+6+M9xudTQ8tMhyuoITrZbxD3nqSAUHBi
g3wbm3Hmh54YpaKMGVyZVNxXkFS3nusCj7wHO7T8TYCEZ0DSDrFhI0FsKjnG
2xHrloF03s3DuKEXPqAXE1QW0JXsiEc0zBRjDgeXfJoFKXShjeZCOA1zWNU2
7QJK09+QYTrW4cWu5DvbGOVUDK1bn3B5MCrOBC3D2xLaJZ92+7t/QUSfMhUB
lCldKz90UiYcXswbbK5f2D9kE+Xvj0UO8XrsOhzFWH6q/tLjsZ30zo9l2PQP
gHghJ3GFbPJ7G0aKBYloSE31R5QhyUES1SwIp4CtM+t9+jSeKxOnxe95gYUs
/BKMoobkB5PGKFIsUJwZcCGZj0Mpq+TZmzyifSMCalU3up20nBZiYYI9jT6w
fCcSr9wNaa92w1d7Kn1OPQ9/d0SgdKU/BhIi+gdZ674bBZm84E7jeQbMndkc
3N5WCm9Gwy/Q/xKvISStXKSinH813/6y1Jbth0iZ+ucypb+cecN9gmGrtOeb
+k5F0HSGm+TPBSuJQGddqSrZ5f0rVFDUOdLtoQtcGi5uJFgKADQs3ZMwLW6B
vGBhG2tSCobs4j1C4AbzUPkIVJKHzGkHJGAu2qGIRwi/vcXgMcdyT2rcpPix
wQ94q248JlaQAAbDOh8jnZnmKtKQImPCCeBFGbNS0lB5LsDAHO5RHPPz4HgC
BwGOpLrvSmlnlqE+fvG66o6D/xbzd3dOpLQXTIk/xre0Ds7l1r3qPJQauQMg
iGl/GmtPJXvLeuatConiiUJcw4UHdVcD0Mdh4v5NpUy+8CsmiOOSWr7W6sbS
VZMPoRGXXcJHvo3W5pN9ZoZVwMUsdGPqNGdYCT19m6af9P3Yjj+AVOSlrDT3
yd7/Q4i14gh9UgNuOjn/QKeq8phLDt32saewqO/MhpkSEgGrewROjKh3dsO0
BvCqXTpGJQpcg9qzqaaB4LcxGr4XhEU1DhsVCTkbosh7yMgdMCeoJPELAkBq
ItopJK1Cn7WGnsZKkfDjGqNuUZQx60tmthzEfguXt50Yo2Iy2da2K5v5bgna
uK7wf8Of8mEqT7y4nkamwcvkw3969jkvBoBQD+JLxMFkkp3ZNlK8KOPq4j8u
O0W2fevx99CJyk4uaMuCr4Yjo6725jb9kHr7XU+ya6LUZBI42NlmnOhRWDxH
PcSdOB3n19OHJvJOWBmqsxYvaN2bPdubWZuI7rmUgDgb80tMSoNgcb57rueF
Umv3tC2bzHI2eU131CfEvIImTqhRFB14qv8djfOoQY5k4lxfiSShbck5nW/3
QyO9q1B9KriM3ANkl9YS5HAtriVsJVYm2w6CRZBcMQ6YnbhEeNjuHn67C/Xo
t3K5Ab5JyRfeTPYdpCCyjjn4g7qDvYnRX/VOkWBYt42IkzqCabYu2f/ejkJM
SAQwkaNl20Jo3gd8RiBh6RpsQtNDgnwsqc4bYy9gfDJ6iELfc6iJUdBveHds
8ICVYEqglo5+hrdrJ5nxe7OlXKxRKuq6CXphplNi/lFF/wFqt6GP9ui1IWgv
s2A8z7US0b1xjRTOBoi9Kszq+Kzw8Ux3yLfdjRgX4MJ7n1N3LNRbWoJ6MeOx
ktydQA1p/pLwJKp6vOUXy1XyOWPTiiK+mhLpbSXKEXYBbtciKsYiz7ypBw+2
NYnjUUqCcZJ0nYDm65cgg1Gbp48Ro3DFLSdWLmRrjw4jh6J4SWkt+5Q8nNnK
GkM9czbs97Y+mUkMAEGlCsBMhZ4vl9P+ZDEWtNpm9obIoEo+c6FsGHHPvpZo
ZqGR7RAZqsI8mPp8qGoVlMliGF5dhyBKqgbUfbxdBLUT1N/DFtnHJ+bR0uKU
xvqVucXNsw6f/72ycoYgyDMDsNUGSJwDueo4jVl9LppQJpFKVQj9BMAfsyJq
ikuWjCv+HG5suMMl9DQA0NHFuOhJnZmtUYCzwONduBW2OyD6s6RcjfWVdGC/
Y1xf3eThdiNkwPuRnLbH5evYwHCD3vUs7t4ibzdO2EzZF1Ucn/i9LSzwpMcV
SGusIbURLTrjwV2iz+cBxvVUDAG58pDQ2ZoYcOXXN05xFp27MGpFcVxnY48R
w0WQau1s0lTKnuRsHweEGMmoLMISbAyU6Rpll/1NTTgWqL65D3YIjwcgUNJp
XiueVDQ6xfnHmILB9EBoEDpjZzWALmSpGQszW6s6r6nHoNUOLYTy/lkNXrFR
pZOxjon7oYGmyn6HHf59tiW6FvINw0UwcP1TQ1R408uGs9mswuglkrdxrBZa
Z5xhTAgGFBWudoIl3O6fKFh8luS0vXbTT7+X3gfrkzasmqaqoFHKqEzjHTJy
5JNLvAW48p0j0KqGUkrEafm9wZwlGuwh+0Frk1e8lY+j6Gqo80kt8I3iFFiZ
oVXJHc+NQiVyN14w7J5Ilbq+DRZuOj5ScS79uoSHUKH7eVgExOKtIzxyZR9Y
m9kh8tYdBp8zxInvxE69fzmkUGipm4TqRBL3IHam1rwOU2NBmKE9ffEUKWSI
+wyS+gewvPoh5vfknEZnVaYG+60LKFUmT4qXQAjDtX43BAdvn2gMS9+zGy5x
Gp+bPmRuqf5QVp9I4+bw0Z/TzayAvykM/Gy5gbZ7i0TDMlPL8MfYGaRBP17d
OUk1ySLWaCRt4thO6YTaEaKbjG/Tjdm9YVB4+r+BZCPGz5JiEnGhjrOPburU
dQrVPo5lONlsErWfsxV6UAh1elpQTICwskIEK5KbWNjA2dJNbGzimiBPpAEU
WqtMAiAUqrOXJxBQiTiuicoIP8VCtxlQAmLarXKmVtzAs1too8WiUuebmaXP
RnX1IM/3PCCUHJl7jX7g8MlKmw/ELez+1WnG1HUO3D5WAoycG0GWPDQTH84j
hofmn8Nq6qcD8zaP3ZG8c8nGJVCgHGJg2Mvb9BH7Og8ACQYS2xFD1b094S8P
SOqbKmWVIWIekMKNz0Vw6nmC/QErFe5+3bI6eAE0QxIyrr3xg/C0omNOWQW5
PwFsO0120QxmX+AGy2VEy6Si9+oX3ZSn9JGNeZsVk26hWqU332tz0jKb1uHM
L1oPy3cWAQWLcfC5U9y3nb9Rz+d+iobwECjU+KHS3vghC1alm1ItqT5uxHBe
UveSZNx8SKBPORi+sR1s9PKgMzmf5kb2F5/wCdvw3+kLTQtBeLiCVbYYGSEY
FIcItq372CyJk2gIm9p9DCpnJq7OvxUKmrjGrdohIYkY+Us6jzRxKPu7Mn1Q
7BxB5TaBJTitJPhG731KGx+vWLajwF27xnyb8aCKPzUFTIkyyBR6RAiqLFbn
P8Rw2n5PfRDKHtVZtjZhxCvvOJsazHCrar1mEwrpJswZLeOzRn0Z5jHcb0YK
pDXSjqi8wiukw+XeMYPbrr1PfSFoUHbTJtkwUMPXQiTt0o4eFXNP4QWvKX/L
M6FjUQtzHTaIkgbPho7XCgOe/5uXIptb3tLaQxvdFrtii21DNtyLaCkYRcW/
HoHhIwXnyh7LYKAv7pmaAvVbpG345dy6kpNZmgWjckbZ5rMpkMf1tcV5tydg
DN5G5npKw7oHFltTulTQbVIQjv/FyvDPWr5yCcg9VM9BOF8ZUT7pxan+bZe3
LAQcv1eceX3sXpfj5Z9ru+Ox3b9V5Lyn6LJ7dixoLjB+jpBIMqhOCUxXQQYQ
/uQdVeQqYnaQNPwwjPaIxGL5XkYLGBUEqzApm+VYcP/+HFqKLuH8lEa8hCA3
JYAXNBvwfw2si/tyH5WFRBt3rF16Scwk2hyLEAoP+t7Ku+lC77G/EI45Xcuz
A/QU+X2gRvgN87FFQl1gEN77pAz8UcM9Ughe71l82z03265C7pCJecwPpxCO
tGd3H1QKTLURtdlrBvbaY2pnUwqcaZoZ7+wWm7wZC0JZOAO/hMIyMdlN86ik
g1zzz5+zU+CrCLtq4dZht6p47nsT7DhlDZ3Q60MH9o7zRlRxl8ugldgQuYU9
JA+OkpMK9boW4lkwVl+BFZdLg6B0ZWB8FrondQeEGY+TPPZALI4lGb7KyVpC
edJJIs4kpL3xBabgnzyhhGSSlRcDdWFtGHQOas0XJo2ngPOduzyjNeFVtzgl
24gdlnJg2/1RYX+4C1/Xb2ReSS5ogSpIw00q464hHiz0fp5K42Ata5JAH80U
dYwhFAebfPC839XGitwxIj32Cu6oAJjfeQKi0j/izNoQ4iZ1GASbnekv8D1j
lfy0xHW6FKyPclJ/D1AFSZsKsA4jqpH6yxuv7OZAzv5f0jOXph9ndl3E0iAQ
x1iyT88NjZZUnNtWvBpT5W7BOsGEkvBxc/ODTW0dEqyLelIYSsv8JMU8waFa
isryWT5HkCnDb/GLeoNMgs4aMRky6o5cmC6l0h2FBubFRay0HyUk75o1CZ6W
n8lBbdvwyaT19lsrhYyD6nFubm8wF2BJ+o3cg75sRPAl0lyzOt5OY/H8/Hrb
0GZBgC7K3XulXqEab/YrCT6gn83Blh33p42PGhGta4LMLWalMTNF8b0MB6x8
kqj2W+18D8fFKYnWtqAWIoG71Zgoxz5LslFc2xWN0zXApFyuPCY7wwtMrRyk
STTiydu0EHtFNF4Ro7esJ3ZCTx5SOS6tL7p5xxNnuC2Fisx7W082Ku8AESKa
TJm2QgunldziKPkGcps5gPgUtCuVkJM8Oy7NWpZa1TmHetQ3z3kpmsXZthu+
hBZSGwbnNXgXkZJTzbfunV2GEjL3/XGAt2GiIJ9sHFkuqZ46q3mRIAKgG3wY
3tLS3NkezYG2KWiCBpfIwuxFLiBDySu0zk+aHzZy4T459zwukDRevC0II47g
nW5Dthxfq1+1qLdpD9r2eSo3cSUgQO0PQAx18k8UdXdNF62qD6ur3WU6MEc/
pYv1obANr0RU7clzKZ7ENoHOoERLYx2sNI5fAy97K83WwRBPGFal3PSuwj7+
Vg+M1h/bQrKexcKs9mieHMQmxVxoGWVFv7WOknu+17ps8O8lCVYG29teYkxG
Ed3AKXMXVbnomyBKGxIFh2cr0OrWh9BmWxU2RttGeXZTcGDaO7NPhLxkQ2T2
9K011+S+SGZh1gfkH6ZK6Q0hxAPCs6vT+QWuLooQd6E8rICPOjIkVeUfZaYl
OTRMHdm/qwiofISHI/3Xg1GCahZfgHwH24D32ZYCkd7EB8cc/fGdmajElj9Q
4WU//IacYtmVvHINs87G0w4BWpKl71jPVuJR4aDfLbi0kFsRscepwNwnWyST
vdEEM1VYak8MuUFAyG1+LMvXH2/uFiN1845ZzB0rK4eJ1NDkOPkbfxjn3eUQ
fG4tUGO/FKBybsLj4L09TMdfGqNhuMZsBu3XHguAzsb7TWwD/cW5E+3PnPY8
juDJyeWIDQnZvCpFI3tWHKvQ3j5ZLV9QjtCyend7GSGUax5OZqVi9nHYgLfV
pcxxg/mhFXYKd24iUHIkJVFAAJM+hWvJvqsnBobtO3l7sSGiKZcUT/tzuuN+
BOn0Plo712UGVLJeG0eckWU+ig+EStcUCVW7Y/9mDIV6+QWu7rGPScuaZiQP
Ci6V0Ah8RxFURCgLmPdxCwbP01TZYNbqKHMiDcyizhiwuMKcxRq62qfyltgE
NpKD6j/dItI0lY76zzE/inMzlvDXn8ZezsgitE2ko/gnEbgsZWq0LK3/E4oe
1YNBjLNkJ8xXd/8HMrgay6IQ9spAt2KVAa70MYhWgo380c4Wp8vEdNSYV34p
F+Rxbg8gdh94BtH30Qf7xKrl4TaY4WxUaISxL0MtXgV0+C80pYqyDn+UXygC
M4TThbMmHO5VaUfjKlJ2VlVzfBKyZUnhXkITdZO54cX4J7IWL9ys/IlwbJ4x
OcDvi6Fa+NdBGoCI/nPAbMvflGEBJR0SsS72anyZsJ8/nmdCM3odPLRwkg/7
qqJ2pq2GTIFo/qA9vmzVrQS1IFcCEfxx1YmCT47+41dab345DTKz97l/x1R9
zwVnK0xQfm+MyAK09cl0NwYIhm4STE8suoQPB/0fhUVBDTXkYquW3+GDm1Wh
V8wHxTefDgWsLLpLzAfyYj7CyiA/Uq5UUgUz5AqaaTdpo4sP5iiM8gq44eyH
XiHUSnUROGA8VJtkNYS0BAgFUvSh44BRdqUajhY4Ql0nuneKXoKujITCCkCW
JZ5BFhCdNAZ2qHfw6wlZxUM/PjdBGTEQ9klkmKMvj6icS0Nm33PwYBCKCyHB
RaCn2p404+9rT8jc5SaMEzsgklrRn+3G2XJj9bLqQ07RX/wZns+bxS92eqhy
4L6cJelsXtrgBpKr0g9iuKkR6yL/4jbdluije14hTnBo33ZMGYF3UHpu4j69
kzUAUPDFZ60WtVO/xpb+D5FMgR5KpCm53VwWZCf+eywQWtT9uoME6ok6Z+1V
uopeu/r+a9z/WbeMCC+uJYgP1QBmw3CvKVNepjpm1CxAZfZOIALAZYzQOFZU
Y/wu8+G/nsj5j6f0q+3FYb85AlMTmV3/+zZY7bxRco6slFbQTG1TR6spUTNd
UQ2/2+Mzzs3GWFkt0OgnGgLPEKUwJs6uOqTxj4QZJFJaaiwYuRQqOD+tksS2
n4FvRn9O/sFkGMVcqv7QTA8GvdthiAsaVVo40nBKy5ZfJWjB6BTfj5OmsRmJ
QZSBU2eOe1inOUGQoZQYf5LSJRnIMt9f89t5vLJ83iSV9fbT3jcQFwXJubVb
GQqLN7ek78DC+H8uJpofG+Bzd0V2U0jhiKtx8Ocr1ZbzT2niBiADikPX5GCz
GyOQEBSu6jh6GomYSSIoTCy2STn19PrjL/bmK309hT9RCQQEx00+H2kakCpJ
SorEu9axnZnMcfnvvuz1nKXWi/Mc32vzc1QPHSfRzxm/ZNrZ+rQtRCVjRRFd
rdazxRhXDPKjclFIn6HFLPk+Hj3n2HVje3H3Y3W/ecvIwVi9zq8XB4vNEsdZ
luRBKqA/wCuyzo6tR2CeTnYhoj6cJGNKKWXDUI5G+HaH8YZ3Pe59Lnt+TMoH
dMX8/uO8TC/k+FIXXKgTbyW3jAVdyA0gPlLXLok3ncDBKHE88AvqU4Zmxmbj
FWlOKPjEUISnCsFEsfYfPfgPQ3ul8qO+UHPWa6EUP0XhOfrMqdjZpMeJsYgx
sPs1cBJEP+iXGtWzIBNZ2YKr0is8fPjgxBm4iDjF0DCFaoE3v4H0oSiEv8TZ
TC0EV3dGOqvtxqmFf/+C9qPKB+crHO48Iyc/i5cUuAFY/BrgwY+hMTFBcMwE
M+NLKy0ph9HE2eDOUPihx58mnYNfs/3XBuKrPCXgDI+so4W8HccXjQAxD4Q4
B+kj69AxgArrzWjB+SK4TIppusgLaNf9PxNJnMAR5Wuq3d8chAYPcslW4aTm
fQvGxJaH9ORIeEPmbHzRTmP78+dKRyaARB7IuyESK1d8s2CpWdP2FwdpM/td
z+ScJuyddzgCY5FFKKgbD6LiaiOl7DYkbNXT5ZAwtCIW3HSqeYt1zqii3bVB
AanUZ/x2w8t44BFXhPDWFQBAjSBwlU1FnXsEiFxdOcquqiZWVuXocyhxvP8/
yURYtnsV+um83Fzj6kTtvpmtKXteucTOEGx4UfkfLcu2W24kAe50E3E4BddK
bo7IJPBKWJS2SuBa/dNh6TkSSPQR7SQpefUs9EzkAlZGwHp4p5ckLUyWbL3m
HHZymoPrinuAgvzVEbHxmOrXtTBED2j7Ik7wJsIj0VZV7pkeZuLhZuftQg/C
tzVaCdznOPk+C+EfSvoXyATUkECX+s/gBwD5UCK+P1B3pBoarVvnpe1E6tTe
/ebNo5xPYEH+HLa5GGVAwmT8M4GohHJvvWjp13c+byVpDf/dWPcjPOHxuSyb
Tb3So0cF+QQVLgAEDWyPKe/J/srQpMseYLAeDWTryj6XAnYXDtKRiEvaiQBO
C7WoZ6LWRbR0PBGHqsMsoYnf9hsKCYU48pFrCHpoLu4KXAAZBhyX/X60H+/g
hEIlPghhqWNr3AaW6o/wvZ1w72Xv/KyYjgt7rvjbii7xxcfAaRvUMkIv0w/Y
PM02FvvdMINcR4lcysLgl2CLAyfUPk6OLkWOs2XCwykE0XpAT7LfyR8RXJzg
JPt3UDT3da5+ePibNFxPV1uDpmhjtIGNsPQwlis8NCYh71CAVfbSD7CvxolC
DzZLJanEJmboC0Bpme9UlhWAjyfblWmnduq0WC03bkPDoXlIu7we2TU9mpf4
YpTHFBBIYfEFBGPde9KKgpuNXU0IwISMZ9CAMLgV/E+2N1CEZqb/6iKg5m8Z
Bg2SrbgTIWBkcNzvN+IkDsZ1L2VedobcD2KunXK/GfskxvxfyBdCejDm45ew
FF3YodvW3FQevqDRnZT1Ay8wUARThuRx1wXbCcRpIGsPzpMu3NcD5SAnhIrd
6AqL5bp8Kd0ZpVctdtLDdApxmqwKtMvW7CTCA5Kt7CNHImFhcv/l/9VUKroo
AzIPRL6zK8blyMyxygsOR3D75j12pBjzVgX9A78hakxoDZDqOBDvNE/1IKXC
EAUuv3KsgmPk2R5HmRmGjfPBeLaFUnNP9kUDn3bKPs+miK3kLWjYcDBbv3Gy
5SckHYeSiWNFpgdVkR2DXnARV6hFd5Lk1t4/gYEqdFfjzXVENBFrfca0HvHd
5b4a/r7QHUeWVEKx4o3NtRPY29myTOvJ7zP9X0mwBns8vqEl9XfjtLE8Z6if
igM60rdO6Po66k1kdDzCtv8kKxF++GkltIpraz/KzBH9EsO0qreOFXkp9K6Z
aMpaUleXN+AeJVZGHc6bitQx0LnOgQLMic/ZiCHl98OidKL23/TBLZnkWgom
H2AwYmk+ZeS4QM74QFaVh/92F+25flQlmXKCRBoOi08gpCOUCZFFZvXzKQpG
UOOCg0r2nuGoBOO1da/d2r7fG6+c2equwibgsA6a9mIrfrWSICZPd01N3Oli
snQPzkQBOAZXru8LBtGsi6MWxnMCM2x2iKxrXSbh8CuFj3+H7LxbZXkUtjlZ
QFtX2OppPtaNec99iOdxCWj93n90q/pRqqeZlJRzYNnTPYssYDec3ZPNkd3O
fJi9mVvqZljqgDkN75VDt69FYsKb5ecaBTMHvChiWkHQIJGRL+9vyTHOry7c
qpgAH9OaW202gLZkJ7oxU8SvoCMl2g/fOT9ks9j5n+s5KWnR9uaYYJjk5+sz
AHyU++YpXBLc89yqfPpJL+uyE0VwRxZo8GPqUMmiVxUat5eu8PUTm6vmZQPK
23D5fof4JuKuJpfZUrnYkMuUO6GPzNKMPOlZ+IYpte2ZtDKV3q0JAgqqS38v
N8plkO5zWeWFFNsuLdM8541dFnrbMcx7Lf55NV7Lw1QlEGkDqg0rM5mNrlDJ
FeLW5Eh1xj4JnMe1SHszt0JhgXdSJtJEb7B6scNq9xcCTkjGEZ6qPw7nlW3X
4FVJoO+MMhYLH+kzMr16XJblqtjhgEMB13MP+eggEVYlis1gYHZdHtUBaxH5
Vuq1dIwN9t5eD2lMlSl8sTOtol181T+JvgaiCfC4epKGaU6L0KOrDNj37xkY
NWa0hrsmvxUoHgYbi9Mw24R9SiMHmNMmWGhhuoXcMCkyhFI9tHlRx4mv9bpD
cRfYqIXD4jSII+wd+E4oIguVByAceV91nx1trOOECNgnlHo1wII/VU0Dr8xa
yaU45FvH2K+97dwFivRqiBdINTTEUQrLCaQ2ue7RGU4dbFD+3Ihsf92uW0eY
P1uqgPojaaL9+sPXWp4ePlqwYlPE+euJenSTNryp2rwlqg2D5Lv0PUKGFKcZ
xftww8XIl8DqpPJ4LuNX+fvXreNzlCyhl3TEn3g9/Gz9fS5sDazva3BjN6hz
HvGVLZlPZIzm3JaMbd7E2Mix0NJ+3REUHZl/UFit57xEkt9m9hAHYhfASdnY
LBC3Mra2Vfys4kOE4o6Ecte+fykIcrXRrhxgYKFoByew5nCb6LPvVg5vEYV8
N9K1cyibZO6BPJihqofIyt4ZU4Fs910TKELVUDPU3y08lYsZhQCEGWsL5fhn
bRkorxgSk952HRqV4T9cABxLSfoD4qhcgCq8DVVyYaMSNKdEgQYMakCqWAe8
uNWD0eyWp2z0teMsW3ZNDx1bSrBPT9B763brp2P0mvQroMfx5bRrROjDJ0YZ
J0Rgwugfo3/Pdn4Pl412p/XaNu6q2TxQQlK9aDmbo6WwNo2XnE/THHh02P5l
PQEF2Kh0zDYkZBLJypvYh7DmyMGXw2/VIzG7WpoPo7tGS1NTm1cle9zUixSS
R6t5ren4aubOcoBU+sRkZco3GmfsrH5fgmd/t8dcF8VRURzGSQWJuo0A/mQ8
C38a19vy6fJ8IePlXHCUJcFU5nHKx8c6RiMRRxLse0zuNZNab2yiz1A+KjRe
kBcbFeWz/UWfTeIBL7q+XT/VbMbpW7dsoESSHgcut8WvHAwNrrKDsIqBfTSd
h0q9FswyVeyk5ZxEx5RWAOHJJp6UWozM9JF+zgY0QLXVrlv0Pc5gAAF+5gCS
wuOC1kMx3TsHETSFpF4E7+ycDgOQBhThIo6gGw2+C3nqcHHvFhIdR4IRVlom
YgcVCjbMrzEd1oqU9dgfinDfdO4+knEmfCVLw2DhdQEXwVD/2cP0yrX7DcYi
bzW8KR9cqaeidbu1hMQDUrc30hBWxwpWrBWyJt3keEl8UXDI2+CknqE2WyR3
eP+JbdFtB188p6Urp8DDDJWP2voojB2CHSXW0g/N3vj2HGASiCvntM7Bqwfv
inVRFt4iweOCNVV/ac1sSuGEqt6H52sYb2mCD77LOndIJgmrxiCjD8sUJszI
oAydHTxB7Bl2Nq1FRe0exnV5FxOfsyFGyn1w2avAJtWjP1a9VYe3WUuY+9dp
Ks6ZwZ34f21Z7nLMe81y1hoWk27fKKyVZuARCiX0QdPbgQxkTY4bDi1guXCa
cw8ksJT4LzNbzyfV3/Z703vEDmdXQz9b5X2c3Ns+Lo/wskzqfZ/L+0OY6PSc
Bk/cRrJoIzhKn2dy1XsYmU0BC9PZdwPQVadCwpbA4ro7C+31SMlZCu/lnJCZ
H8SuXr2V7FS6JGCR95xJet/xS+NMz3P//zGsy0qoMHSCTh4Veqzl3hOC8FAO
kUZK+tWFXy5QUEo1BqOcLwm1blzJwdGBPtEq+dftRUPxJqXAs1IuExpqBuin
+d3X3OKBLRyyfij4fOysGhT1SlLXY53w+mq1A/5IAFp/+rpW4JtG/EboHyLB
fviaDCftKK4pBqREXAhCwhRjj9uY0alFMySMEjiueWa6qCJRrMYptLHNWSuG
/inJdTK0OTTlqOAzbFxqUN/elDFfVioogTokiQunKOyVNnppcU4oI5U3+aPd
VM93ATSEBJX9slWXmVPKCWeBeatlL7S502Ieb224E6Dai8SUrrqJ6FL/X4Ns
Ypn+GmvRf8l1nHSP+cLgu+RyaJMjeJhQPvT/2NTozgmDqQtTspmnPvxQCnru
p3PP8OzTLVYaZRi7yDw5VM+TOklxyheIX1+zO3W2ypEbSe7pfq9WlmQCdBGA
TJ+oSxa+TKhybCSQ2OlB3iHnBqD9RStkcRJ4jh85dhRukuK7AQX8IOVKKTZJ
chK+R7p1zE/xGsSTf/QrGO3Vu8WljAhoIVoA/XzjU2/y4wcfgOmt50kfqX/s
eHFKfjZRXo5Mb/Eke2hdLySxg8z9sdtPOQJZkApek8rOfiQqBFmjerFFpOu2
7YObJ1GazvQ0TsGluJZCFzFn798+h9bt5c0eN9ty5nuQV9gvzu9P8/irxPlO
17xEhLkofxgAw0fdEMX7Febnmvauw1RShDZ3ibPoVvXJLBXP/yXmgZHactrV
ZbbLpMB0bs0ukrrPxoN+9Cy0g5kmZ/ZcBBMBQ/ZkkAz6V1ofdz+t2DFwg7d5
LoO/nLLv8Qx/W4VxnQRmWp9wvCdKXQiTPAnuG4oz3GVWnE4+qWR6ZbcOqhkv
Rg+LWD13qCSCeU4khgI26OY9nsFsjaeETGzjejL9BRTLjnmJhC6G6By7zDSD
lh1DghzY6XKN71fn06thb3FkJ6nsf48dfLtbwiBWcFdexIMF/NU4mcNlMRiG
1aHqr9tJ0W4BRgG+LTCJtL2J+bWvOLeaOG3vfQmBo5g6LCXX1blp5OluW5YW
l+UbkjgqLRIc8is3op2FjMDcNqaoCzrxXgxDdgNJMG1vcoOJwdWwm8iuVtWQ
JsT+z3ElxQ4+LK2+ieBSXR44omCKT/zzSYMbgg5vqzqDNDLgGp0dWwqkQ1gP
XauuyGmJWvwXypmxEX2KUQ/neRH6/mht056U66v9gGSeTDyCJsJBvdlT43CT
/M03eCxH1wO5znHVKTNgxJb/3H+rFgIm2vXFcINwYoAkv3dN0ekXgeCjNDhR
+E4rAQk8MMQ80ASAujYy2SzQx60tbzKycOil8RpjCHZm0va2LGbbfXtYWb1U
3mp5UupT7jrge9rUVLwHW9pDSRsyy4y47i/zpJ4NLIoL1KLX/puTelLhBlGI
EaElCkSUTaUF1OQTThAs7stp9Sf/3lFAq+15x2DSRY49afJE58ZMsMLMHxCp
VNTopsdlS38VUech2HwRF1Rk6jnqcFS/pur39pik438tmqyNG//TPJ60dbxs
K95e6E/RTb0RK2ubsJTyB6GQR6gN3QwOG4DKfn2vSCauvDIFGlbthmRP2El6
kuQg+TB7R9JqdC+swJ/zw/zEC3YKsm0ivWHwBXLpbcLBXCFg8bssa59o4JHn
UYOj9brmDxcEtLP+q9vXfeMF36V+aAAKHqZNOGlVT+kUdDWX/dXKaKgJqiip
v1gDwp/f+P1Y/OvgZ4XN3/ZIONHm8aGtLAaboRvzBiKAdGB9U6GVWlAQkM7p
OXNC/LE6nRxQxSobUuub5FuZocwzeCatHrPyRQfl7K5PAdf2uww/c7n3kDgI
ih7rGBLbvBMbKoTHNZFyOvRpBnqKPYR0pbwbGBcK4FVK18kmKtt9QWYuXhv0
c1+sshTfoY7omwV74LsHKBy+ZZIAHtvSWdtwNQPMdRrUnk0LwyvFHVCTthha
Gij7UkHfO1jbPLE7EW/kw7xAcn0MwBndChDx1XI2q1HsgfkSI4vqikrvW7On
JL8baqP2t7iHhgNoQfBtewrJAU13FTftiANvTSfnAxJ5cob3B9gibMW1+YTm
vq2LttP6+OdCZKPJPQ8b/qViWaaAKlI13ukYre6g89h+VOSztlR/nGaWcJK4
CF+bI5R9fxbLDluUvq8bo8hUUpvsp8Rf2jr8/BqV06J4HmqJqTUDe1ldyG8Z
RP69IwhUgFsFFV8dRe+ZfxdvBV/3TdOn9vwJ3986KPa78yUD6Yp1nGGFWDrU
YYi/zcIPJ+V9dzN+a3NHURManH9KD0ydfOGKlM6r5S7kypoca5UQc24OXQ0J
maJFHN02GodQ0TMqBLV20W/IBYwtfscIrsQia4LC4jEVUyN0ntCGXaAlxDX2
CUXup+cAnEdk6wJIr0Igj2BSQ8YBSaIccR1npMFhwHwX5VOGw51r48CzN4BF
pbbek9ZEhrLJb3q2Lhbs+DFl5cmVg/zbnAFd4MV7WiDO3QZ2yDWAkqOVS3HH
elCuK5W2wfWTXYwaWHesRSAmJeWwo5J/ldk8+8FS8+YNc2Cz+HKnTtjLFam+
+BvdiPzor/5FvY2SitoJO0EorGBZZdrA52g/t8Hppd0PAmr1o4iEU8sMw3Un
98auVtTHzxQVgyhKtnzyNCSB8T0J6eqFu1Y15ata+ypHuUWNugds7D5SiqaS
UvBqrXqc69DvqJVlwDr7nWpJ0rry4HHRoj4NqW/upTFMqVccYFAZcO9geaMd
Jyfyuhq80bQXECDlYsM/DpyEk5XVuClybehXXnZ8IKvg2tPGFpNFcy0f2ENE
ZHAvRIG+w5KuwMNg1mUV3okOiWy22V/faj/ppZHj8wFj2tmpvoC2j0DYjcmW
Rgc7tQMKQsgseiF6dpHzfM+ZLuorlQl2vTO6sl++Uixc8UFrTlL31dVpahR9
g0kjFjUaFzkUGGVzMonc0nnFWICaDjSYX+XImZsG9/1VhmzLs9ZmmEqkVqCw
FGq7uvrOhzplqJx2Fx7yMfmCMtLom/eZ339xw/0x/Ki1F4exReiV9cKs2WN7
xJK1dVAPx0rd3+XtqYvrK77Cfh+PgBOtUjNi10h93s8tUbOs+/3+6zzR2kfT
t3y9QJ6XT5I/q6H7Git8u1L9Ti+ZYwnCi0LOzzEXmQYCMAGc3VQRI0/MXnyq
zbvVmu12+Gh7bl8wHkhl4Bafpa9oQiuyV+8Ycw+x+Hlf64yvj6Q1127zLQC0
WWlqBBNu5bH919EzQfNsblp+cGiDojMt0nZpT1lSOYbu8Ssajge8N5NawK3w
CsKQhEmes5j5/rhW2kkT8K889cnqOwYQ8bYAywjT/5+Js886nJixJJeK7LmP
j0X89CKLqDfB/vSwH3p3d1prznw5r/BNWeAE27ziM3zmTPdYMqoF1AOm/4HR
EeLqPliPKOXIplIN69CdS2L2K7fiQwBlHYWSLlPI6CM+eHsa4mPDOxsnLt0K
Lw8hAwBELjv19VBdU9T+XoGk/Qid5LoQCW0yRQzT/i8G4xMjhHVhs72dce5g
W0TN0jBrN1YMSC8I3e+kMY1/OggAvVeFVhJB+l7pRflLYj470by0eiCWeBLM
rulyUTHzNCcvJQbU3+xDXxUu8YSvZWEjWSu8KmqpbWzqdhZBJA5BFdVrLQRZ
T3KPkO4w4UmwH4yVyaEzHOQA2ZY5dVfbQJV090zqZSFPpAa8Q+6hPDcgGihB
75yu8jaXm3rUBcQ0fPxqRxoAr4e7rvkuA2Zo8MwtMXMAdgwcBz6O6YiRJecv
JoKlnzzdTSb6PoIlpNcK9krZL7WYQehkruSHbGiP+9072uab3b9mkZzzrMiS
1EKUPhJ5JfNmxa7wpmUITzHfVoypUZhovLymyPz2LGXHuzbGdDYfuizIXXYH
3FWt61U9ExydfNt01LtMtnWvj8c4PmrWMzie+tXx61D1ix6Reqt2w6zHwObM
Xt/toTKEMr4ocqS/aINqpaILMLGCZRa5FP9NrvKX469CRu7sMDl4CcwFU4nm
VEMdRdgYE4BeTTNmX+B6eFCabx56zXUxwHjZrHcg4olEyuedbkp16kIwvT5s
BwBcIbsyCZfDhNU92z/JfFC4SdJCsUH0ZFAN8IeXrSMIka/kLP/VVy6xHuvt
/MkKg4E3uqnOHAYJlKeNYz0cfFWUqWgm7eOxeiFDQpiBnirmgjZwl2U39O3t
hJDDf4IALyPqatOQ/9GmQjZc5y5xeWnucjQ/cXItdimKchRTIL9GvG90M64O
eOAhYwqniHq2QG3ZaBxAWDtb+HSBLAD0lTMn2i+Dus4TJStG9xqN0HYuU5/v
r/zW8OAHYgWTTtx5VZ38joMl7x3PwRZkSoq3OLDYRpNUzClBn/b5o7O8C1gR
qi33bypwWbMAbMY/9nTFpr5lL1yex7+ulQE96VazLgRQd6V6ymxs3w5IfE8z
DVKca3hwGKUNIn6HmVgdUQGxy9TMEDpQEo1Apz/EBE1wtWK30TO+UuWYFuoM
fqdDBPiTvg7qnRlBWOfbTSmq5vZuq0CsjCFwUJn0mp9I350ZDpSoJmacz5Or
MO+rgIaU+Jr8Bcj0x6bAx5s5KQaPWzM0eRPsiUaLCFBt83vbpYpe4qq2B70l
2vnqF9CCUMfRAnwWwKJXZ7/QUKmdZPFfO/LeaXu8yLDG9mqjFoa7tSBUcNMo
hSFwoV7e5AHEP4jiCoXqIGrl0tmUQd3XPpc0z5M/vvmb/pfMWx7aJZjBfz8H
au74DRaH9TXo1S12ppvbqcDA5J99Tn/+lSNyQi+swREULAubCQnkpjff/GVS
yewpSlQCDFNeMYg3VMpVRiGctArXDaBmbPjT3C9fL+M/7Q27chc9n2bLsBcf
CPF2pWEDbmBiNkZEX50LvOXK6w2LA405NIXixR2LSLQKwN3+XTyqONse09oZ
ANIPY0LPJO4icqc+KRlbQjuuMRQUlTuehoFUdQfM07iU8ocnXuDKnX1Qk1yF
mNz9fc9LTU+ym8lDL8+GFcnTcybVRiz7i+VURRPBx6L9C1z1xoyCUfsy7fJV
8SU7qXQQEY0lNSjLePK6iMyyS0SFm3sef6vwtQACA/87scG+VbuG1qqcz7CF
HPATSKULFDn1Jxlm4tUhdmt9hypDDgsfiS1Fm0T8gd2OJcHvFIvmXNMC5POH
ge63gwaQNfkrlmI68wxB9Sm4HwbANEx2EKrSOKEyw17KVg6wsKQRo+Kkef8U
3/14Xi5nZ2hBweLsAg3v87P7W3ShFK/2HOJlVa243L1LRAzsGx97rcDyxuU6
M7PdAblBW8yIe2zqjOa7ooBnOZyURyVX1uARRwDR1nZ1BHwcXSjlocWo1FQU
0sUACcTKoA2++NdOG2P7UGOy3+Bl4eeyFCCcZO7GHpKykcczS1+k5WXRnDj/
pmdL++xgFOtwtbYYK4RH6dq4ptCToT3j3GV70thOKHrC2vZtKXoRsZli3hdX
srAIaJIFuO6GUg3uhgbVz6mJBqyGjqATgl+ClslDO7hHxs+9hc14Fvzv8xaC
0Hp1hFZ20u1t0kK6vaiyGo4fhpg6XkMKM3M2GnHlQCVxR/gAEG9BFfrtzW1T
t+u9ACCSY9koP67mO4AvQD6HQi4V3wdnxp1uEn3gySh/yMoUVKWGT3y+z3y9
TH1SNK3GjVuna9of9qiglvlteSHuzmsmkhBKCOFRy+WqLL+ywNtObjiM7XEZ
o72qR7P7NUuann2nF1PWtaPODlAmmqAkqPMc0iHa1zZrgFyV3RSudpSy5WoE
VWoOiF1SwcWfqul9WwvlPSMqzhvliLULUKI+S8dhhoYQluuwhWmC4vw5aAEx
t96gWCtmkcvPJS3MdpJLrjSFcU0Rrl5vcOigmpx7AFJmYNSwrbNL36LC0XBs
o7AW7EdIialKzVGGIRd/7Kj2xXqNC9cUkURy++k9UzPmYUbyookkGcjEp3SS
5O2z/7zrNKLqBes8kudP2eS0H9biS+uIvEkARWKtckLmiZmUWO7k1T/MkYOq
vZyOMfknoOjXN5dkiRpovLVrL4RWacpytPEUbZv3ALKFhVesPHRNVRUjZXq/
6FumUTRwuGikdtmiDVHxtyrEmU7zvCR28opjFhdkSgURhdUGfDRmNCDh2Iwg
irYB1bg/YcsqJ+6803N2g1IXjgPLOlKdIQoV30iht4w2Wm2BszD4lCQanKMO
kEO/Zfh/u700BssTRWScmaCaq6/ihd8AC11RReN1TVsRRDNESNOziG9njmOu
eFrlrIAlJkBqK9taJHWX7mj5gX2SLjpRs6ZS7VlGTUJ3i1AdpPzc7DHS/+KJ
DkHAAuOPV9qXlr56QiKpzRpp2sJcjO0FMrk3ENDZ6jngy/SKovbyOi1Egvz8
CFbfKezpmP9LUQv9uPK7HUWKKl1VcDO0ESlyjdm6zMbV29abhTBkZt6JqlRE
EZd72RiRr2LP5N24whGksRc3FvMvRK51q4sjt30WRwtNSy/b5ycLK8aBSQiv
O0RLsB8GgCHRSoaXidLdhnK5Ral5wVXdqWXh0K3ax6coSZaIoD2cP79tCQU/
RCNHqzU1PjSt86eOc6AJbzwOzp05QfMMKzv9jakmbzknWnwoASo6yKzX5RFW
sWDGoRnWeRd/9Sra7Im6E1Zp25DBqShGH+los/uJ36NSdqIAdNbCagCm5XKs
g6XNvDUIWj+YBlBlJLJ+KQajtd5VD5HP78QV1+3fJb2VmB0Y4dyAE0L507rD
Pg6aTYgKODyVhIgwrgZRubrIrPqpoQhJ1CY2szuALyo5clyZQxwJrphyS08W
7qklSe/ExsEUtK8pvAE0ZumoSK4AJ28hK65zRY+QVhvLvuWFxkJgmF7gQBHV
iSyIXulqGdi4L+0OvusEwhRPRicFEO5x/aqxDq8Th44q++g6amdMdzMD+tQL
pu9l8HBLrzrbJ8I3aCAkyFElFn6vu27ZHTI2VSRd2MrtT092U7/55qAU3yqQ
orO6Kwu//cpA1vLmfNtz5ITWRhhshZwZWpeZa0/2KYxZ6b2n56K0rnuo+XGT
hYzrAqAieCowX8XOqCVw4zwXvO6ntQVx7YshYDwnle99fKhQiPtb8MRiH2cr
0fHVAa2rxuIQ94ZBNnq8KfN+2xLsHFPl6aACuORB6+hz1LqUw5fPiZuPE0MG
xrkUY922M3U1pz0Ik57q9uLVIGwM1KM2w2Tn5zdGAa+OA/RcZxtB7r7cuLiA
GMSx5M0gI+BHwGl14bEYRo48iaQfngeHvwKj4cafCuNkxyMZZqDNiyDlwFRt
FFgIMSSQKfndFshaze01ovQqPDjFAIP4eIB0NvIEfOYZNqa7WhBISVAqrgMr
x7qoOgy76t858p6u6X98Q/wIFHMv6xIY+ZZdeXWQShJF8FRxpJyw1Q7P+erm
knV4uCAI5udZkC4wHYd46D+om+szS6nA0n+50N7+tOVs8os0wXTPwBgScTU+
zS5nrGh+tj3P5ISEUljDuQzmePOcmGaIXwt1GiFqGjsULCE5TpYRU3Jjk3+V
mINvrjEZlMB7CwydG7yYdqp17Gj5a4p7HAVbayHDacNF4WuMwQnP15VihpMT
yr9oTI8g5JdRfCEQKhbXVBqwGmQLQvlhcuH7k0QR7kVvskP0gPkbMNxsYco0
CrnuMx0tiZWJvqS467DBxFE3vbeITmbGs9BKx7FOvz+L4T4M0ALq60ECeTNB
/yPoAMvayQ0V3wgAWUSTobowBp9t9VZNSxyQDs01moU8RGimX/L5xzM4NG0w
B9+P9Y+2AxPtrjhFEeK++bB4qoSolGmhZn1Xg2rkqBDjRjmj8mHUG0HYZJgN
++YBnJJcYxDzCiHeqST0YDEmPplamjLhA+/CUfu9WL6eKV5wFVhQZsbqEDB8
tZ0Wvb5dHCRkQ1vzkY0/xi92p5pBIykUxEv5n4A7cPhh3fHOKMHDjzdn/lpy
J9EXQ0HRZq+ztdQqYQv7wwPxWcQdjVvyY75U7ahypNEcD2n3J2czpLflGlnd
AQObtArO/0pztHU45Ccl/NKEtJDfPHUeda6GmMsdQjgWOo8Dt1qrE0Zk80w4
EmIbYS3J4t/ukQCRoS7xoGpuYSHm1wS5cik3jX3SuITj1VuIL+wG02FeNrBE
9LKNJefBEX0kLkyb/bSt00IgjhHvYutC0Gj18MN+lDMr3B8Du9EK9t1QwC06
ppmsWu+9O5Sytm+bJy2lkniK2Y+NLm81C+0ap2he3ch24smouuAYyIhcpWWw
5sjKNQQv5vwA4PQJ5xysDk8bJwExgA5TI2dM+46TD5tvhNCZQHfaiQajOQYB
8/SqeBqErdSOZkyhdBheAojtfyep+nHVqLEEWKtWLNjBhJ266/J8fGOaU+fj
o01pMe+wvIp1SsBV88C9OWEFcuEO1Wuvdq4gYVhmWmB7ePjpxKAa9vqj7eYR
DA8dwi7gfbfZVbp217Ab2ezEm9TWqDjXex2254Vig2VsTg1Q//zF68lQuc/C
cA5sX2VWRKlAtnKKivrWlIt3HtmU23rhbXOWPctgK17CyzTjVzv/A8m6WMpS
4JwTHiFt43/9eYmaXHc+4qAEKIuE84d/V4kIw2uo7Z88a0tx/BQURQ2imNyB
NTErg8uSg9NhsNvbcP4HRwn7qcuQs9g2G1n4QkDJVqGQ9kugM9EwiHn+tZdt
D+bN1dM6yr8q6fu+ixZiG/RnaU1oLrQTAS/MMW9jAs5FLXKIi87JGqQFZQrA
woMgskLuLxZOcOprY9wY5EiV4E83FgrL1rIYOFAV7t3Dj+SzcVUhUU0aFcE/
aD/27fw5TnhXYWMU+GsQ2P07/eFmbtDnlngcyuxVZMII4roK4WcTHIhArrNt
4fGg+wg9RRofCu4BOAvs1SYP/hbyhY75iojvk0uklgD1zPaHfJjsioJSxhF3
bkjlLpafC8ochYmkOKXMyed305oTFXG41ap67Os0v4ZN6IZKbl4fRkATjsZ8
R9y+64I7QUlBlRqH8JODwrKBgDeorRJF7uJ51JjJI9ZiC7mkfsiTn0yRaLew
5/fvOC/PqE0U/vFmuLLfXnKxFhC4oixTK6PoDeJpdLxum1zme6KqEpYlLYuv
/PiqoYOeTThxERPYDs66Hy0m/oAIpTxyvVRsDT94QGmdUklCaaZt1FWya96W
cMH+RKRNexSghFZZ2Ldk+atkHr87pP8K2/YeF0oohLysMPdxtQR7p/Ry/jpm
PCetsEd/3YwWz84bOq5hpbI7QDADvuT/slig3IwK9YgTgDFDf1GMKkmpWBuw
iXFusYXKdxvSznM5ZZLdEYLmYydAblSG8s9QmnUThZ8t6Pry+Nwk4CCa274+
5RNV6bD87Ava51TGJ5GFV9YNUcJMjl8GaMMfgOa6kp0ZB7XvSftNob6OOsL9
IakiPpvc7Zaq83uXfjC6eEeMkkWgEIYf2cTObtT7Gj8CIdpODxkJgoBsnaaa
+gK/LDKXAoeJxc/LND2qy5XN9GkN1DMd8Fcaf9cewaMr4qsJjCw9ItnkVegF
N+X8i8HyPHxPqtz8L4ENkrgyTEa2lBYJ/wlx8a9XsGgMTZvD/N1w1AyIMLdP
u/JD2pnMt21WsdzvA6TlMJb5232awLNF+DFL2XGbGokpDpF/TYMq7yfhvoWM
2s9020yO/C9Qpam2bN31SqWi47ad/ab0iJPEpSAt0Ax16HJU8Z3WyMEmil9G
YtdrqNqIAMHlKEaaj1+2GMjojImS17Kr9o/cuOx9miu91QdpPDojVJvlBWz3
ygwm7uw5mP/tzVm17gMorSCnlOzrky7UvnLmkXP4jmZAAGDogsZ723IdDE5q
SCnAAzj3acl+WymDZNrED0QtgKkckhEwY90MZZmDBxIInmFSlYPMHzSJE4qj
bc5h2vRoB8kty/KxGwYbqMUcQzYHyHfJYS4KS/58vXQtURKrMe8jhNI+hHMR
m5C3k3+ND6LR6VlEvlQ7Gcm10HAsEmKuYuLrYmAjrTwIFPSzBtVduxcYAwmL
Dw9tw1YQkspZRkXKXNrS41xmYKTzwDWs+DGJlH2Ckar96XxM2QQpm5OtpCge
/v6hbJA4SnznbAm1TkbFJ9iiWbBqG1PpiFM9ATNDxIIwZvxymZha1gYQALgk
XkyVD+fEk4bVqoclC46wak4cHKtIeZ29bKNIkryyktNo5diT5q2QHf/jorDk
/nURKXnCTACTwV2N+VatLljovmNUqhBEuRcJCVCVsMuCTWYzLpv/6zC9BX9G
wy5pA8t29XUnAhpNu+fQEnC3SWSJsPO6jf5F/lpYJc3KtBItLaoKU0cMVFYY
MFd4yOR2a2LLToESGhLqWJ/mBwtkuK9QChv2pOQcD71kqaeV1eXLu3R9XTxI
5t2OL9qSSJORH5XlGtM6/E3w6CLACLW5fkXZ8ijYLWM/axEZmcSPXEEkhdIX
tWW3gCC47eGtzwBs+zszwghA8R0jN6+czp24n8W/1bHQ75iKSRNBBeo89ETm
NY53Uwav5uPocLqQoMPpZsrTsaA3kSOifpgr3M8u+5EDs14vPXar7lWih3ZI
D89XWlQs7W5bJqillU7SWkB1lS99IBJyeg8gkWe6xpgx4HKcQuAaLVZywWt3
NSkl4k0UO+AmUN3sLDS3zU2iX6stDe/RCL/wAS+upOSRiK/rDh6mtyLY5MlK
84OFNGnH0pqyNMSHo3Uni1OovzO0dBuF5KNe6QKT3VReZfpo30FFVXaqngZb
XU8hzsw62RtS4qA2zgBhxepIMHPys+F6fi6SR1GdJ9rcum0Qhm9Ahc0cxmFZ
sETF4vicQxP0OGbdrQXYAnO6Y8+4htoSfzg6ZcOIYhL+B93x/8QJjjPkt3q6
rwdWcyyQHS5awsJ6XtM6cqXkT7OhpJtgGRjkVK35ZlpRGieXkW+JCgEfeeDY
1iw0EHxS7EGHFD9Wffy6PAb5+OOXb2jgr0Rc0OrmnHLzomXjvNiAql/eOt4x
+uZGKZGF34xoLrCg3BE/tQNwf8uNEqeH8XFWKQ25TfcmlT1xOa70ez403aps
/qY2q3yeHBl0jhQ9YfpHtNS2RbujWNjT8NW4TMd9E7gT1rEhXf9veka98vQA
qS3W/ecOPdN8leooLVHWEO87E9KH+kpKatoqh5UVp6cXoNojBGVHufNcadpA
Kd9l3xaPBD22lnxXBii/huidTmAJigx8y1FUPlZAap9f18jU+cdxllF/wE1z
swYB+d995YjVhDjzHeToaq7ktJUAQBd94iiQMqNVtkHaxxSBhK9A3qz6dUvF
JYvbbQ5iabyCnEypUSgIzmSpT9K5ISVaL4nH6bH/7uah+q1ohPE4Z06RapMB
GljHjJeIAwp3Igiyo4IXH+nLK2APj1hJKeSCaQZDWrK20UiAG4rEPG2fbyEb
UHam64J+iKf/wrKf04UvpLWyKTOR/9Bj9kfvF+om7Iw5LnYoJk4w9U2dPTKn
WaIup0KBDQc2BhSAH0fdJXJC/W1H6jVcO7xwM/wlx1rST7aGkBJracb9QKeb
MlKKXPQ5+0Lqy+lefMlESFRNQqaas2Tyd/F61mTfX0RIb5L6hYrLZP/E8cHq
bbSxDB4/pcp10OH7pUaWTuDM0+2TMRUXI2MNKyct+niDzgf7sJv4wcE5Bztc
pdZHA1cFDLKf6dZAEnRK1KCiWmqi8L5yVy+DM79HhNGIzw/rHxcrUq0QIQ3e
xTzos7er4hgIqH/q+/MClQRteyR/ONjzloe/vO8dQdF8cL9GJcVz01e3RJtK
k6+qBlhttDP+xQVArtxm/RgrIzcTdHH6fvifu/vkE2Qt7NC9tvLeycQ7tik1
9x7LVRAjfwocFnU6+cLlsch1MHzMikynzZFTILsFcA+mycgcxq6dIM0B1v/0
xE2Q8c1q7L3p0EypySUJAhCWf9DF2ZYzvMUoHpya9q9mu9OGtQdSRUF3V423
93sB+KQYaW+Xm8+HzNXHUWDKJMvyFD6RD2h1yQOCmzwHEGwzmSQbwhfLHpNe
RTcLDDww9Q2asZwhyubxKyF+KfZkAdZFqFghCd/OMN0wICHgRB1l4FjQWVRg
5UZEaVaOxqM9m0PTWcUlRijES5LeLJjUFxFBOn8fnojmN473431L24YFmC0I
HZHlwzwvF4BIUDS0nvUXCb3FrihBdheGZQzlYGI9rCNiWTtaulxarudriiQ6
OqFksX4TkOzYhag20puuMYb5+2lgeNd4pGJl//l0km6z3RjqQahvR6COS+0d
0Al7gOESaZOfYmob9p8hCvxJXg/l0qnxWa0g9la0EpIZfLA/rfh8iDQ/ITp5
p2j0mF9c09W/pMtMuJs8nq4nXdqB+6aS2nUbvOq3Wbxz6CO2YlaXB0A19aNO
5Q/aTacQBmrSaK0aPkzGrJSACkuhTTxQWNV3qqEZcrAd1tepegFEHlFXH6Uy
Y727r49GHx2HgVmFva+6r2hwSlVYcTNjTIX6puAoUA4d8BY5FXzNHV0HzNJh
hrlHO1qr7KSrNa0H2bHMw4zQlLodSFTE+JCEwRNq2BoFFeY1i7Z0lerZh/jB
uuQSrkl528pWnpvElVJ+j0Qbefh95jJMAfdXRLFpotSOEfy2jXDsrf9Q/JuL
XC47Gt2EoNYd3nzYDfpWA0WFBq6h2wB/E8DNSZ0xix5EIlSsdk7Tqo1obDdv
a4LwkzP6c5f8SzScC+lQQX31B5SHtS74NGOtWExgz9QtQbumDOASjV4Z8wo1
xJYgP9ugzCA71s9TzMBm19RTdQGne4Kui8fOIT9DVVim1YxRdO1yBxqqsrJb
/vKeFM0LJ0GbajHRQ5usQWP7okNMJFBU3qtKLZqHgN06PQ9+q7PX9A4cl2wz
yXOKPXxUMua4KmINY+GGKMX38dUvb/6w+KHYEaqlrtmXYCHyRfyKD13stFy0
kFtAKGhjuLRoDKimfOIWOre3mXBuO8EMRRal5nah0rF14+3HpPNOOYWwU34W
H/j3DYipJx7ctz1DMi1ergWJ1G6Tm6YWiGEDSKr4GMahjOQVQCmcxqok29jh
SZpycath2+manGvnpvTAh9UONzmfMzdwx3qXpsmCFNPKTtsrXupDW3rvYsMJ
r2sl2Etv/4ILViNV1anSIY0XB0nc72qdL3obAnlekQ8d0m/hFMIUFumirm1o
3qR7aAI+/nAk9i+SmI/Sp0joiqLgEAfS/ZlC/ZEDRzkLAeADRi7A/VI+vedZ
8NQ5CVViVaB8oStJ0IyOY78O4jrhOexOfIqkIpxWiKWMUsbR1V1k3gJNIIip
xfvdYcJAJurppGuKdlbqfiS0ctcSFzFNPwAMWecDBTH/xbC037Kb6jwodNoH
MpQJLC8wJcWXABxh+UWa5EexKcRvxyUms0/UwF1puoOqP30QZ/i4fxN1R9eo
7szIJbKjUwVA3i783Wao9oub+6OOrtwHamU02W6Qo5mWfsbB5oy/hkq1csFI
ovc6IEQe0qEwRRuV2fIexOZfHlrRTYAdfGTrGjmPsn9JMsyGE83vSGj8hOVD
SUPnMKji590/5AFoC1AWLBhyPFIzReBOGZa8yNJp3fbjFakQUOcYYd1dY2XZ
4sE0jLXz6SiZ/g95lteprM0jvVoIUOb4Xd6ymX1Eq86lO8yjVFLp8hL75pfV
ehp9/rCcKNZqttuXbOIcxnl7R0mxawgnLoiYu+7FzlUCPKONWYnCAOdpSsX3
xwAFPZJqKcvTzscL+hlTuVEY5J/JKuStb6hop7c/psjPBn+uP0eIa/h0tQZv
KkPEHB96/2qy7sgUkIpVY08iLsKqnaFvXwu0U3NBmGc9j1o6m/gpdIse2xdG
j5cnhiLVoKrTDK+qsIqN9FekO98EskXfZmlIqHaApnlquusZtcIUGCUX/8tn
NE5m+znjg2+zCUhOnUewIs+ZcKMmwnktEB2foj08cpP3oUOvZgCl2aFoAYk5
C6tPenpYKMFr35032+b4wnHRO/i2+RiJAsEV57HZhz7m6z5O/x7Ivd9otIWm
IcUtEnNzoljxVLJWKhGotobq4cktsvQawMh0d0KbnrC5ZFlk3ZgOWXfCTPiJ
diOjA1a2H+JshK97Ka9OaWi9mbHZCTs38ZyvSoy50vzIH+wA40IX3Mamq6Tn
GG909VBjEAdyGF7ElMh1Lf2g9kTUdLnTsq6bsKIsZgISO48oOT5io6EAqyqi
4PwL3hFoUZWyczzvB32vl6NCAG8e9ybAwKuj2Rj54P+o3Bf1uuBvryDq4wZU
E5Q/gcS5aMYiYRKC/B26olvEQWtmWr3jNfDwu0Ay+K+mqUrNrDPfu/r/pvDH
sjw/Qijb60uqvgR416B7+L39KPGXHN4XF4fy+3oz0ycxZdP3lz3jfIeteWQZ
DEyg8HbDbrfOs1ZfdvsUgv994hCaEANHlaKkvbutOVSphIEV6NJXi2vdaYVa
6ZBXhbhxw3cqiohngrjseNHoZ9ZK8IEilXe4A4RzIto9+jgaXoZMi+W8Eyri
emwb1U45gEdo09Qx9RFabsfMbFRiSYxoqEE7f7XR4f4feCyY8mjdamEDATdp
6zZB6Ww5GR3IAwAPEQiaQMKi33lA8VgdgA/a2uDgpRAzJuWdMTFerT7jUzrb
hzzsU+EQUkH3AusVOQ45Cc6Vr8IYu8eAQiiBqJn+VSZdjzR8f7qxQ5wzDDaD
YaOmWVvhiCKN9IE1G8F/yJNylG9ax2F+Ic6fIZPp/86+YpqseYEtxDF/QOAq
2tb75eVr7KGP12RYlYZ6TvqPamSjQYmDphWpP2QUh+txRp0obX1n+aFsLAeS
0DFvKBws9Vlfadf5pwdUHDEWchEcTkcVs2tHf4VXQdx/00ow0h1cnrLcD/Za
H0o0u+4QL6QoQT5vMalUWgVgS79jXjJji5oNNf4B3XHIMUirDN6IvfV/MMkO
LdnVDNNvZRxAUfpaIq9hYZyFnhpJlg5vhiLJ55gurTfXVgPuacp/h/8Ziq/Q
HEeB6cSnWeATfoHRyedJp5dPlFOS5/XLYkIS4yoP/wNteyari0DB+5DYibox
x9srWp78QxF9Sfiss0KK4dWVI45mxj/Z8QwhZSCy8ZLQ3ca4yCX67gXX30eD
GpnFOHeC26slg/AWMiEkdU8v+2H2IFxGXq2pBeTMFIX4atCnYPgrWC3ycu98
H6P4wsoizA3sXa3oUxQOQI8pfmGsXpWYX0AlHgCDTLRLvMsHyc2vh6/KAcYE
Y2D0evFis9YkraC7DIdar2SntVevlwpeOZPuAxtJTl/4tTT+slH6fvImFzvy
NxucvKkPW/d8ZmiQwCQ688ylSNqq2VTB+PhzKYGhwh59RIfgU2TSGjK6i4xx
0z3uujSRleb19zNEnRQTVYi4LOzrpYkivFLwJJ32E8YNEyMuT5YMC60n/0uU
RKptlRswhTumbnIetOxHiwpUF+c4078k83wFWNlt6Us5quh8w7ODAC7gbZjU
wT/V43BzqKfwivC2JBNyYhOxXc7BjBfFTS/NmoSF4IqRKNwRz51cgs+MnxaI
kKEfCW4MiBlBG3+3VWtkD5uh8BGZvxOSKwwTDzOPJKOzlGhFEC2SlKSa+ez9
bfwBAbMwjsj6f04kuXu1J3O7ni0JDiHEfNlHI0jeDSdTvScgGlWkO2Vjvyn/
EJP3F1sJ4kncbF4QBQjIl7g0ddlnBJLyqmy8HN0gtDDwVIaJtEH26DGTfwOC
fIWphv0T5C1AuOXcTcyjsLMxGCdNcgbKwg97zqHR0aRtOc2JYwI/HlI74UkW
BEldZkkwmBjdeKBbvVK4uwruq1/nU0wZYrmYtbGgDd5TSiRmsJJE16jKNjZC
yGKhKBbUbmuTVxB2JbvswOreAKJHnldqQ7RCkOyK4P4X0d992y4D4zm4uljo
sEWJvrSrST0wnS6jIkhNhs5tfKDsWU+dnRcuUeO90C1icg5DdRil/Scx8qVd
wYTFnP3iXF6bhXNjHZfV1qJcZ5yIPK2+OLjdEW7gXWYYQaHzGcS4mlJrQVGk
Z4OT6DgfKC+4IUmF7WVS1YV/4XAjSEYR8p2T3MBktacniDDLm8o1gg6IGVDp
ZFXn2vEwzk93AvPDatL1uDOzVH20FWJRzJq7hTbuQD3dDjLr41Rsmh7xsq8p
l6Q9+oHcY+jCDEuw46huWZWV/2AhEyo3WvkDtQKkwG4LzIszcy7S4Lq+XwfL
vnextYsf4fEqsewNU5fPKa9MlajcC1cQyJx9Oar937UKcDBLbZ30pWpDiJNc
wOyb+tczWoILbqM7//sUbthfU+3+In7/W4RiEHW5l+2qQI4Efu64BSzfoSps
DfY6/FMfKGIMt0CFOHFOqb9c4O7E59K/bGUpV2+7I6Wsbo0ogql5Q+ey/Bxr
gD0Gp4Tqg0/PA582/Zta7x5KqoyUX3MEXSFRxiIXw62eH1Jb98ykjquQDwH2
0TZBts3+9/EM8qa+xxFCwtNnTc7vcAcIGSI3rVr85BATtTuwL8UPyzeOB88S
jGbD+iMUN7QsEl8HHofH1ibZFbcZcISrYVS81qba6t02FQmKtwigkuv2tonx
CGR45N7XcPPfwpYZMjZ728q93r3AK5FoPc9/fXWKrO9/Buz7o9mCzd7MtjkE
VngJ033/+OTk96fhY/ZZO85goIJwzO/Q9TcRDqncHzo5CIZVzUzaGNCb598f
KFXkHzpu3GIkqZCBJXKm8xeroHLQmHdCcHRi6nUF7vdszB8741TxuoWyJykA
WBXxkFbH3WPCLCZl0v3Q01NDDiAvQT9JuYWeSgJEqDt/AtLKCH0SCzb/nYi5
aQFSbKglWwBmJ3Uc9vuj5pfZnhdiYRbD2dKiMK93ct+aDIJcWQPzK+bQtQ6i
obUlWH1FlaFCVakYXiE2N5iBlXTvcZ9cYHJQrAVlBRmpBD9ZHFNe9DlpY1NO
6qZOOAMV92OV3S0AQSDWX2QYYjyBSMEBjVXzuMeERZMWqmIs6FWFeSk5gY1b
SpYY8xCGIHroz2vDItSUa/oPqGFLSThMTtaaINqysdVXyt1ug0V7zdFDj/zd
I0/ocqrJmmwZFpFAQqcfURVR+FOjm9e8A5HWN8Wjhz0AIci78BR+MTMda90d
zQ7JOjiO6yZ1Ynpg4PvGS/khL2Mlf8RljaQLSWVvhvZB3qnMCSVpKZZBZSH3
EndiPZHoNSVzvbc34Og7HJfcOGnb7iMnhQjCYuAUiZXTj1HSnEqDtiqfdJvk
Fc0dEKJgbvLHNlzXj2NGsnTDYzZtg/aJLz39Ql3O60Ew5pzQph5nUQgNUmSr
6ame0NLz+GZEwJZTxvg/8ciwcBr/arI2fHNvvHf7sEVQZOO7GP29cqeLQ5fV
+Rplp17NnNcfDoUKZ58Y8FVgI2iMcMFX9VZrugc1JLtkgDD6y4SR/r9u8gSj
60+vcszkY+7Ovpiq5NzAtku7pmB9D9bADAx44AlX1nHsbUv0ZZCOKwkIiV7K
Z0sLayUpS+xJOrabAfnZiJSuotfb3N/f+xcREAv+V1NirLP4DLTgOB+6UVNS
px0H5AEQhPpZCJbZi7DslRRUsoYYIjEJZbay04upd7D4AToaK9N9rc2e01bp
TT/r9Ezdxw98v+tV2cXaazjOkmREgAmuq50LPyPY5w2JHk8SJcJyd5CO1TWX
DxL6LqDz6+Dp1Gn3gFCX04WLEpBW7gHSIuV+B+oKCwtTUcD7w2eiK5wk6hN3
i/Mlx5BJbdaPtQYY9E6Eh5dqPKIkCA6mXg8iBJ9xYIp/KLjKAa2yBy33WAuF
8S/LQJBJoUbOosJUttD07anUmKKEXQicmtrPFvtCsZU7z0baO8kvoWMricLi
LFn36qf6xtDU8IB095kcRak2JIwIIaJZarx9IGm+y/7fZA8fx1ZWoUWAwTgl
LgETbl17lu6n5iOiYQguQX0jYzh8mjV08bRtpO6WPbEvc+MuZvuAVn8sofk3
gEvaA+IOg5cBB1PfJf+ntnn4HwtlMkwf3JgfjimE4Bj/eLElqy0J7fO82VY/
3CSWnOCwprawqPKpSv9hB085+Ao5WMSl6zfJeK5CMNDw6doTwnRbybT435ix
hzoTjhwLnrdkCdbA3u/FX9s1NTeAlZKgUmr4y3jB3TY2WWiF9Phj8OCLTWNH
87L+tszbCPRlevoGgZ8NyxVfMJhZgj5C7IoSNSw3OObvUmx9dTukt1y8C36U
u4k5imma/6jUtELhCzAUUxHgyhKWF+IOzlkCnjHpPjIKIwlLc231gARNoXNy
doOWfT2pg1+A/I2SDljPQY0UY7wDAIUIlKThPXM5UYHAmQllFHXUMKTFyoz8
a1Ib+hXPm8gjgnOwgB9SChNLH/nTQiu3MyFEfA6EJ0/W0zvXTvOcrx0oNTKu
lJx+yJIsdcv4FpJHROb8+iiYwLgHs8/oztf4GQqGTBKS+jTnEfm1BYPvP1Dq
Y7QMfzJA+bVaFPwq0ElRMfRjdI+M14mPvU01kKBcp4NdIR/PFLoplpVIF7pU
tnEfvJ4qsaummGODSi8q//QXSkBQvB9J09abceLgmfKttCb62eHV0Owm3UKF
ilacZUWZ/My1mh1bCtEsJAuXM51TrnyMCeRdCvVN2x1JX62nOJgdpywPuRPq
FgvVCdun1urAsR5yQxoisKl0i36Afc3AQJqifu7xti/Es+NrcJtGfWxF9ZNB
0BKqFAqLIuTGhLcSOlaswnfsHnlN0iozx6ShyZZ/WPE6sSK2enRcEx7YlAUB
geTt5EP4sB1rh7fRpGcYQ3nfbNVdI0H6WjiT8gv8icVqxyJIT0fVkT9ujdb5
KdZLudSlKrTHnrGm66vw5viX1FV/dkUiagFi8cqN3TiLUiWmG59QrBh0SCmu
LODDrSBk2bHkZxR1nGgb1NSOykkvqERjFLrpgw6wbhhFKEU4Y9ZvNCID2XKl
6mq/EBdfkkbR/B+xPHkvB/QRKfD3pOeKL07w8a2pVhYblLpq/DmFimpKifFL
zB2lIhoRkoWpkxmLMIJQkBJI4xs108hjaaKAdDV0NGXmQfxjkxYrkbcvvtlw
ckGAMvGJR1JwES8107pHJ2SXoIjs2QwZoE5c7R4SP6kJR6YwIX1ztOFb2dEh
kiFRGmRl8fgag9LmAqIPuiiyAbWJoHtrWXOnRT+jIbFeon05ZUb318SFrJ/5
JgY+n7m3JJ/w8NJaC5y5Sdnpny3Dn6G14bVJ6DrFBdQcSpFeit57/csrm8NB
/s0bFTAD1VqIhD/D4mzhFgfvQexWF6VUjMnYgjI/2vjpquz7Km+Pf3vpcu81
AwCcZ7la1SyUN1wUbDM8n55yi6NH7zrc1+GBltxM+GmP4n/P9lGu96XnscZe
LJoey82MCvIhqyyvHjX5lpLRC4w0y2ua50KfMifqCofwJtVJqrqZwDbU3Zgu
IaTBU003K1/9/nrBvShmakAz5R4FII1BsVE+61lgUoj0aPrVFGgfqbNil0my
EL59BsDM4CcPeydSITZNWsNtscoipr5H1xkKqemlzCLtKLcyt7hEurAKFYhd
1gqG4moP4DBho89MZU7FvRAnnN++I9W3cKTlMA/+wu2SOCzAaupWJgUS9wiE
xyJZugbFm1tBFYH9iV8TQBIaBk4Aivjr77wTzfvNqhSpCP4T7/ovrhv6G1TZ
w4W7yED6QUPLqf2GR2jsTfPrjzu6OCOQXwn0aZjTz2mnAPwlexw58xUpOmLn
Zla6s3odfhdXlBJwtls+SVmgvHajQnHDD+rTk5QqKLdAZwChB/25xGkCjXUk
CarMGAk6CquQnh/dDzptqDJn5vY1ZElZXccKdGRZCLVMrhMynKcSByQ/jsiJ
UwLAV56dDHwkcdxy0SKLtfxzzXpXFjQVCt8ZHrMq8zD0yJMmbnq+Ydmzrtvk
oNuifGYXjtwVC7XzdDxwLHDe006NrN9s1NXQqUunobK5jPcVuJJiL43HyU04
jZ/0tMP8YRYqsqnfaSLnyXrMPWEh7Yhi0BwfMMe36wFsgGed1HB8hEBYD0Fy
sLoI8+S7yN00CnxLq+V6lB+NvzNblLAAx7jiwYRppvXOsDbC4A+EaLC4un5d
DPeDqnP0XNxGLzhpp9T+K7b6JhiBOMOUnE+pKyfcyp3H6HWBFU8GOnANgJyZ
BaTBYK+Ru7fWQlb1vXPbFXkvTG7MP6KL/CMfCmCKe6KLt+vdHnV+N9ur8mSV
Juv3rPJCc7GIOb0IJ/zwI4brKNJ10X8vi2bSOMQgbbuiwt3ijMb/LzL3zB5+
5rmJv4+aE0nckjaPpppHapqgUxRg/qZSaELCa8fMDRjPj5VCYelm9glLFStg
AJwXtVHEZfxd+TNZNJUnTzNb7WGiXeT8mbf73b15pWL89sKHkIxy5ufX8mEV
C+zxmoALM6KOZzWqOUTbsVPDBSa7IJmiVbunJL5YB7CZoVBAFqi2npXL4K40
/gn3ttpE3yI6NrnGwa3mmnmHb6k71MG3GFOB6SgXl6l3/LQlrEWwrfP6KGH2
ghxzCYgFWVVtDtaftno8wbU/9IknojwOB5V7OHvVlQBizKvTT4bpxpD/BvTl
+VfS/HdWGLwxXXeOV1eTy6xQrC0NSvecuyi6BY8tE8B4uxzy1DSjtzWcCSZL
1UM3ChNb+tsznm+WQeS4LqdMxFB5E6Q+XUVxNNjQESQVug5qmZGD0DVQJJHZ
tlWqKE5AFL5DVI3woqTFtD23QqVXtHfqYdLTOH2f6mp03gIG7gzWe8GLEqLh
NNjMWmuoFSq/+Izp3RC1s5aAvRHtB9Oy7bmrumHKy38NjDmMfNs3oYVg02t9
UDhdFXnbDCQeKFUTX/jQxC1nE+KtVHuskP5cHtsx27ZhUcCpfjqesaTWcuao
mRin//tmaUhIvJPX5Z2m1hQn6qLOlVrdPYoqly7pCG4hnJcV4Rs6OrOmuv+X
YgTg9C1OBTxwa/QvrRPsPii1w5HEisB1UqxT7e1CWF6kPKE6/qFbRyWVFJj1
eyCSiOSJxEI9JHQ1Fnt3cdDc8lyog35wWB2dBeU+IGsGzVJp/MMf+nFJQqbF
i3Cr12w3l+U9R0JozfQWTHM/C4BFXmA/6YNEEt2bUYWyYtmglj/H17nKeOnv
9f9/ITF/kskHV0ehLEPoR5GqBxNRzvM1dN5TXAyJA7AIqdp5mrQ+uDZozAqR
miK8uU4Wc0lFYjTPs9+veQqPVmpq/SI1UwZ2iMp0ES8n90l+34xzvlgSJnlD
WE+XYJ33gsIA8OPbpkM4xxGC0jM2/1umNqelDDFhNk5RvIPuN5uu8mEG+bg9
XA3PMd+ccZUy8uWQ8OUZJjZagDbGYpiBo1T/0bsu0/jDGc0HBSVaJZNz5VOr
9615oGgMM5YAIhF7TRIWGZdNLXGTb3aw7dhCFntcwkOwuitdE+ueG4HJWfk+
9lJk27e2nEffm7r2bud3aZ0rFl7a9JHDz2otVL+fkofktTjtQh9GwQwbVAQ6
RzgmH5vPlZJQHT8RNyQdn6sR+F3F1SgtJIAlWythaTw12wL3J7cAZJjNqGwa
eiPGGPQt6aCvzl/XGAu9ZwPucZwjdFxu51KhEQ0jW/VReCK6/s5ADDKc3NIo
6A6ije9dVIBy6UWTJWwoDB35gOMtBglZXo877v3gRVZe4RClBdK9erWN4Y5h
F/1QXQkeZw0GnVgPGijKo/aMYg5bnDd0I8mbvKGJ4wnvTG/jOR8lu+tI+dn3
2+iPDDMAxcPT9ULZP/ljBT3nX+xQ7+bzwBtafcmlne8ZUIQk0QfyNC8sn6Ke
rnJk2GihpjKd/gIP1KUCUc4B10oN42ftdxhMZ4IJ+oXqh2bbcHOxj3LFA+D2
COPJjSKGw9KmyNiWu+la/TF/vUZ1H98HzfCq5GYZJZkgfaCl4g65zLt6X7XS
wEtkXW0wFKpu9em4qjoMakFVHvvN/kK+ROI0Q2XT69oOkAGrjEBU81xPpdc8
QTjtB6RMPcGuRYBDYyBMZZJJXB9mQpY3Yb29TX90c6YJYeHVMj0p8Dv6scHD
QnsJv7G5qlBHLsMZU0KtcbUx+VeXxsNw/339P7fDl83biscx79kvV5tZ/1Jy
n6EzOKBrY+kL1UrbGuJmt4gt/CeBmxa6bNzbRDwJmAadC+6X5ehRy5MCXBOK
jsjBE3iLksmfqJTnqaE2qyHRFkqwMZBZc/MK9nApASIHIIW25E0AfhmjAXsY
GFrauiDSn3aPG9cFF4wUR7LzCG+1a/v00AS+uHlscROcyjMwhjcBKFQ6vaYz
V3uMkl1BXmry+N17rE2NsIumhdBzqML2L453PDBThOQL7GzT/vfdrabLkA2u
zfKEhDpssS+PCfBfhLI+pAI5jTGl3+pAYaC3kJKYmrfIZeHd78m5RVItFY20
dxtXZRIZ4sK4wgbBboUYt3irhmjm4NaChsFTlE0fWtAJsBw5QbOiaMWg4NQe
1ekrESqRBuG5XmC7Fw9PeYAL/PB8M1onEd0mNK1E6dietu40N6fvxurNB6m+
s/iSh8XebpUQ9Mq5Wdt1OvtP0VZHgTis8rQU2eKe1GyQf0WRTpgBNQOUBh0O
OqbznTTihHMPFH+sbJfiKTUklq9djf92B/IPi5W1/yPrJ1q5I3MtMZGk2ujm
xVNfXwFCXPqadwxYifwR5QiP+KQ7NnvO0KvYNGI2fdkf2Xh5WXXbcwkTvpd4
68GtNu1EE39PHldtdpfNzbIP24PtCWEX0CFiVP6wE9OgYaWf9KEasVuZJlQs
2+tAWdnUGYwRJT3au5rwydmzU1Jx3dS3u4ZbtNrfVTc3fM7KQYM10ZjanU/B
gMs2pymb/t4CWaJ7izFMW32PRST8gUrJRRBvuPMC6wDjhbQFphvzqKmoRy+m
RhzacnVFeo5PO0rhLeqpX7QD6re6GCDzNqHUA5bcSqtnnNRLNqGIWgoh5KGJ
4mfuBYOwIM36SdEF0cvndNQT6QlSQEEUWQTboh/dpIhDoa+/x+e4sVFGtTwt
NYY1TlxHxuYwMtkr0M1VC3B5xeeMkUqkT/V1jucmcPGOnNqE6M1LO+J+d4yh
khpigoHyZxbzE6ugbLixWm9vfSn6i9gXsOY2pxmSpRmcmJK0KHNEgROpceYX
APdjn4U1UCrJ8uvyTdX+PhNQk+zM0c8Xa28IZs6O5hnq360Qj6UM1kyoUr9R
ZZJN2X74boopVx44Y6jlaRmpPkjCOEo7kmeLFisHhznYuDc3GK9LVxAoj01t
axYo6UlncfKA+FxRs22922/DEiuGd+EQrVtkzNTHXZds332RfdrsoYoqfsNG
mlRvUnBPj4y3NFCShdF06ri6g3H5xddxOMvl1JuBeLFS556rwM5wF8dzHHIh
NJBDtnW/lm2oLZ46wcyGuxi7zjAnLW6xJAAj+Ji3szXrtybLQQ3XwqQfjLhj
rPbZGkoixsiHuUQvEoa0tmyKHDm0YbEhIj/rkiGPlntku+Ws3bqGYaUAfvHi
xmS/qISeYLL4lt7lOBfvfTmHvsV+hqw8kKSJB1ogIyqnYBMFfEQTRsyTetzt
1Z3SJHW3G+5zNCoiYpMIrxsQHsiqrl2dSd4hAyQ8kDhJ1LHqa08YwUWe4tnv
ktKb5PEyi2A3OXT4ves5l4946L6EULUvn7/lB0rE5ILKRUy4WqUvZ1SMRtAy
3L0FRP2Xj1QG/mTamX7GkcwrK3zOKnUmtP2sjbmEPL5T2HcpKNEa7ISQWq2P
woMzQlmmVnUCVy2e88pWvjv4j6RXTj57hiCV6FdvDwESJxuU0YwUUyoTKLMs
JrFkS1JMySyWLV+SvtZDlcH1yxGF3VgQXFYm/T5mIrsSWbBQbpT1Z9682OCM
8zQUQCL1URWANqDDwKmHlUrZNdi1pxhVQIlyiaBt9qJrfoXa8rBVooxXdQTz
9rcSGNxqZDDZEPRjhyWrkjCNY+WT4aD9znpXNN4jwLt8EgU81CUIz1aTCWwY
eTYLcAfPM4OF2EImH4GTP34o9eYDDM6ovjOmJ9rjaDxl+6G/25zcpSVyHums
kVr1sMlA1DOfJPn1R43b4UABlmwwZZfTtNszYIcD7mBhQJgC6dyV6hh0LmnP
uREE3dOe3p9wUrwnmQDPnTqgOcGzkH5MAvrS3C4Qtvgglj7Txm2rXmX+asXZ
gD94wBR1tOqtqcqqY0+gromlZjPZ2BhCuH47o2gFXXWI5fAXCYeq1fOLVNnC
7VW5MdX12LU/eRXadM8qcj61GWCYhe1sBX6Cpc/HqyRWIPn830d/56XOv+E0
KIQFALnmtYDZ7DrU/jDTufDfSNpk09wH8T6DhmpdNwZ0PaLek1LKN9oRzrf0
7qfqWwLs/1Eom8EzaolBVbcv+J0lfe0Je1tZ8skEv/LTE0Ujgf2h4yIF3QM0
9z3E9hlsCLwBhzwU8MkKLIle2T1iyNwEjtqNkj5jN9saC5ti91pYAncC/kA5
WNYyFDSKwHggcQifSs5rYaKiM0skW7ujPWthd9TExe72qpqmDZGkc9o+k3dM
MJob53rUWLf0a0OJHmZink6NHCXYpERhcwfkPkyK2xOB2mpTVu0UWFL8vDU7
ib3QsqDDtSiDaGVGaiSDkWD9iM0Rn5yND4YTWx5aAXGZv+FAYh9cwbIx6hUP
Gqe6CKd8RRpI8rPyEhwmTvjbWWOgdoXsw+Hae64QSFkBeyAjdl12aGhshT1D
KzNkk09GXRl/DQhWGHaCFUNM2qfSwH5vm8QjZ79Aeoy+2DvfU7LRA7kWUzW8
SsWx9kt6FWlatcLJPHZjfi3Pce9LNIfr18Escnw//tGsEXKVexQ+XEssR6dq
8EkIbIBmjvVOuO9LnPiXF1JYUzdvGyX3TdhLxoX/cJk+mmUEQ+twmnY2kXk1
w6N4hAom1HvB36fqeRFLutnQoqgpqjl+065GN9uLGLKY4Hd21+xFAz0XGsmG
CdvStYuIJXDKx/10XXJMBe/rkj7eBokS6VT5CvFTEbydcgkJnwpIPrWpwKHQ
m3M+tTrJMQBiGDSeJkrHOM5pNGyuJyWF7agRufKslFj9/nQ2S9d/+MzJYfTy
7QfBhrRLy3f9e98QSLgvCZjrsGoz1wqJLMftS2fW5HlFO935JDDXh+v7DADg
/ApPg3CB9GXpGHAYqdyntvC2ZJIvEZ6U9tQB7+v8NC8R2VMNgi6HKijh1KPa
8nRXADFRrV44udYCJWA3VDXaiivTrHnZeSQH93k/WZuxM2VLB67K0qGxSW1Q
u230mr2tNzssAPwe9sHE900UL6k1B6TnrMr7n4V51dMz0zI6cg44yXrVseL5
Xtnlmtuq6yAE1H1S0IFT20PKQsIh4hlYsofWGAjOiDZRxx81yTTxhCrTJTKn
ZISGWiVFyAWWzSBzbrY/UWCkR3j5FipAV0jdtm0L4cjcRONZvW8v20aFIGUC
SsVQ/aLNuXixaIiZmIm2Y8/tLTZCa7hh5rj1vNEeknXCV/AOlYN8HbJnkIkE
SAIX5Zy1tvkxQ1KlcsiOzki6hdH/1XLJ190Q7EIYJupPztrPN9fUDqlSmpGG
DpCi/J3VA6/UNAx86X1NYCU++cIikALzlaU7t+R1U/UWsgm64aEan7pv9o+E
hzQby7CVO7TtdF6hMXwO/eYXmlQB9cSCzBOnjhEvrUAIyH0WJTvmBXdkVMpd
0eqf0QIfAzAMXrt1TAaI3ar0M72OoBHhSdT4AWZ/yBd1hfGJAmdupaCo2xIy
LMnc7QkW6fkKK6wocuOUlmUfbuFk/LpUafCz/oO1udJPAH6lxt56EyLiLH6B
GCZU5K/6hhODNWdp5iEAAHEEiUUn2eH7cmDOndIaYRPmEo6KXJ9twK7ky8/T
ESTaiBvGkJfyxjweRrcHxh1L89EAfmXZJyz3fZCHMe8Pu7DMBiWs9M+vj77T
t7wGuS1XHNGV+6BLJrgWmDrx0VNQoNmLEWXtCvBycZ4r5SGC0kwwXAj5bb+T
fFby0Go9/azCcUvTBWHnRvx8baGC0MjK+J7/kQ2Bzs7RuChptSs8eQgNLBte
f3qFJfbB2Eqjx0noUC3zPTce8n58CIR+OqNO4AKxfqdjB6+h6n3gTNiG3D7C
9sc5U14QBAAK522rvzXBo+6sVWVaDIkyW6lw4JfndQRxWcwl5yvMDo9Xlb6f
mC1xE0OP2i/tfTtlMdhokBL2gkO0vs2E0ZKq2WdtOe2nFJ6xCVPcJzvC0MeT
gtSepfpmeueWhnDHtT90DYUJ44c7KWLWwNUB6HXuASnlbXKXQXeg0B9rn/Va
UudvpGdb+6ObtpsfdUy2+T/etzpDIYsR6nCMvT16i3SdeVDb+o8FzMTVd1B9
98zmnVkxznfarjNEMVp+qZMttoAN7CN3w/RSm/RaK+5IrEnBHgIBADfLrvcm
CsDO8YBWFCNJCsPZAJmriOYvyyrXB2S4hdzZRfIBgUvROTnfGKoAUZTV4e9V
tThy2sK1tLrrIFyvRXkH9LRyILzkoLuuZDWVCg0IEDa2I9L/0qsR6ymiRNyj
t35FOrwSypqHb7eiKPvRlIQbHlvF3846NERJo5O4YAGLPjNLW1rNyPbtToEJ
MjiTsvbb0ijQRjaFbVNY7vgGeGr2WwKAWWwNaoNSyzqeeRrBzaSVwpK7sNGD
4s8RaJzWRXk+q58Oq75+SkKjLJY7usB+uZNWLQjILEdC+txYPko/JtTf+Suk
wtnHxeKrXTBOrMtVHulhmrEnc/vZy2CiGW1ctk7sLPPpALe6ileZgAvlkvEG
bnibaV3xzu/TTvgyPOt5+oQxNmNGjDY0v3l3rQ61SRE8cWp89zrjsyXX1iwW
Fy7mPEKtLpmpUWTUPLzLto62YiX6T9UE9kqNDSx/4XpiRHis/RvewZ9YX72Y
r+jrQBXVjAoG2xH7VoL3KR3cmMGu/KXPx6uLuo993fLYPRvCa/SKtTQV7pwc
VMDimuEfC/p+ePepoBV5vgHj5DY14BWOZkqHnN9Z/DHF/uY/dNskQ/lgQoY5
Iquzp029WqKzA0PAl9sQZBvPxaofPcWiOzFeo4cpVoF5yVlTzfapYnIPkWEe
4pa75u+2yfuUXO2oB4AfwigT7iJO0n+0PkmpbFiETiePwfQZQKHQ760UtDh9
GyiXL9fbPls/GE7/z0IcIc/t6vZJdUFSWE4b3Pn9PzCNKRIIsfQU/sLy5qJm
EC2wYx2YXxrhpn0LfLRZjcmqGgBuwQg/xkUQKPTjmGSHvIlJZXmT1Y6DPGhF
2IvDIsdeN4vZl6aSdUCUT/dmfQFMlBws90/PtsHJEK+9DuKv/6P4BQtzNUFg
8nUvoYputhOCb99aUN+TPfHH8QDHMajbrhXrlGjbOfkqUSD875IJjNARXfEW
ALoz5KNIkWEXan3ZFS4qkVBVoOiJ7Sexq17xzye8FMHoekwCxor2eh4u3D2M
CFO9vvFUl3eLFSwks1QknEpvNp15mS9zwF6sUM+uWeNd5jY7GMrl3YEO7Xdo
a812OHpVAb1SSRAHOcLXg8/uNaj8pERwdzjOYwARWDHcQn3Z7FPlVFMc7vpf
OaMSl8wIcX5v922F4o0nTvykWdoKyucTv5Ms3QWlECsgdWS1fDBH3dgXNpES
Vbzd+Y172UhWf/M1Twv/bp4/mslL8459GsfJG8N6ClqQK1Ur2y851qvhLZOB
btZKW1pqYS9Pamkyh4Uo7dPvE/TYm/Ud079+xoVK60X5lyP6Ykh/fqKR89Kg
izxoTcBfSXOWoCGHMHOSnFwB62sVmLaIVpnrrcTI96QiHXQ8qSl4ixE3FWyT
QgpWqYBCVtiNSYWCr9ZctL68rNXK/zJEc3i+OprSKQm34JpT6iwxlVqJHQns
JRGv3SKkmE/rthzJYa29n53vkrmmQ/kTqGUn90cR+9Y5Vw/2tj13qpKxnLeF
9K3n9PheE/tgiHVM1OFPsmdI9PA+mugk9LWJqISjfe5jh9NYbbMQ/7xN6tLB
wTrSTa1G8fYj19NTjDFnhYnkri9ZxMOxq3DnANxvUOmRcTODnzqUWsa+GQJY
iNEnQ+tZsWvNA9Kdk0x1lTW6Xxrt7n/lxhCp34qq/2Us9XKfykLtq2wK0+aw
SX/EL6hlCd46qTzuMM4Im+yjvHxliwfiYsEkEkX6NROZ2u9vv6R+VjJ0h9Bu
uB3+mQt0zoAxbcG+2JT1NqGzrQteOqBxpfEmLaPnbtgUEO123hRnAw0NoM9L
tB973yQArI4BEISAAQ7qEVEvXJ5ZvXwkRTWgPen57z3Qf7FLD5TzMNPe8XjO
v89Ttv5w6HnKBO/+GHSoGlMz5ezknZJccvzTan8dK5GKUIoNRLZsLX0vHu3e
3Vq7VUWY71H0weVh1yXtyVPJ/fgLRdMkEzWo5IA+G4HXUa7sAxwu2nRgpmG/
oCFeAFXZi9po+c3b2bxw7ZMqKaUKvJo4UpRGB2cN3iJOcgWqkTpFM+1zFK66
Lp/LfaBEC0c20WZKLSuaPnqFlLCb89XdNaQUq2XZSCFnKKammDr5/S8QfnpJ
Ajr7oPUSKMJRSehSGZM7Bi/EpytPRl2Cs5wmEoeOlxCFg1CmR2CBeHKDT2zA
2EIaZgITLNFP0gm2sqwcJSP5jdLvi2xr7HgbKJpkfElGagr3BxtHjg1vZNnG
BKOUCujquZjun9Z+4tV2QbCjaFStJRQPC7pn9sOkDJspakawsj49xcD6jAId
VamwCatkwDLbObZ5g+3ApK7qhxMemryc8xjqOBY1vu3HoHu4LN783fryqmfq
++6G3txpZR0G2ZjL61jnWoCCVE4fb4HSZe8xAN0kBhV6dAEWPpuZfnvgbXF1
ag9Wf6Qk69A99lyvgK1MoGaqvfRjPWpq2m2YInLNedgUqFm/RtCFAcUHLruB
0HxPtiX9j1dEJmvAQ2H9bKZw9nqkfhRMUtQAm4zSRvyVBsAIGg6RW3mjtXSR
PPDXjutRj6gqhYSYkvitJypI+2f88sFRqU2sVLhhMnbU8sCzNH4bx4RutdRZ
IT2y/8NIRDBx+GWsecBz1TbRoT4Rgq9BrT/TdTO0O/T9ZTxxk03eVswN2kMl
Iw4qrNAkYerjxJbqt/+/+emxt2oeCU+v9A7Lauj7IOkG/3sE1HGCUlMPg1rw
eGTZIIV6sP6v2rU0XuLhiGczJ+pDiCeDo0SFvyJyhZzox7BDtGBU+ulW/TWl
QsUeUTnaOBcNv+gs/BotMhkOiWE32Lw6aOJBAuxMx1SWv2N8aECfQhCbLlxr
bqYq8efYYatzb/pMH7ttU0VG2C/zgrUbJKgCLi49xsLsOOaf218ZlixhPTAv
iXz9P8SEq3WoJbemdEQ5KOP2KsXmh3EW9E6nbaQ5IXsf+R1uQbmo1K1kc92b
JWquv8H5NZpladneryn92gjNplA9rwPXP6dSjTojp+3trZ23cDwoWgwB6mSi
TFmn7Yhr1dbmc9QaQNpIAdRdmISe6vv1NB4HiD3hn9YHL9cNMarKs3a5oqY7
4l1umMglm2H78CbSHRGyGU/vtJb4N5zD0+q7fm6+5OX3qUjmif0WugbOiWzV
FeMf9lRvlVPS8u2/uiwoO5dsEc6tn/87tU7G9ak11igMPVP4nkiASsv3wjE9
+8hvzMfjH0jqKkf3GRuyxqey7xvFVaBTCZwDPN4LOYwa7ZpO3arTREcC8Xdy
R8u5fgkFc9/Vk9eWdaYVRNtnn4vCkVCHHv9xpdeaq8W9TLBp/MIkkop2zDp8
GaIOTGQbKWdNdQbg3TrmJKwXIvEpWelb4sGJWhAK1psRp0PZ+DxQJXpkDsHl
tWlv5znegS2t8yX6iEE783yLPSN1vvy6jpYxZhw2c5vZNE1rhos6csOSuMm9
8n4weorA+YN5/XnKxd8T+TEsRF8ch88qYro5fEYE8RKZ0Xxw+4uLGneveU13
nedGqwWzBDKA/79+UtoFHajoRqKKpfwveXkIh5QQKjBnpDxYA0SoQvOaoByy
e2PkTCYZGDJpkZYkc38l1/jCITeN1+5J/D9gQwuFcJe9xAWU3YEWo2WHlMSp
EJtut+jVCUpFLLHfK1bhJdO8p0k9RK6JFyzYN3D7HO7OOaMs5JUjsKOxFzQU
MuWnH/AaT7323w3JztiMFn4y2P4WABzLE9wU4Bf97Txm2etp1WeI7YY+8qvH
Gqza0NxEgW/yq47yS0j5nSaTtWxkKUkCgv4Jclxrzhi776wM7xzZSIXUD/Y1
fVSZ11UCFxu5pqN3502qKiMKIujIVq5QmfkTdotz8uKjQWBdQ0LKLMj0QIl1
hGEYFZHWmPX69cvCV4rH0NkquEf15v/FsVBcA//jEIhv6KZ3ijlomMTSLpn8
iYtQS4zcy+MTBiV71gjL0JjPFSuKU8f3GmCAK9D64NxiUOrrF9mTg5UO/xwK
cYQ3gc/TCN1tKfk7Wbs3BcwJZLImRKV6e4jiAw/1ohf2iOH7TSQ1IGZQwqih
wTVeyjqrbT+20no+cuw672ymOrK0vFNwKU8TQqQFRXXl0u9oeYpT0InVXLZn
PdAt8Uh1/4yh3fJpYtu/6AN47waQfmFGpe+/CjalEFQP/6YHYuYbpnzI+suQ
7ZZUK5bjkZvghcYFWUuxcfmbGnOtIDz7hokm2N/RV8C5MvY+joL/35dWvBh8
CuD+ulDhpM8NYt9dK+OI0kEQXrchPamcs8wC30ssP+YknKo9JQ7CkKERQtp3
JVAeY5KGJgENnkP8BwnN6b3KoZQrOQSI4sQoilKsdMpsYP35jnyxqwDRsR7M
T8s10J6sBeiEkOOGyGlRy15yPGm6mPLb5ztya+wBXoGzgVVxC6Oeo8/4NNkd
yb4JWCiGV0y31ToO5oZ0TTiOHoP91D0dlKEToiWWy50HEap2DYOm5bHv+YXn
w9SG8UsWGNjarmw++QRt6zFsy47Kz7+BsCPTr1Q1vkPPL4kErPIeOUyK3wO/
DpigDejo8SzL0foPdXEJtqc/5U6P5wfCCCfzzhU7wsDwFoMEXto8molkpuXE
lqJltdzQ5zAVlTT9Q9kaIX6/lmMktymS7UrkGw1n3CYf4lhujpVQ/RvURlXr
aIeCAueVx/VfUD9vqxRauejp6DWqdAxdYZQOXLUQxrm0gW7y14vi02j2aoKE
mcV9anoluIpg9c97Zr5bym9j09zEG09b9jMoHLMzQQYumc4J+AAZnYE6maiS
M3jkLVJSXhVo6/ywFQU16v/rVFG1zoJ5EpkvkOZb4LaBqAiJcQzke5wEyqxI
Zf9dh0hyCgkyaC7303+Ld9lNp8HwYaMFy4OYmhHleKquKhjLN6pr0M/MVIc/
IzIYi+nY8CJVGopxHC4XPn7ZE6uY54jUZ3NBx0asevCYHDXn45NdFidsCCKK
x3t5QmokI+Jlg8uIgT61X4IrPChgWdyo2QG8nGOnjX6f7xbh6dDBUGyR0ncu
mE1MpVDKZkgQNSJVGTayms44+ziu88u/vJGNqW9o4YorJdSo7WHe86RNY3i8
K2VQ4+mtDAurQKPfEGXGRxN9Sq1jlR5bksCzI/NDmT+9vZmEoFpfkmsutdNT
qQmZTUvpNeJrYhQeCYGRjE7rzB1soe5Y5gy9IOfOxt3ig7RqdtDpDlwR9yKO
a63t9LmZQ6VegM2jBJQOImBmJTuR1O6uu6sSkDOkpmVAHArpW45OBwl4ERVS
opw5/MDF5iT2MHHgjQvENk2K/Um0DdvfNTwsRmpYiOgM3HnFYSlLzHIxqeIW
0R5oF8fwV04nxiLinXxIh6cpatcRtEwGyFPuu7GmvahXhf303AtwBaFJsQWH
kkR4Hugc+X4FljrqAN1FvnmG+NiNHQNzFmv7EGluzwZNZpOj86axEJuvpWiL
AZmfjiA1Lnd86E3vC7ERQhM8xBtAqKp8Z1Qg85SOcPdwI6d+u7lL5oj5ZNh9
2gv0665QKnX6ubL0ZlerSWw293iaq0PuivZ7QWEvwu3DaLbGrtvtFfzAIQnJ
NrvP2TV6VEw35vBPCVGzCiAjAbq7RptLl1NGgngpibg3MBy7OreHl7N90z5V
fhF0erngg9smm2odtuwFevDeUBCnEteDnoaof+LOyw49/dZkG4vqyPx67HjF
3s6FeNtzHPwE5ISz5gEaUT6Dl3cAzBKLv+xSlTQD/UeGhPxyvo1GtKbpzCLh
nnaYxB41Dy6jcgZkaEWUuV/gNhKxlEQfcNaHg7ABXyauYqjxbXRoCaKbfjIR
WBiCLcW4bhDqJwd4yKXTfQWkigg9z5J3/wuNVmob949fhtBWh1kzZGr6jEWC
a+IRDxeStnAoEsz11luSDLaSuouQk26XkUOtZcj5KA+pSsjmKqQ4AjwJ7QyX
ioxaFo89/EgyzCrOiQ2GA5EsCS0TR9awWdjKeqMXzu/HZplJeULYkwv2cKPC
1Kr9hIdBvcwQVw6OpJLOVPAXb/wpG4ufhRINaZzGqEM1xG3kiauIp87rhqr/
CCYSqbct/QhrfrRefupAq77852bQS3GFMEh3rerXDchdLHgKEOOIsbKNOC2V
M+8PpfgromYftA7RaVaRnPQT7G4+jOe7uQZVcsj72x234gLSSXy9KEDTrLIb
etIVYm+Y6Bl77sZTi3+rsdTI8hxljrBHOtBh2usYu4CxL6smMaofKcK6zj8o
a0+kmL8ZPrQ42fnTg8KwdQG6X8IDU+1xJVHxgObUpTJ9aS4YTaU5/uon3NZ9
8+kCTQh/JRJHrEdTvPadDfqSSeDB614Kl9FDDQPxiK2cGZGqc7AX2aL/qhOw
NLL0QOhkaxShcGyMVue0jHLpmPCL4MeeOsdkJxk99hH1ZeyeKOFrujexkqb5
Dah79ew5IkhhbW31ltu8TcC0GgJ0eiL9tVSCBvAlvyDwHiIh8fj/zom03tmm
CXJVz6tIm/2sVTAno/l5xkMz5jHF7y8pMiIf5hCdY/REF1uzKGRwu67VRiDo
/Q9GP3wvbP1iAABZ6jVBKfIeYpDIOmHIWAwjIoYltRz2tyTGq1Dv50bEDRF/
vUKO1dAEKCLYl+MvV0cN3EVfZO+hrK6qYIS+4ipjkySQ23REB1M8ISfRvrHJ
KE0KomnkiPr+Re9oNIK2VA1xyy1cSaxtVq1bjF6u0CTHnClVcC2zuAPRLoQQ
YsrLmFrR7UpBjSIkDnI6vst5M2lzIPxdzHp5mZiXjmFMuVonTvyzBehdGJ13
tK+Jv0lDXOsWeBGdLCIu5GOwNyK762YvgLyLxcJrkIKP3liXy6QXIwEEaVl2
5wu3xXA2X/rQjSkBgH6VX1TmRfIsbZGx/u74NaceXDR+Q52bV7Il/v0KlNfW
YjVMHiFmAHc//M4R1uly4pssmouabz9WS45QjAdrxZpWToECymaUXWxBj1L6
QBvwJd9+8keHQtuuGRy08acih8OGpFPbm70E8AWD4+z3Ivq8onbKFnzaWCPO
M9qVGuz98vxYqH6CCx6Wjz7bN/W6he5V+AUCD84RLAPdGj4doYsUoT6SHZ02
gLg/XGQKxXZPTtCkgpEzF/arZedOQWC3iCI/McAY3He1a5qWGGIagOYfl95Z
tYIIJLhfeyQVn1QLQ7/UKSQLx4vCJIog+SF7n4MmDaw11t4vXU5IbGL3f+ev
GcZpwJzm1d4FZqVW7FeNc95L/gkFkEQVOh28NtEp1yFcRJkWaKorO56H3J51
gcoIEkfrV5YWFQ5q/Lsu8No8aFzU/uHUGqwy2Ni/NE2QFDrLmp5mpTrChuws
61sHOOZTgmRr8WutDz+56J1J0fyBlgtIUumSgm/ALU9wFamVXNh6U7VGMBTU
eT65QPKrTPAjLLinl8/CLDvYYuLABCdnk+eU1z++v4eKeg6JapVYPaxHf4q7
gckS8LKmVSo6OdeT+Bgc+dgKWBvVo15UxxHilfpLBSPQYozPh2XFZHlKfFMJ
4jE2Soctgsk8rg2jG5tL5UGo7JdqzbgSZXf8dzxtq8ztQUjanqbShc2jPgYv
s+ih0/4uKmlTUHNkLui2hjNlcYJ/kZzES3/Xqf0WfHaZwT3L87QZwamLq/TG
1ttYwlF4vFKX/D8xcPl86XJnWArqG3g1LNzW+Oa9WNOALllbbT75VUqBF/5F
+ornCIBE3RoX+C6icg4rj5urvqBeJKjt4nsf4hnPWA3r3AGblnJHGUcmQcXU
jdv0Xz6aX6dp+36R87SV0/TT2bOYUFUm3OxWHU2+mwjy/NjRa/5TisWzTlNQ
MhJFItDxF2yyjNgDk1D4PwK+7cyUj1e7ataKTC2wvedm0+mGv+3u6eu5SqUu
tfJiPJON2FJZS3FERu1dfh9Zqcz9te2XrMoT60OqRvZDVgDNwljf3973kUwo
gXfqIJOYPhNA8CeZ55ahlTrDLujMUWKTK5a/psZYMSyOWaGnypF3oV1XoEji
in3qP+4RNv9KdSb3L/TxQgP9U0hWtY8C40fuJHX8gPgiwMVyQTC8hsT3KpYH
z5c38WHvFFuq6dPpJ70SVIxUE6S6+sxA0rM64Rqd7mFdHRraSolCJjkyrG0N
CC5ojq5md/F1sbdLgbmEIvICFqHIcNKLpVb/7bGGHtRjJ1PnS3QqzHlNCNPD
qOAxECe2/PaAwi3WFDNYM1zYy2EUd4YSUWiw/fJZvBwgo1MbZLBI/c8Is6kq
dlD0k4zaML3WrVDIXQQYcVcBoSWt8WzF7Iso+7ydlXPvNYlEE0zEXZFWHKM3
FSuyousmF+fpseIL6SAbD1OzK6xoHfeT4Y3LOCJGeVdQigmqfIZvSwSsJZ5a
/PLVv89+Jl5XHVwcMO31JWYfhygdtxUrq8xQ9eowSwGvjTpxJ0DRyJ/C8EsS
yzFvaB7JB8ustaS/CQTVXwrwPMSkWI0W5XGgtdFT2NF+MvEZZlEh1THoP1Jo
WIw48xISjfOZRl7JDEA1JiNiHMY0xGVDBlldZqWIudUbP3yQc4hAUqvL1Pd4
FwAPIJvdGQ1hBMW0TFSFXshKXEZo22EREr4qAI73Fku9SvxR+4cqYOakv3hc
0pNyw/rSWKWup8QoJzuU+bNjYdauw1vAv6hF8GMLP3wdGfdS3a691FdVffLd
dzOrwR3pfETgLGPSWSFdxKvQT+x0UZXN8rPv2xRVTaNXO/AdHudTDy4yUiST
dYB20y3ggMpqSfpPke8FYpFlNnuN6eoF+Mpaf+ma9Cv8NAj2WlOiwWDp/+Yx
cOCsoYLICWz9H/+Id1cCid63kKyOUQutrG3jMUnZ0K/votn6CnLM8ytt+Uhs
BcWC2ySelIsyJxxbx8pIzk7NZSKc9weyocfPR1XzVghrerDvK1PCviC366Wy
7PaGPXL+TGumvM4s22oDeriXP2UmvjCYSozoF3qNf0lMRdnF9xN49tD4KzkD
D5D3gIjC1M8/KIONzj/kI+3HUW8rYgkCMLCCbYiD5atXHjjHmCz1h7s90zVg
KCIh6gTd95y+ogonqA7dqmM41m8owzKTYWVpjXjkwb0IcSKK+7/sQN7HqeVz
fhoTHY0XmdXTvnX8zvimmDAPO1LcPn9JPj+HwP7ZV48mTXZXa/okjjQaP0Zr
iAKxvqcEhbW9Y78iL0myjwjxNjHKlUMA4wDJP05DDKqf2MZs2RXgyuNmuXyO
rQAPp1fKcgdf+FPMF5W/72Qu1UNj35cQHaPbhjpYrwLhAmWFrVk0KfY+ephb
JYLzuFReIG88ElI8hyIzXn3okbBYXwxTqU3dFV9OAiVLxbsr6vn7rvnMXo07
UpFVy7HJcvypEThtriGdTW18kNa28TScaWArAg0WnXdCfeTrLi/XBcdfe5GU
xSBSa4b7+dym2DUAMN7OIu2BuKTZRiQdvMWX/4goxX8hBe4+ctSO+DI672RO
GdkcSg15lygZcQofECiteNGxjCgm46l/iXmWZ7EAwNc+FP+9KECtm0CLy/1P
0hAKmaZcifHLxSBPu94UC6iaoLgq/Bl2hg6bYs/cxr6x433RWWQ1i9FTUEuD
EE/RyAdg/gLH/O6kwzF8IgZLwbEPdVWTgKCO7NbQ94v4cNzZGXDKxwLEBqK/
Bg2Fzv2xG7EYyzVVlH+y2utZpjT7EQlkRukWyWOLs3OJwF4P9aVwQyRcF2/j
DYa5tJHdyLsqu0u2wAUouyoLFLVYqYUXR7VPDwM96K+B+gL4zyY1bhe1Vx0t
uXLV/8RRRTXgwtpbk9XWMr48mWWzcDILG10tXY1+USwBJqr89GTcFvJel+ou
K0gbOqVMn6OY+ercWBKcNFo9Wt9FVfydWHmjHhLntplufZQ+IG6IF1qYQsEF
zAvZEJrNZWH8hnzK6En9dTJmwcu6swCFN52JhVHcNzwoWi/O1aM3Cj8KZWFq
yxrDKMv4MYz/tUQtaI8AiQqo+82eDIyQOOhECuSEN1zZl3jD3DCV2zHRpXQM
T+ySWWbDUREkRTMMIS8QmvnlSGNb24rqWTxi2SLVg1Q3QEogT/M91SnCS4PX
57CI+35C7wZM+TC0qeTFUsOuUInnur/AP1Z6UvvlY6jiRcDdJYmsYYcHuQGL
31m1feSQ/nuNV+Ka/haLD4AFnNuou0yXA30npAogEAsWZdyrfx87NIpOC3pQ
TgaWfmY85q51nU5gpSBPFWB2vClN/W/TFmV7I7FyxmS1IoQPijriipwtzUc6
u5caQuMIUfUFtWV/n8MBb2wenU1kYF4zAHqf1zJIt31ZKYSilrY5eIWnjUsY
ayakcNhva5KPbhcw+aj2mPepNoLs8B6omYb8ra3bhnyaKpD80Evhqni/ByFO
7WSWeNcwYa3J/Ny6eJgotmTdgtN+rxexXIGMlO29Cp841hPpogWB+VzPnx5L
gzXP1lXTIW4oN5WX8oMncg0Ve28TKD+fYODKmOU3yV7G8M/Pwla147WWOPSE
a1feX+8s8BaLKdeDLK9pjXJ4yzhjU34d9QjgZ/BiWefPrO4jWrwpcIE+r86t
xMBx13135ycRCI5PVB1pfT7XKzrHxbjd7r6UtMtcW3ETXsB5OFBmAXqu8P1+
CXSz/quFnNMMsoeRo+818lrWVDXmwbbpwAhJRYDpGGtNnmfesF/dLOuikZHG
XLMCdfvLtIY0rz+TG7NXHXEwc8LCuovdVF8FblkoZy3z7V9GzivJ1LIiZG+T
3EvOLJZs0bCECq0V5JfEuDT7TO6AdIA497I5XJEnpJ1u8EwZyFR8k20eYOgg
dZqdu/QcMmu1YvRR4yhisTDY6z4vIGAtjGhLR3sKVKKHowpICkeTf0517/e8
g2aEVc6hl/SYCu1yaRUzbFrVCabmj4mC8OaEelmTAtr3E7ajZl+cO6XYnP7V
Z5BSQVhMgXkIKeCMheD1Lq5n8FHOIDtctPGwDR+E6d07aOszzDIcKJgG9AZC
WmnSe1+LUkDDgnUaWoSYMBmF2caMls2AaWfVueH8l9VBatBPOdHbJ6BE0k2Q
ZZHpsWrlw/xEogS4B9uv6ZZlg5jUFN4S0+/82vAqN974X9yC18ypxl2dmS1X
Fa8/7da4BtuvFoKp39e66T8hfZ5QNxf3pQlXBhKV3No3tpo9Addush4NXG6T
ArEtyPIXSN9v/NmaymuWsZpkcbRtS7ap61yh2/4WCERNR8ltK1NPsCCrKX3t
35Y0swS/1NtPPa0SmA7kkwhANSlZ3tKYyhPt7dWKG+WNokf0wu2f0Wa8eCR9
rYwZKJ7CPuEgBjNsDR8ipKn5WkQfszmdlxvmTe3fxGl+w/ZhA33N2MVw3ssJ
voeIlPGUghBLSPg0GLzeAQNDHpULhFbNMMia0WfynZO/6j2XYl5QWFMxK5JL
ar+4ZG5cQ2+xM/bOoqnG5HGqGJq1I4N76eF4NE+o7OUYM9apewLB5WxMwBf9
dvK2+mUVyn/+6No1h/6aQ8z/EQhtzAq/8Z/buabULFHWZ/NRiVJ90Om/IxAP
DERvHJbVlkzrg/k/Siw3SPcqgUDFf1TJSKYTMUpSjJs/gyOmlG7Wm//2UI0T
9Rxg/I+PR2pogX1fj4Wur7iDO/hkQSB2UTfeCt8NOngpfwLIibC+KlnHFMEJ
Vj9n4bPISVN4XOiSkELQBIvKSsC3n8iJAXK3vZoRLEunKZrU6zJ21xjkcbJT
X0Fvm2XA8wNZSHkwZrogAZB2qtmREceLiTJyVnstPHH3F3SjGl2JCiXBH4m7
ys73fIenhStJaB6j0rpnkeRIffE/jyXU33znMcvkcPrJYj/FUCdHdYsZdpdF
afJXCUVJrJbAhsRonHE5/nBieSTF1Aq2anIlKUEjbyF1KB+MitpS8/RULM3Q
jHZzA+KHigQLzNBPbPs9yOuo9iJfRxLTVFXCYTMyiYKX1ug+MDZYGWmSUVHJ
rFN/fvIkqIzXqbRlaMAGNIRiZvlhGy9rg6NgC9wAiNq+3/hTIFGgrcLDjCp2
UV8ZEkr2mS5JlSZsqmLCPlOXrVrRDAr31/6ESuGwecqtbL5eqNIt6/TlRsWp
J/T+57MISmnez8fxA4WhcrcHr92rkxbJUHt6quFuNmthO1NAR2tkEkVFQ5Sv
inCt3LDer2/nP+oCxTKUGmt9/MMeSp+MgMYttRPNNXHpj44YTUgdIzQlOzv2
qt02BQnYu7DoM6QQlcYpOYYhRVHOEHM18tEaiiIJZTLfbiVlJ/6E5g3A3DqX
xua6dZfBXEiUaSdgHBKfTmXqpvmuipHb3CDfgF8kLTGg0LRJMGYzLF3Sf0wB
VaInGfBMp9dazqIyVlYlIzAUrbs1rFsXT0Jtd1oqyCOVS77k5ctLPS6hi0Uz
LcyXvPpruDE3yu9/kiTN5wqZuof2a6Pe1Wpy42WdCxoqUSvVMRXoVJG1n0Vn
qVTXAMBs3G/aA98IvoXLW37RaxS2S1RJjziPCZvslgx1Wd7IoJ4yeeoeHhGa
XcRUDt1LNIhirLqddTuhKTp5yxfDMAsQ/VBwGleMO5rgh9NvYAvpgPMXUDzO
rpMqLwisNg8gksInuxwmKwR/gqVzv4TCvhZR1L4EtF2qsbG3bljUmv1X+HTE
Z/2rARfNQlPmqJwwRWqNwT2bJkXCsAXIoy5jAgBLXGz1+ZZqdp/wz+JFaOZb
ZCG6+8pSbFEPjDNWDDHrkwo8AZvhIvCDI22RG2yaKpFEFkAzC/Ftjz4lG+3N
0fHWXDDmm4B1UxcXesELg1JU0XN5Nv+8GBC0TsazZVCNcw1VtVRLt173qSt4
WkWTaMBYy52pyit8Qv/Qe60EDr+o7LlY9WgrVXkBLE/9eEFk2mZgzXdelaP6
/lOZsLs91OP1LXdmdAwObK7l0mR6G+qex2cAf1iLQpAG5pnL3/alq6Wvgnak
4S0iB5HluCfjhmVQ03ZH4Bin+k1v+bPTS0zIeZAy5wfGeKxweIQVSDt4/Qt5
R2NFIyb+gUtyg3Xtstfo8ZC7QVXgabL2osTYXlNVwppw1xfEEqxU/dv0/cmi
hhW6TWF+xNf6FlzeRYsykAx2oUko6MPhv30nbHHGQB0J/pstxCHn69PC00Fn
ka1OLG087lLGS1yPEWPByUq1mx1x8n4GdthY1kUOG6RoYOUCTAA8vsBGzcEj
5xRFXs67qttX2tb99mqeul7r64e8bo555zhlaDVA1zCAy0jTAthBx+ofKSsS
TNR0vdg0YNyhA0xcetGOyk0r7zVKZo8xf1ZHm/dxHzibupt9zBOZFbI2KX3X
cTsipDWVD7oVqbB8k1rjFZrzFJ1I/o2M6tnq25NdZwzJaBiFp1Nw5UIxxyhY
UhQvHM4He0MYiUnjv2vKE1gij6VKhxrWT1Asnebsf1uHrUy0MLMEKfovVPpv
QL8mLDmoAMhyc7Cu8JTsbWW4S7bLvK5F5jADthTs8QQI5fKzfKdtayI94n6E
ZFxjRQCP37QBJPf3Bz97wAL42iMQgQZu1bA4KSkOQd0BSCbrBoLW9ODsPlcN
i8naC4KMHx7xgxvbzU1yiUAqBH8DBnl6uGb8JKHPXk73secaMpL3eotmE80r
JD9lxzwniebUHBENj8NO1cTyY8IzJSMMZoWhAhBlb0GRuokRfhQC7d/WZKRj
5r0S1bNoMaicMKdjav7ttGL3+RkJS6APgZMZjvTgXFOcvaPYaxHop6FZMNfc
IMWsdD5/sJUUCm0muC+wX6F1ksFF5sHaWbv3HVwK/68yOb6Go5hKX+ZTxKwb
zDgFOFFFqUafPQChPsRB2txlAh7VhNUkrMWO/gLckMudu/s3dPIJ+ecToDlr
tjLxhadyMU0ttLHLYOQhpxxjHycByjKPGPGiMX0YYymJ8lo5szrZS2iNzROP
L+zmVnAhdQXUQczaey6FRD4cN4OoXYQQHzGeSdACqJOcjBnZEShWksT9ntLH
HL5fdlhWQuCIgL4eIgT7TO9qcjAt3WWUWV2TCWCUl7W9EPbWOUwhtEuqYof+
3orU0MHa82inYxT1fEa/okDs3vPjjEtyFJcJyE7klnhN0MVga//IjGiOQ7aT
guIfl0wDIwvjxcDWuZ9D494KsLCEP9xDzyYdNwx4/Ny72aaQNlSBGEcBHhIS
fyta+Iz6R26ay44hkRdR1ZY2dypjreE3D1b+uKiWiooWfYfQs3RLJgEDi1PB
l4eLVjPWhjPAQaL6KiC2cxJkZc36maLT6Af/ArXZPtJZTO9bDrTh3Zlxl7Al
cCQOO1u5duPUtqLDEDzkaocCNbfqlLiZbpl6Tm+g8k59ERnYktrnO1ZfrcWA
gQb6hCkYN+XN+iiRsrLatvxAcYratUTb9AFD0C9+7iB7j+85tuh5GqIIOPy7
rsUPi/o5rfq0lY3M9LV+XoSKiNuihNuvdP/ya86QlY2pcKfJMRHNCG/GiVo/
qLeHYqcW4XVeGj+0tCISpz51qXQDZ01KT3DC9wTf+ivUl1kmHhxt9Bxkpvek
Gd//YAc/wH40EkzU4QtMWPPZkS5OVs5Ep2rZTC1EwkQM6XBYtZlEoMI5QAtS
608Swk6EJsfI9rwLpAs0j8tR9uDGrd304JVRjprTPbX2kpn2oCJIbh1z5agb
/THTFeiVCJXFN9c7KKrKH2szSuwvO4XE+kw0NN1E8ZrDUJXJMZZSQGMEJuGG
iIGKMpgItN0NVEodZZhXXBNYLDHwXD51P8YrkfVEZ6OFel1yk5Fj9Xu3ns0z
AqqLv3GMUIGpt9nKxzvb4/KW0JncYrgNdJeoUfCRfeD0XK1acnQatPUTl1Rw
haBt92baeqw0isi5xoN9/j29Nd6gO9ng1BPDGEn4qvqTK7vH9CJBXQavJqL9
13QY8KxbtSSD+886Fy+ZDEAbmRcPuwSxPkYwjqDvtbGKJ61zyXEOZtWoT53S
5sEWFoMzt32MFl+TtyBcGbL7l6gy05vSOOWKQzuAxCMCei/fPK284dKFm6We
mf2AW2GkdPw8lLovGD/+kZQriKTPD3rqny0QNBef+smxdRXhwX6vmfkYKKoS
c41Pi9Es8W72DMCypF9yEMpGshXDkqzGh5T7ZY3IPFKmyts/KnkZsWgFv8rn
mJhaHd7a5wBIyP9G9qHFMQE0Z1ec0871oxhKg8El781uHkg0iNULV1cW3dhg
AZsCp3BwiQ/qNlh+OJxVbGI6zeQf97zb5h91dBFbY3TI0CmQyPLS07kuX0IF
OUkxjCfHtIXeCvIrhxJDe6qejx+PXDzub0aNyTE9vmIoktQJfMFM0taTiBmT
4zotVBS2JlOFVuwwB5cBK/uzPm6D3EuVeta6dJ5v3BZaaTlhq9EsmkWgcjxp
4YH4tvI6uNJpeKLeFnxe+eqNy2Xw84Zf/ej5Zkd8bxyDT+0QLpYWoGbpn12s
0oauuuekj15Fg6aPpMAuW4mQLa10WY0sPDGwg/7MZVZHe7ggLP62xYiKUWOc
pejAK6ka+Si2x2pgXvyFMD4480fzGvgKfqaOOu6yTJBfk90rcLBCEwaF5Mvz
f6m+W+/KbyE+tMUcW9G1CMjUgMvS5ks4dTU38IYN1Z0G5rpRat8UsSvAd3M9
E+O1pB5HJbtfVhcDb+gg0JSTjxtB/MF43QLpYadMXcKzn6VKOL6Di52/AQT+
jli3l32+viG/idpPX+4Gst+yQ4xTurxSUULzF6a16vMLwzS3LqMCQvlgS+Hx
TsvO3ApIqjZ5XZBx5/TUZ2f1tpIAUX3sL0uww+AtLsKnfeNwDEVMbYp+n4aa
dRiOgPirSOGvtB7pwT96BcljTy+3ayasAkHkx9uQRsNERxcvRd2ywkVTpJRj
djkxNxCaPIm579UWGQaLo12/u/Z0uIkAMbVN/ta6RF+9NcrIXEPqK5Cr8H8P
LazbspSoc08JWzPLCtdWrbVo08u8Io2hF4B8LbzP6RSW3mS5YMVJNoS+NSU9
kgDivpdbj2Peo5sqW0abUakUhX3qjkg0nGzjk6B5/cj09rKx0R3Fq4V6difo
NTMIx4ZIKc4eI0PymmrTqFBZV7utdZxPQJyiWJsX+eRUSS/3u5Axp5kFuSqX
F5oWXrgUdY0lKsUSTbf2N+UjoK8bQX3LWosEESVBom0FhAweyfNcgJIzrPwt
THuDYBmsazXvZOR30XeqrbuMK0FD641Kfzd4L3piXK6oC5Q5R5tEZEIurX3i
RHUr6l0GUVon3yg+IeRZP1OVJKj4trXtvrzLetq8XSau9H5FfVw461o5/Yde
5DayskLYZv8rOK6y/3o9XZvWSHL8f0uC3JdhGDDuQVQXET8xrUYMiH5pHnZf
b5/y0cfWSzsXaD9NvKNSN7t4m/xTFQl527brs8V5ecF0o4rlldg4lIPJm27w
NKHkaCd6V8MUrZmNS9EJuL9QtacRzzA5jWLrwNXjEVDiknzrEY+QulokPXto
iTfkhJcGV+zCcu6eF6TWbfV/W1WOAkv2rOfvINIXgqqEmPwWnetjLlqCorPO
UL9NQ2/LkGnYC9QgZ0szUEmEysSY+EwkeALW23CHQGz9zRL0G4Tw+ctrP1w9
9HzejRo92fU6W8btowVb+oN6cx6Xsj+lLsHgMDob+Uucc1VmEL9VTxvn4R6B
pz0V4wItlKhtJSca3qpb98EUj8Khep24YMn4rYfVK+uwBCQ6CXoJ9RV8Pu0H
gLUfDD3PVFzmk7NrR7BsOmWCTZjKl4LpGdY+KFLjAhKDEjem4dZiAFeeWjF8
GrLGZYpqP1svNDXr00tURS/5zONw/1V8NIDPbZOkQbuBCy/3PVRKyOfNRo0X
MsAJV8/a12JkKgh1J1J84Nuyr2dx3bB/Pu3zNWGGiPMkPzcBiZp9tHkqKk8p
qN8PgSOYnI7h4BgZrUhc6ZCMDA6rHgyKUuEakSNBvChgoP5YYktUJAR5XDF7
ZKXb0OmxbD53DGbKBGzdqT3ETenxRW7IV+kvnflfxWENZdMBYrrzcVdWUMqP
LVsCm1mZk12IfWLyJGA2mfE7w8NnOlD20OGrl2mtgC+M6g1ymQ7ejgdE/Z2Z
CgSxBX+V1yW5+8bVoXVzEvxU22HS910p77NYTTzip5eCEidjcU7PjalAYs9S
IWUYEdUuzCmnB48Mz7zHqFsZ/wG8oYoa6n2khbco3bE8fNybw6NdJtXtwHLA
sfgv6/w0wievzCMdDT3nJVHo+tWj1iRx3LqAjnr+lV5JD9cfUMj155yFsUz1
rkNqAulQ0nuv4spF2/kd4s90ImcXiof26QLlNQMIvNzv9BGWGq9awfm5DRY2
fLwOfJ5WGm51oC6CWYPUDkAmuoHYBq3NksKO0/8/R3jf5pTcdkuGQKktLwPU
YVuIuUZVlOMVUvJ6+PklhMm4Eunw65xsvtDiki2DuTfD5/4dFHCp4sX9wkbc
bYQI0yydjZh94sASeEeMGYbMaParuHL2YXxMgxRG5P4zHyT1SLZjxwq2cG6U
rUK1I+cK/iQEvYo9Ks6OPAMXRPpdfaBIpJMnzjhFb0nMk2VjKIbF2Kso0s/S
DVPh1atxPCaJ3/cHNjQVLrmzNIKdkIM8HJJfgVeXkIAK1Oky2PyQ2JQGns0E
k80mE36fOwlrN1ymaSF3bmygnDGan0Zh5esUxHrdbVZmmiLEZPr4YwYRgXWi
YLmFDd045R1308/SrgXZrHjMCVajSwNwNc0qZDD72kGVUqdLnjfeV9dyRNX5
CGory8Kb7CHRwCrzE61soIUAJwYZgxPzBi6l/vNA4IBYM3xc09SUHyQiZ/u2
x8tfvCV1MGPbWw7/gTLQWhdLaM1A1iRuno9Bj/pn1scUi6BWpCY8d227wbdS
+yKD992BrwWkrMMBzfN91YI756WVBLVBgqq40hHOpVLavFdVwrrrtJvY/Suq
IMz2lR1XkkEa4dAbWKux39Y5NgYGuFNrDklSrWvvoVmet5yshSGXVZjgmOSL
WpklQikPvpWTO79x9NjO6aB0bnfNU6neCgWITegK7GSHQUp9c5d8mYrQJrlH
+QVi0fmb1XflnD1jEJwX6YrFQK1WSKOAMCPsJ7Marhgg0ZddU23wvX+HRRFd
CYlPqcu53ocjVeEZqgxRy5qaiLfJpHWmbUvsj0dvzpuKLLYbk1HXiJo8hrAN
5Kzb0X4A7+ySxd3VcHl0SRrTAV0WmP7F0ABCRBfwWqPKHJr0QD5mQptftvMN
O860Cz2baoi75bex+bi5n0cts5eyksfMuEIQP1WmFBhwKc6oFg0mi8Jb3gWd
/PuudovzUHipRBASFnyLD7dCkWN78wo87o4ZlgttH3qddFtGs4aCnsbu14J6
BVX7P61wD/6WGTrriIECvfJZjr2iGMy8g8zdYE55n0Zdo9pKHGeX2IhZKEM8
maJVQHctADMNctY08uU/uBzYIpE9HwaWv5P5JLwERPbGWk9kmjJI254wl9og
114m1hkXR/IxkC3LMunTKosBlxCGrqc0D0Cez3a0osLjkvA6YCWk3lxH48jZ
ZP9KgtnSHUZUm0NMKxJrHg0Tzm5Ww7JRT5LYf9pOyU3SwIuAS1ay8efALQ5P
NQZQSq/Nlq0IMAFBjLhptDmDjW7OGRTNU0OxthfMpwrpV/OK2UD6X/LaBxjC
ZcUrey0mEr/VcWicUFsZpMfjclXl9c7RbvO456UQ2d4zr9l/zMlVAqG6qJxV
4YOB+Su3LP6QTZIEToEcTSaywq58r2Z/qrG/BAM/lA4fQEnfbizROtC8Gp5L
Y/G18DNjGbpyE9n34F1JFEYao7DSJEn8iH79hQAp396vpZYGvj2apkQ8SuO2
TO0k6+RVKRS0h2bNy0Xr8Wx52HbO3FCYPUBRISi/fVbB6fJukH2fHQZQDK3k
+KsHVWJaj54Admu2+Yz7fSRd1IrhDzamGTMmq33LwUpuCzp0ibB7YqenZMp4
+BYGrH42T3ziDfjKBrdRMal9VFGFVMApeCWphS9mJPnbkRBFnekC55/m9Kzv
TrX+O+e/MXXsiwdyktZxrlrbDWw4Yh3sTXsZxEx/t0BmHg4LwgkJCYWIbM/U
oovRbqycloY43DvkU75B1yWRAIMeetBpYdKMoJcnazKKc+TWzzBiP7UzRHE6
2egpaV8G0byWmG5FJWbI3in7ow8NgCnSzbIty+v7OVVQYYI2ByZO84u7t6dB
9FvaM9a6RKm0Rq031hGrAqS5TvNv/LZRLHi+V7ZeP8fjMbyGZ5WBTmpS+c03
g8p2ZJ0KIzP0HK8xZB/TvJ6pcfd5yapC9gfo8A3P4S+XJVPbrC+Y31z8UjJr
MLvl0NE4NVl2dAgENj2VBpNJJyPi6HCbcWzQCJ+On2U9KaX4hMvtzsvKkMtQ
rUh7Md+fSavZwjpKJ+ytQbJ9aN5/wMg7HgUv8MMEwP7bRc7ySoSGoamhQxQ2
VN8fUagkl5fpITylgZNIQ/fxYPDG9zEGvo0de+zI9KkJl0RI2SLC1kUSNstW
xalvrMkdsg6YrsLvYE958yH6+y3bRzQKYk9wYF9AwEsc0u5c0EY0DiaOLQ52
ONB0ZvFCUnVX0KzXwKcPlrVVs3CxZmvumYa6FLAfQTuFPh5z0j/s951cCIUH
HzTuzzw4KI27XQy26WGhxysGXYPwaUrBcT63rjZnH4isw8VDJZMIrP7qbnHB
YxUp3Z+pxt3UrmAC77yoLOT1oCKooWPXtT05EmolVexwM9NkIzuntx69lhEI
E7RfgbC/lqiDCDLFWbdP6CL42LdhT6cCmQ+57XDD6iP0ft67A/9dZwa8x1Us
WBCpk4cD49ISQ6AonJHsIKgUFPIU6BEEU+qL6ID5s/cuw6aoRjTBYfeofKgj
TRYKukf2yehFHFD2sNGxPGsQddbuCzn7Aj7Ac2Ldm/CaUNFudis1QM4eGilN
OzyocDKxtpZhfBFMECRdByxYkrlvJ+tKK6Rpc9+UQmrxu/nzsHkERPFa6WCd
567iS4VRBr+M9KoQPE9aDypQmg5tWb9GZb76ijtB46TAg6NTMeWedEUrPQYt
B2+lKyK3Omdxigb6fPYtGqtg41fa0zd1ujLjIQWLNZKxzQeaGM3ODHiiM5Ff
wkcM6ADbu+PJ55mR4hJeKtZpHcgXBqtggeIp3U24SIU1ZNXFjJSUqNYsEXiU
wO80o7Q+LTYeihE+kke1co2Apj+s9bhWD3WtA5wyNLgqArG1bafuJJLc5Sfr
SP8Gu83ghIX2r/23nVp0G2+WzpXG9/KlTjQL+gli1vG/1cLwJAOMSacRhGCg
9GI6vgSVNTCaVnl1+xkcQ2BWxKB+593mAaWdRUkHMMYWPSsAhATJ14hS7KqD
C3Nm8V3qrSbUFQgKkXmYPZthcgGKJvtzFfi7XZ3H/N+fXLoSYZc+P+FQa+kO
/TowtHxuAiriSLaQ74x6rvnPZGjjCFxYf2M7jxKcmXncnrjfdeiHxR2AuBBA
bpXkqfo37IWXzZiye+TIk2xCEJO02SoeKQdwngvvbhmfAlvFkrObQIZSMXfw
bwfn1GBGHso9q9JSWaKSacBt2nLdVYkddlxu14vctjGjPJ7+RtsSfW9+oF5k
+1V0JuaCzLTF2vi07qrE9zxGu4Suj4au9X0PQshZU2mbYoNnIUdg5y4H0Ld7
9aZduJz95pNrPE62c5Shhjy25xo6d62nWxpA050c/g4+GtWN6ZgzC7pxCZUE
WWlSevmHsjQeW30VPaF5PleRD5B28Vha25PXMNNeb4uneN6BaiZ1M35PlWPG
0RplLMtd/4/T9yI0nY0bphxaEqEVLfnhe+ZK4qKPtVZqyyIyBfIRgBC4AA+h
3aHm4+JChU/BAPTILYTsxklFjsO3xFPXJ2R9HGAUd1OR+7gQyhg3PtxRRKbI
XQucCyPyIVK21r8o5kjco6w+bNy6PskaVtKmpsVmNcm1KoHhsQawrF2UiaN/
gPE8uT7v68qZEaU9i6NpEE6eK6YHDE/DgYrcB2T1t8Kc6ziE54nv4esmyqRU
YKs+0JYNxI9RW7K4DEmVTIM25mrQVc27HIc7AU+EHe44wsM+wbVtCxVqDphf
Fw1kC9lUxEicFD25SM5OD2+7GXYylX05JYE7yRhBr4jCaXooCtRqNh29TJDo
2ADUY8rn7MFrZ5VZ8YT+vRS4mI9Og07pqE7m2mGbvpAiDLVkrgGTRM/NmHch
ShMqAMeqiGDxmIg45fdpafR/coH8BkpAfTWvs4lvie+aS7CYg47yBQv31V1p
4e//pDXrxZGORiHtIILKnOYrbEpfL9t2vwqezORryaEFYZfKKAMQs5/DTuQt
2yjhU+xF1ggxa53zX9vzz9/12kb9RZWC7SQC0srKkPaWf+pOOKQ98njYZ6IC
uQHB/UkOWhVKMBLdtXSNqzsSPUxdwrUgpSmhqxKCqyX3UXstumng/ORXx5y/
x2qUV68KPagWbSZlqMcdPCfAghGW9ejeU2YTvzJ2e9y4TIplHPnDWOVTPDj4
HX/3mjV2J8cMHRCt61lHkiTV0gFRUIaY266YpS098vivmc/joR989X/MVEt4
OC5o7xGKNFTBh/ZBFT+rS/juadmcdOJudt2z+yv4ipTp5Q+Y8yuykLgKaVKo
jVU/QibX14jmLhTtQoduxmMn8XxXLxsx0tv3ytsF84JAHFjZrYqUoN1sL/Md
iTcD1zgBPbYRUo4FqGmh1KT5rUMcVMbl3Z68rCF+Nuur4J8fc5B0z/Se6rPK
2uk01OGw5ZEmeMj33pbInHwbYc9l+vWTjyvY8/pcY3lEtyPee6V8yuTtJD7N
Au003CM/j4eNbjBN/BYmdJIC+uM/d6SjwKvYoGYEUsvDC6IzPPoNUj2HHOtV
7BC/I5fFJD7ItQ1PO0bXiWwTcoe48UKrhti0MQmnFvIcgq9HyoqB7dwBvEMA
4zJxpNUHBVVLa9pR0IkapWuU008AVsCcIq+CPIBbPmkTUOUDnte6/w5wrNvd
q2OJM5qmxVVzJowfEH13f/3w46jqdI5QS5Zg72oEFI0tVshy9f51c6soIdZ8
ZkBbThdNnMWUuLehGaILibnWqbpt2P93jisBHZH4AJ6jqegl1LPaAjKt5sCj
hgdzAiSOj+RfC70VPNosDLKsNHXal+V9Lndd2YgQ9qaGY2hrUuyZpLknEEDO
e/Pzse+H8jwn2ulW6zjOVCz2/6M+AyVZQLS5STfhAYOlp3afD1uON26It8dk
1t9iR/ap2rI7ImSSX8JTbplSCskwTpk5CewnYR3VrIt5zUJONlYVHk4OqqTA
vkolyzUY70cPZGK/yqCkz1hEH6ZPlWYuemSUkqJgBEW27ZjO8QgnKA4uBDuA
cWi7nm8vq5ZIBMMtrBsLmTCTvSyIjmbSN2zC1JFFRMZ7LqFXNs+eWeNSYFcW
aS6BTBzaukjm17iPg3LdjyfUozLrQSvye+/aN1RStA/UD8HUOgn2X8Xn0eFQ
pPOMTSy3Fv9Y8uOdTx1/+auwAheXYQPJ8gy+8D5/mm/MdkZundlhpxPmF07a
rio0Odok5RX8Ej94ta172cLrMpoNDm9SHAFQdwR0NX5hzawEpenzElBY9+op
4oBmo0qS51vnho30xQNhk8RxLIFNaCOeyTzy/jFEGuOxG16fpU4C/xj8yHW8
PlR3XE01GfHzBVjOnr0GS9Cuevh5QgORQDMxe8ZoQTM6blqZmDlOmE2i6sEO
qfoViXLmKrUc9uo56WqEGm7+YXleD4wnAkVJ24LHNKjkd/PhHXLOoEP/iVFF
PLu+MHWUsQP4DwFmyTqsmUIfLhHSfNdoe+gkzEnJhXMzoWXEXqmjSJaUhBBC
8vnBbvhTgdjc3CkEkhlkAuTqgJcRVQq/xY8CEFebP0iAdELANI7FV/sV2uFn
sxrH3Bw3VNNjfhMFQqmyRNc1j0u7RkzPfNNTTwonn1JTTShCQUCx5AJGBz8e
Pc/Bx7Ef83X5gCUxKlc8/dafeOGE2FbM1aWkcmANzB+8FK2Ysu/qfy/o5RM9
WPu4/KKUZWFtPo4EbHD1a+Pc1OIt90YEuXPqQ2H2LlBjYjQN5+BVsA4dbZ1i
uRLQ20JtefYsYFXN69vf5nmIcdWyg8mDTzqLm9KmP5ohr7WA4kie4jlaMFKt
yVjgokxMPvK4YQ4jPJPYAEIxcEq70i9GcTy4ExM00rDt9AMM2tjeRojTxJwO
CKYM34h7HA6Arj6wY9jDgfzTPfaZF0F9kYW8Qp7AvpGZqTu1kr1vTzlTqmqM
/CIDYBzLVWRU13D2B286kwbqZRzarQWz++XY4unay18sEOnOUdiAPCBfHISB
uIGlfOkOa3cg4lF++mEipZPAhajRQcuVfQDUJhTPYuA3RQkJsGSQC8GAL0nE
K2oSRB5SPy/xpdNVOEL/e+phjxdDXSpmdkEy7McyWuEqFvYwj/iMrAWn6qYU
/KbvQ8sZW+b7wThUfE9JOY3GJyo0QxioeJic37zmJUqPG+59HqLSj9+u1346
YlvSmhSVRYWpBXGf1ixDVSeIedHA2WlredRuHt+pCM+At4jmM+UVFVkRnJk9
wcYQZbGLop+MpUdsQvc0F4R7i2LwFJ6/3LXb4+nLrvyP6DzH71fKFThUg/zJ
mdGJckd9bJahSVrszMljoDpprgNhVGUD45klqOy34jacvRPOsFOeFVIRyzop
I/y5ob1a6pNjUdG1FrlUeDtNoe55khNpo9SZrwuZ1a4v8Xw4h3zhq6v36XFy
S3sT1NHDVfPqMVAcDCFLT2gHfHvtPkVTUYm5rOBYZjrCAdk3xOIx/7RhhWgn
q2MWIEIx1JSt66vAGmH8UvJSpPSXI7fkRwcLTGtA9gmJBEty0RIrtMT9pjt3
Ox4SCGwyKu8wFvephITJ25fG1xzGCLCpu4KgWFksfHNZYNptEHNjOfnEARsB
Gd2czCPFLpAWoCG5xM6/5Y6Mro1fFd4Ea/HT0FGCAgxnLR7LArq9t5dOEKVP
VYCjeA0StdfoBNJszcxLDFFnTMrJOEGRdrMLGJhNwsxGQe7A+Gm9Ay6PquNw
EDZjIqN/nn0mQvsJoE62n+ZEXraxm4etcRItdNh5oji23RSZaU6pJ/G/2d/0
EfxZSgvfG3FBzuUI+2ZKg+j8rnqshPV+UVNDRKd7caLJXALj6bKKwCgqxkiG
AxCm8YzkVHMh0ZGb6iRixLsI76OBGXFiUoLaTd0IJfd9RFIgNx8IXtAYvIYS
uC1CVPs9+Lt3gltYw6HtkQv+r0kfTkIVAFh8IBulal7ePLx4o7Y3Ri3zjJmh
D92UQcYmbZz6ZHg6iww51fY3/llZRjenaW4vxPFrWecxVuhRZpA2cu7q1e89
8UfppNCaj+TNdLiEOIgSuSPJt9geO1QAGgOB1ZstBzZBQj4H5W6ASbPZZr0h
9I0XKOLmrbzOuaD5sJhUajvjUTH9Ty5UQdTR+lPiJGoAssmq9S7k/I46BCty
F6w6ZFYobirIucD1B2+A94wSRn0ZHrjEre+cvu4MpTvMB3gTioK48nuUiqpR
sLQhUBYYFTf3JxfOTF5KPGyWKyZVO1aLIWOQE0nJEiedBOvuBScVPR2UtHWU
Pxeb+pN2lpgWlnzs5vp8lY/AU2rAybBiQIqFquqS7TCtsFgDwg6wH7zpu1fD
o2/RWwwSfmeQpnM+D/CmUXmAZOo6D7PW9DNZ9ddJhHf1vLBx985M/+ooMMlC
gtCF4VTSMqCbu6Ni/kJ1Lvq1fs+4poQoPiluPeA9T0vFNW8FGdu4YPI/YG3R
gaEhyxD86ErY6bdz9ejJ+4cmy5TG/3S7d15soFuoFPw9tPsMSnC6cJOHN+D8
p9Rx8pfxX6bGf4ztF4KmOuX8wHH2sfqRVH8ONFjwoH/eXEXWK7O3x5c2WQoA
xlPLaQX5EqdmRAm1S3wQlslEXTxP3K/m7AtyM+OFnMaSLCZ5jYUv7cFe7VgX
RegagY3HNWb/QRnTyhcHjeUlMFAWF+OJJIa8pNUKghBTETD2D+Rk9bGTPhNx
qQg8/bknwSLXwOAXvg9atjuIGW8Bt1ZGYXJ5O80SbTCcX36QMyVbk1l5KnGJ
IFxegfF3AcAKcjIcE1wmlMe0dcVGput77dzsl/UVJp5jMV/Au+e9sDeGaRZh
NiVGFRUFGLZEn/f9BWjaovMvJXnWc9yl02Ii5M5JcAuPFNt7pGHDBKmVBQwr
wSEDiLbOBPNHQac1BvADsQ6RZu1KUeAywZz+dh59VzTf7ep675Nx5EStyJSm
po5ZxBBZIiMtxzGirDGn+BkyAkhiz1VVmpOJC2fWW04HnZ+9OPVOwMiQNUIW
o5/ppfu08Gvykb3KTKLO33UCwxWOLyNofn6tXJsLBqu+TrJa4owC1xNQC6sC
Jm+Q+n4KVGownyOXekMI4W3cKBvFThGEqSE7zaECa5egMVi0Ntab5lcB7FJo
Gx8V9UWvDXfQu3W+eDNUWjrWPZwauyEkgPxljs/8qLoesrCxe+joVV9fPGxx
WTnIYuMxSEVJxvoRlnPcCCy6E0rnibIGsdWEbRgGIa5BKa1BWII3wuxWGeV2
i6JUsWb+17hLvFlSZQABigZg6DqHWyjnNWfG8Pz2Ca3fG2rQRvV5ZTVSXRfQ
XMQIX9fG42RN1i9zIDVkOby+pxjspfc1O+NxqgbIf+o42kOQ7RltQJFvlT71
9DOqj1/IRYaLdUIIDc9L+1b2673exI9RRocCQPsi3rxAQHukeJ0Qu4DACu1g
3HZsq+Gil59IeNVJBSa4rAWpiRCm4GQNEHCoPlDdFPxxn5g4tT2t8hf2xZNn
k6pZzBrCdutKn0mErwdqGq+WcV92JmJpI2zNxQCLKI2l2dnGYbzy9Uq4gSmU
FGCu69TGt2net9Z5ROFTqgkd/fIwcBaXUVJQB7p9XnJmW5PoBZa953j3ZDh6
ATNuIo7STHXbOmMq4NBbEpvongqsw8ls+8oBaDx6by+XauUqjjWAjwFnDrMh
CjtwLYX9oGP/sdL77t2zlxphhY0q7A1JIS2EMQJBnCgiE5LJR5HfXlBW3Cxo
EZubP+RgWPrm1KRs86peD87v5uCeLul8O9NeKAxSRFgrWjdAeDHVAT07pYK9
JJu7f/xgv3a/0L2uwr8PP9++7Lrj3I/TWmKiSt2baU6hf2b7QedwWBMR3KRI
KXclXjK5UPPfd1ssQDuHEgP4pJ2zuvsRWB3IfOKME345jWVUg/svkpm3G4Ne
ZXURwSH2GNNJMg9aswK97HKlH2F86bahZFt0YjbPX2C8jcsTSBfWAAnHwjFb
uJUIFPjrbBS/giV+D7jE/BC6kOp7bGadiRcjmGarpAHFyCNko1sOurZHuwGZ
ldyOK72FxWngQu15+s2Zl4wyrKEwFGGxXAWFsqH+1UWYJntFeAtctThauj4d
ue4nEsnfvevvtPiPqkldzlqaN6FnO9JypUpTWIuGEaSceq3xT7TrCBXNkxBk
NlbWXbRzywg1rvv1n/z7dgXpXUmv82zoTewHBtqMXLxg98MkVTz0JaBZsFFn
VmbI6vLIbYqXeEWhE16IWrp5DfF9ePgreOuzf7OxnvimLy0dgtikRJ104MOJ
O7cOqZaz4tlRfgO1Mhrje/UfmMG7ERdGNz0ctknfQVPEuuEE7mni/UOJn7kh
E78SjqU1Nci0PTDXgRC+SI9sWWHsNc2jllDC4L46flFZ8/ICt3oxH0fl6kVr
mEvy3zE/RBo9I3UDsJW8DC68ND/NLqyf7qQhTZ06aCViY3f3ZsaFQLhBxYWD
aCINN9Sd949QGCLPPFblc/DbSoWgvVsWs4o7JyYHdb1fTRBzvm/wzQt/zRYn
0fHffti75W5OIAXdass04D6RCzvBsWDH4oc1+D6R7EN1Mkv2QQ72gMkemOGA
r1sZa0sXQrWtb4KryR2OuG1LH1jvUirZ4SNTUivNAryXue5n0tBRDZRJqGYF
VZqUnBnHCVvWB0107Nek+0n/UOG3GE1ltbY+oyTsZNDSuZPHuAjoHCFEQkmV
06MYfwJMCaC9tKammknsEzei3GBWMOmd+0oPhAB2WmlR8DjnSZvuMWdp7deJ
Nmol5S76IbucwIlr0cpaMkD8RgU77QxPmyZDO1Y6ciZkE+jnrIO1o+3rGoMM
gqfJvODpHRFPJV60eWM22rH4ZUs8279GogBdyOVXvcWD4wf+4nFoI2Ue+gqJ
dZMMitoDT5DJV8QXxSI4aeGwDNPKne3KftbqhsR3q+20EWFE5Qpok58ePbf3
4R/nWlzLlqGSheTf+mx5v1ewIJ07OAKbobjVXd2qjtRvUZ0Qep7WV2zDvCn7
Owe8S2ZwVcL572/44cbJteR3YGXXv82ml/+ty5CKlulq//jyMMpFIeR5/+0b
M74AZtE8hMtpbyQJU3frkJCGDX5ge4JsCcfm20PxiUCIbT/X6HprU1FSQHgo
BWoRTfZ1cTtOZDa1cO4I+imGNAxefVoZtFVNq28Xx6LGDMXo8dQECaPiJe5U
z42ibAQpZBAA32Gb1cPghLh0vgw0ZJIOStDAJ8KxFiFwjRYZbql8KReYpisx
Ins8WwohxP0x+0fnd2S6szm4aqIjWopr5vAPBe4hBcQmGx52bTAMphKCNzVs
w29gE4rVmo9g8sWuPvycuqCGOhWTWLTbIQawh2dIWZEvSr98Ho68ZoZV1Em4
sVM/UidnPR/02FSTYTRAukvDvnHk7dQj06qaiAjXPUX4FprnwmDVXGb7aOGk
4zIiFFAfPwnx4z8a5DRshH3djeq8Yj9WTMPIVJbXKjSoB1JGPpVXKSDQviaq
iCDLl/I72JtIvqJ0p5xcjElMNN+dC6r9X+lqM74Xq0haZCkgMuqAgKLsVBhY
I3Fv33KDzO24HUpNwqB9m7XNYQpvIU6HpF1LmtYDqZuYJ7fUtN7X+yjb4qs7
Tv+0s/c3Z2oTfFinHFIQQ0epDkg9QCLtzNEzqzlAE4mSHuczZsPGF04z8MoM
6ras/T51vb+mdtzJKACx0e7AbWJbVppPK/2AR3RzlCPwc8GYCV8iBgyGDQVD
9TKjBDSimqX9iZXYwFMcwineoU/1OimmWdBGaTkv4qamh829BPRAJ7wQcn4B
LaLWvOIsuRzSlHVTZsUQ+P/nWTsRlaBLcC/CPRZ1ak7wzkWoNlCLEqSMgw8p
A4BKTw87MVLMyyKTlFNqESkYm4HTuDxopYbaDAegLgt81HNssv6J6rgwr8Ix
TKtRKcVo56qd1v5xk5qPU0oM20lagw8Oks9cP7X4Z/oesAOfG96daMmVptk+
1mheZ/MAoaN62DnXciAOLIFm9phs8Y6P1AfV7QNAiS/T8gHK+e0FaRZ+NnYu
gtjgJrwYBjQW2j1UyJTOstSVwMkMgB1KIEngmFophUaxL4OiYx6m0V0wRrtv
E15c6NGKwU3gnfK59VZZUXL8nVtofatb0ZPscJx80Trlf/StBz158zbHpHRz
FyM32aTHpa+C7Yjkskt4OVuFeE5kKuqKhnIuR7OijdDtUXSpIVFCIhP61/ba
8waDBxf/LGiR2hmFueMfIhW/befR8DDElrGEHZnXv+G+RX7SttdYNhoOoF7M
BSER4d1CWaZOHyR7jYGdFWVD+dZtN0OW402XjKLjocGgMQTlanDGc8Bw2wic
zSZwo/r3KNoNVV50DSTaDpvmzjrJtMBGnFL2KWEWELlB03vu0Bz1SbCs903/
7ynuZvy+MgNhrH4t8L5Kq+gYQ2nRH3PC9/zVqwf7+frPkoZXvoWp00LAm7oX
SW1XPuS9+qZlmxNdnV0xCuL/YPQ/pVFwCadHl6g8UGCeMuyUj68FO0ZpJfKU
djSzlmgG9zEg0ES9qMv7z9fJlGQxUoO25bPwkHimY9E6mEGeghMSWaDoKe9G
WL7tzjutoJnE9DYJcWaCvqocYxiXTA7o9vyw7qpBvlvEhqqYSz5e2HzBm99d
UlJexgUua143oRX5eVs5eTS8fc7ZHLGPfMurCUU77nMm2jSkKTOPpZhPl0AR
IbOR2UBMiHZaeNTdAVIib08VL+fmbEodT8qn7mBT8nZ6JD3OzVoRPe6+Yc0q
AC+xn3poTAhGOyEVEqGtSTXhOrXwqYjc8hlH7TQrOFvzjGUR4g65G1khIlNI
XsSGHx7NDobCvDj45o8vLI0uHylvboqFOyWCTiQzA8e0iSa/7lqW0Aewbhqg
oaUSgCfpsxWLfF/HffxI6FKJXqfvJQAioeRHSMJ7A10+YvbR6HCOrR68zg+2
c2e3d53mflc3YIv3G114IKrjYoAoJ/PxXF1f3lEU9ZmrJuluVzSBztYYepQV
O7aK9oJY1P41DQJLZa8+nEIXXTFr30k7EVAaTbxr65x1cY7UWP4Jee+pJql3
yjwKpPQ5ktW8KuuPWqr28gmpVHNF8lGdJw2Aq1wJLXKNm6j2NcI9Ml/B5t7e
lMbnuBJk6NwVKAoQdLmpSx885U3tVaFGEOwN5iGR01sRKmugsHSS9WuNjruK
ycYG9oHvDxClUs/i+E1+mpsqo9i4E90fFWgOza38PaSFzw8FTg7mwSfbOHDK
b70dvrTUYqgsVxH9i4m5SFvBbSbGjPEbvJAYBtUGl359xYg3UvdWgsmcISaC
Ugi5jgAy9LcuwVz+/ISVcebI5R+Q8k4YrvA754P7uhD00u4Bw5l9Z73KCTYB
33Y7tUdg7fXSqYb56webnw48/Ukqi2wNmg4C8K5kiwVws7wLr+OkWv2Vl5xR
16QQZ3uWixtNwYL7ErovErZkS9f9/RQ+fsV7LhGlNwAIQtRiCEUqSBYT8d7l
Zi4Pq3S19NiSsePWqDfRWnB+8t10avI9R4+I6SBNEbcX4ciaYri0JKeuIf6w
OAT4cnBzs6AXnsWGrwruCWDPAMLYfF64ipCUVBGJccRdHW1EFAXFkn/pRsl+
3zvbJpbvJIhoscYcsuuokn4IRJKpogAdUsylo7MTfzPasHI6rp/gdEWU2rey
ttujffhYOne+xNWd72tFl03Lzz4clv+sLxSJ5/JEGtO0+m92GBvOEQbejHrB
hi079IoZrnNTrEFj4gS25c59bAyhr04pg8PVWFLLU+6b+5XjioE0fmnt12Bf
WaMeJLgGOWmxC7ci0/q0Dh/RzJ4JULSp9vr8JGPjM3TzkH7dGbCI0eT9dIba
r3a97b9UyPssAa1lQ9BYPGdNiBziKaX5DqnaBW2DWEwuz98hOi+KR3lU7yh0
WYJVHmZvt4Qdp1+a2Lkvtl912A5KeXLIz71Kd2Qrl08lwiDYnlNKqauWDTIb
ZdiEqTLTbPGlYLhzRUyVEnmMFUACuckat5Q1+KGsONS1FbexRdbxdDiaQapV
d1Ya76p91Ij8kLEwuzlI7nyGyCAPOYfNFXjuIo7CEBYpuxEMsAYbnAAXKDXA
gMnEuuk8eNz9QDBFLj+0SO37UygvKzTGYS3qTgJDucg36i5R1+k+2PUv6If7
X6h+OqsiK27jtQel1Ow95WUFcDRFadEjMDAzqCzsEo7xfxXH46W1pfeU4kDT
rjvjgZi3mYhNVTmSS4U/F/nSlz+/T2jny5s/6+85r+3FrxQrKNCycY6dPVjU
5Squ1xbMf20KXc3uBS6UPhA9Z480SxOjoctzZHFok9LuNcfoG9wvQJHOhlsY
v0Y2b14fAqDN//AEnYcbpFoOvL2lgyLD0MJ6Kena7kUrlp+bKGvkfYtbqEZB
8aZrs5hhKeAJuHKeVU/2BEmP5RjRYMNx30WjdPRwPYQOjqGHKwbWzLpDuWof
PYyxJZdedkZqE8a60SXDEe+ugFLMk7nAswQQKPhQO+9mH+kHEQtZQeINRZDQ
llNDdJCNaz89jZ8FDJGOpv73D+hCw8jHOO4//uQlgU0pSBxdZwmkS3H1sjQi
Hkz/wZ8Hoqt8bdDp3VhIuMcyjJ1aDDuO77Cht+sjjGZxZa3HeLySZfEqsOP5
AA/YsxYowASSZImgsPd0le4WVyfLpixdzn1N9P4cEBlXTlnVnBkeod1qGHAK
tRm9J/6y4uCGk/H2Ca/1A7DOjlQGAl06zLGLBW6BMcsddI9GA5Ls4AWBRfVV
jpQPPymrhDWA/3XfBLZPIqOY2p8W8qvrT5WL/zAZHU0wTrzfsEE/uBcLXYsf
hF5rtnVIamMBlHe+Nrv7VwYTrnzpFC2vhVNffmWq/bsULCu/CqNWYs1LYMA0
RSBcDXz8LSZINL7swvecs34QKR56zO50YEctXvOd4fSnxQWo/2HKvMAVter5
MpNGfGaPN7kLAc7pFavTlbNakm1UJj3XEcLyvW9kfIKkF+kDzUgomuaAn1PG
Xcc41YGDZ69TD3sfVH/FYcMzlCVrdkZIQ5BGHg6FuyA8iBWS42Y8w+WaP16E
/jVAKFPdueWjdxD2TWXdjxKpuwfyXhABrUqmoM9LMuNbkhjP5bxkAUu4Gigu
8KPqkwFZxQQyRB6Oev09+NBmK+oH1PoSqBrSog4oCJ+AyXgv+SrWbB0VYeJ3
iwJJBd+qilVDNTsJu6lUL+X3HuSljN66Qc2+xFl5Y29WqfEKjlP6MfKfQwEg
hCp+bdQRk0i7+qmnfbU7nh+Hq7zShhtwZdwe9l5BQscNlqmnDGpgCZcz5TIV
FpxiUIdG+n85yznX1f8qipK70NFkjXkxoRXQUZZ6g2WXwllOsSxERBbKNPBP
dUatto8jfvmL3Rm3OAwVHvomHSuRWJ+5fPTyAlrZ5emKk99qult1LR145EyR
NTan/MfL+rB/FqZYSnvihM7WfA1NuhjrHwtVZvMV9MhL6uEjpucrH5G4pAFQ
g9Y1T6DWF23Cmzn/JSeBnQWc9BasgTkKiHGW0gYMCMA0+NsVk+i3j39q6YsW
vaE1eomrBLhqSLZKK8IthDo2FXBuyF/lYszEqGE4pwjhIhHGxn54q62ngZxO
7TUIZhqbjayWqO7c3QG2vgpXvr8C6VRs5IArhSjB4+4l9njKfPi8zcIf9uml
h3CqdKOmN/WwcrH/Az4CJ51FbYh8XYt6bE2Ni/IG+LQ7T/jzYC3U/RMyU0GV
pN7FADMatZ/ePeQirIha6/ZhDL93PLLAzPbaoyGlb/xHpcfAd0A5LbQkM99P
sPaTzCwh4vkBG6i7AP/1bnrGRaUCLMONYIPgM/BDsBkSOh6HKxXsSHeNg4vy
ttP9oHRM8UTmFuhOdf2YceP2r5nszVabtq+egNU+yLBptNpe66C/E+gPAJ4h
IDhrPO0CbSdwLV7hRgmxsaJjCMrDq120hbSwNw4K5T6qDgvjz+HYujnjfcn7
ShEOOzyUCDXD7qEe3rSN9s0evCqkv9k1U2Ahhz3jRWlwMb06NRhVpNeW6k/4
dv85F72uHHIIyC1XONVSRX6xIL0/dDOueqaPAuuVQI6yr5zVL8SkCAssEtDb
vjb++Se2+o/Te4ZRu17loN+GEb2XkA1JIWEptD6Lr9YEyaYPkG5fjFI5d82y
85aiGT7RLA9HV8ux6WbBaH1xrowUptjkhH0vQSS7TWmXiAI8hf84VOxnjwN1
mzI8oVdmHhqY23L7XShunU7PVuPGeWC8Z/g+dHjShXN3o9z7OBDK+Is9f484
ceaLqno97LyZ6gH9K3QuLiWtla6p7VbfrJY+/PWgSwH0JjlLmsuQlkaMPzWe
85e33KV2DlXIsZPrwRr7AqyCMkfmn1775j2IGBWtp4nX55M1SvEX+kuS3o6i
WbIgX07xXdKQ2UFatLQxuTB1td86FAPyaPf2nheCxmcjds52IGIhnYwSR0cq
A5dwxgjBTQdepi/aqKxBFxVohTArVBL/FIIoWMxNcaF7fUIFv0amtVS6YSD1
JOnOjK52X+JhplH5r6XFcT8t4a139EsXIAwxArypYt/2Siy0JX88I5/AcFbL
L44sfXZ0ECvAzzsrKxKBpyurWSaKnE+uh11WqB24NcyAipi99KxrhyWxGZgO
YYMVoVJpE3TpbpDjTSl/xBl7pbePf7SdSTUKkEqwc/VZ9uFewX7M1Sfn8c2V
RLFOhnm88vZ6S0/UvWjjBlEqvxJguy0JVZO2Nj1UYWoK5S9AiErsnSFrAfAU
g/MfmT5T6nWTjwxngeZ3GyBZi4RI7bR83S3Y5b5XC8C+mO6kAoo9W5FD+rAb
G52vL4wyP2oAWdoPHXo8z92b89UUIU1UN3bkRXEBfi8xv7RoI1AxxbEpUxR2
DV8/uhb58+8fRkg40V7/Gk3sWCVmbsoyuwYaMWgFQIR5PDm/Yp0L6r9Sa73/
jetpPgMQPWr6+WS9tV8egb9mmIUw5VHqXTqaUbpexeo8dnLTj+Ji6bRkagQZ
hko/Lu54Nvv4KDIZ915g77tZ02wCc0+p13Br7E83riNG3v403uyNzWVd2oj0
VHDA5PtShRn0BmlP7wsxBf/wt8faINB9EYW+ZkKgxIXEPaAUMS7wbfbkbKer
MxUkGAySy2A3RJJEWvF92bnNMzRbV47Wg0AqVo6F8CPiQTJTBzJDS0KbtxoM
jgOS50B17rJZijqbdZQVlybOUe1Y/MPSYLI815ENJ+k3/HRpcOHhUWeWsM23
L3tlAFiFvSHh3jp/2/gHolNjsPZD6HfCvU2k/t9H5BoTco0J6OTaLvN93rZT
x1pCfEJhXUAfPU1N6C+aKsS3GcraruPIZ3g0Qd6fm2ZQM/IIOUOe0g1s4hq/
NgdbJ8YyF4c04jqAYyCM9ZvcksB5RR1Dz/keHK09wkVLQMcXUeZ1KAJUy/CU
XubuJHP93V7ypVLkD9YAPqrU/rlmhp68+OWjOaU8YPc6iWZ7tAtfICN5H/e4
Qm0epSlhaw4VHtPWaBcPhmXjFhaAokdgAONcsCENYYKXOrhavYPw+z5q+K5J
M8YQQVCswSuxhDCvfddSGJaF6c6zxLdN8bShJ8hLEtsKB4yziq/VV14YR9tO
PnwGvMI5RTF228zoHGyLDLTsNkOJmUqC9yhn8DuJynk57jMYWxHxtCPq+Sx0
AO0+A3/IY5NUjmr+43jkoLKSIE5XB6pfuc2lVylMjL051G49Te9fJwAZdA3y
QcXcOr8P6STckPBEGoRD78imb7LhM2xvMnpZ3RvXbJPjvVT86So0FsI/lyNq
g9QPpNhpDgYi8cuz0DdUtxynT94sV5qX2hkfRd38DeKRf9ins175LOIwfSFc
RTrK75wfi5Ln2mDzzYsLL+aSlcgiNHssO+LVosBIqVWvYDnkftrChtbuWcjs
thpzHtdtRAgaTmZrgmbQYKju8Kn/b2qTawQEtpVvg4QmIVfzMN9s1oN7ToTN
iY/JVJeCE/rif1AetWV5aFBhzVD5BxvyQzNBe8KdBbcuraSe+dyMAH8zMv8d
C2+E1wT2DfcwJ+TR5YNA5dVY0nnKTH2IgyErHS/6Q4rQZD89nyXYdrSjVeSY
o4PEf3GBmNKOOOSbRDMWaIHy2KXcN209XxXiLHJNe7xTDuqQSFA4BB4jPG3+
JE1Gq5WuovH45zU5eOaoakGTdbcWMTqg/LyGzg45xdLiI2zz2Pu4y1PyVvze
7E5PMktXOTtehi/2pF9sz6t+z8f9pZl19mzH/D1akIkr8mORi3puE+CxUmQS
6g97tmvc+le6I2/yTYY4SlHBX3apHYWX1opKgZPRsdiwNAXKJ94WT13lPmrE
neMZRfqDjvc65HDsSjxQyhApno4pwNFnKz8gVrSG+cMfoG3xMtXYvoJtgGaX
CSOawxIQhRIGCS2H5/VZ8KAwMQt1b1INgTiMijg7Kq10WqSezAcfS1YN5Snl
e5TLtGRna7xXLsN02nbGP8B0WD4BvUDC2ud00MOq+D2/KROGSRpACf3H3L9J
oaHHRKyKJVrgs6YACCjy++lyDEJpAIkjPdjbp0fbBggGdwWu5QqIA+7jgcWJ
4r+Y0a2bsWFZRpG2YDEIy16/PLChJKhpaHsw7hp1hMJt2miIsQAjGj0oLCGj
0D2hs0i9K0lht49s8EdGtWar7A81HOncX0IR5MXJF9AE+SOClwOpm21I+WxM
MtcPSiosUIEcmshMDqI1Mt9kuK4yKcl+g3JEbs7qmzB18nfxnDsiHlmd76Xb
/33fl3E0aeRAHzAXZ8dqlR3DqwkO2Hd42SFmg0MloNHsg6EEcUgkO+eD6gGA
+bZ1cGDvIIZDKt0QL6Rlnwjab+iPZfXJxZtAQiGXbc1N3dRBUxAS2u5+RMFu
xKBsfuP4tl8TDjtwWuPpK8OgYOPgm/fZ/sqW0vFZSrMAd0HQsjLJC0EwVo/m
PxwBCtQeUaSl6DLeNSL+6aGDVPfYjONoaqWKp9vT75mMc3tqLromrQwDdjME
kmsbyq7IZ8cB09TCR3Iz77u6KyJkAqrcL/laDMRoTIODH/mhDhrol943euvT
nXZMUNUaF3/gYHxM+9QEODC7gwnRmCh5oiDoesaEsLuirlpwlghH6nsazX2Z
4p76bK8gIwTI2O88/ZJ35begQBMardNrX0afoPhJEuRVUNyDnrq0u3lTtd7I
kIcNG4lnbkQRiJzAc3GwfNW8X/gcMStnLJHfrUxfi618KHhuEzLDBpG2wuY6
T+Ctpk/tK9E7t9UkpoScnWZ/0s8UdXzbE8/RqAJ84vZHNZvJvLh7wfsxp4HZ
QKDlVdCMIKZXo2rr74cG8NVEG4C3LjZW3LHtzLpk1+o22ksYSxsyTxHo+rlX
gPOlNSQOydNZlxovuxjqwfoFBeB+EUC/k0B9H754ELZB8ncP09mzviDugdjJ
n7SRzKEbldJYj8BbNweRaGkrgS3J+tnbKW+fGtTmi471ukDfn3WzsdFdcM0D
tiu4i0VOn0ytrmgVZbCM42dIlioZiZWpoQuTE7kyv09lwr1g7vKHcidPuuLD
jrW9JlVD2dwbp0vBn123r7rgv70D8xalbrJ/5bZ8MH4Qxb3eJUKAGUxKfck4
2nY6YaCmv3Knf4uDKWHRMvYUNf5O6pQiZyF9q0IP9UmGEmPhyJHAGy9AUow8
JaqtsO9ioUwtA9Hhr5/Cujff+hi32cGY7ODy8kQ6YPrNmmK2zBlg8iemjvz1
YJPiNdkew0CSPHd9z5MybniLnU0xqTpBCqBydYK/oZSMAYGVLESx+8+f71nh
YdmKrf4E8EJo5ksyFt3yP501n/pEdF0tO2RBYM8lRYGdAgsiFVZG/c+qpW8P
0nCxGaImru9+YNLs2xhF2PBljCfN490VZZtd4BJawAaZKYuDfuUaNwGnBkvL
SvAddRme99/U/AAeEOW62hNP1qeE7HOKXh/haxfH71Q55S3Sb3bhzCl9TI3E
eWWRmnYOBpNQmA9nWSo+Sx5/1Iyg1Nk/muFwdluKdJZvpDZilO3ptc/mVO6k
6/5wu1wZt+rnCa/bF5U8IBrX98uZLRevjjtgWWr1f8HNlgB/8GW/c3Q2rVWv
D/51lfVoB72xzdSMjBbsEYb+FEX0zne4NjEtKGr+fTl2ytMVp0fB4R+bttYx
uXNkoRZUXC4Uv+dNqgmnORQ9jfUd0/GMkxPC2pH0k8Gyo2/e3ZCugafyr/a6
wcDO7eaVsfpUnMiif8gd58slSRrxUPBMMiqboChSHQUVRb+UHJFOeUivIV1u
sWNCX7ggqviuNH+0bf8460kbfvetwWQi2NZryaIi0uhkWm4LVutD5DnRnCCE
RlQtMvzOe2CVFmdIgTa+QLoHlNOXKXwAfyrcPeAG0ABcZgRX+HrXsEe3Vn3i
lm5gPj8mkIOaquTCf+pPxMe3n5/bxrFePX5bFHZuq62+irYCyks4ERVZKXiZ
GKGeb7U2pQjcj7627hp92YG1mzgVIkapRAV9a5OGc8hxr6A/eB2Av69Sb1V3
OObQGasniQdmW9GIaqUsCFPvYKT3qzqsYH8m5OlvbWHdK83uzzLKoNWzNfJL
amRWgAz7qMFyuDpIWuTytPGB6Bf6ZxeZTB7Ft9sKUTRhniiH0ZY72ZEJq9y8
wf7Vuwa4JcJuaemA8C897dsieeNQqLKpjPOXf909xE3oDfynmgZYviVVRNAm
hJEl0Hr8NilARykKm2mSd9UhNv94JWbyCxuuZC5v3zVXpZjhvQYz4bFJtX5f
s5YLbD3uexdawy3tWjpulQHoIEOW8xLMvpHp2ad1vNh7+5GyCi/+bvKDULdd
Sdn6oVu6Qc2/wvPqSFErOe1+pGnLwzunJ2iGZhnGk3PPUADalkyNrfFASdw7
t5MateDgHFSVGuN+dT1neZBCa72gQyPQTIjVqYE2UUYbb9ZJeG/IP0RNb5kk
8uiQgqR0Nux8Qg7miOkt5FKaabsh5/lEwVKBg0dVMBJ8pUCavVVXz5XKYhAO
iQWPRr/bXL3qCUKWigcXcHNsWP13VkPh8+6k+FPFzWMp8z2QJ30Ot6oPAMHg
jAUPAIgFLvHi3T78Lo5x/S7l8oMUNSVu76FK7xMd2A9OQCfhZpMCMLX+uFxi
xJzC+uylPAtDpqGlPd6ZXDHvmgZ1TMxhzHX6x6QSlQIQ2wL7bb5N4Fpj4da+
zAMU5DYGJwGop5Mwp8ZH+UwJEGsnyexpZ/Erc0LBiomjeD7hDRMbRg9jEoGo
4v+h8JQQGyUXOm4FjZu86zRPDexvKm0Jgx64JDFVh5xdBS3r/ySP52+gOD76
SjvMvvRpp/vTaxA/N0847//79jIsa1TXoEM+5LdSDFzsv+S7buFW43sIpVfy
PesAkQ4oxmS4o2wVC4zzxR9NJ/N/+x5Nks+Mhzf0nURD+HPL/bIX8F7XfuNk
3lTDwOzgQ1NAAecqu3fldOBTSH68zHQrn8iBzDERaQjKmF7hS1ThAjO4jSoQ
m2tWArIzuUSLo8xGXsvz56XgTiERE1m5XRB1H34OZtMlQfGWyhcEW7f8jQ9n
SYPh9pJ1cwsDpQ28YYngQsS1NNXz37UFOFGQUuqiOs/FEFOL4+5gA3LoUPjo
fAMj0ipxNg5UNQWo6YHpnpowQ1xFCY07j8zw2d95ZDvo6/C2GNpIRd/vm6zb
C/5zL7mduHh7r9LNwrPCRnc/YeJnF9Buic2KQiCm1dFWLb9TZy+MWM98miDa
jff4/rGHnlGitbchK3bJbS6w14H8LNLKv5+94zGujUvT/VRkZuaXO+CoVjmL
k6UxH5AixPpj+mbLAeE3b76px1NtVLQbKOQxmyAMsv3wf5JXo+ExkXlv/acu
aLCH7yfFAlE6B4M0GvoIOyw7KiPTzrfLnknmEWJVQNH3EFBDmmhvlgLC5Q4B
RdPghUU78Jw27wdhaNrPexpeQW3SbQbaWxtNRSmbRmbsaSLCstiptTIxESkC
XWRHpoJsXZ/unCptAmjuEjRJwObQf9xraekMofZQKw00f7MymTpuw9QS1qQ1
ZxJglKEhdfIQl+OeF+u8KhG47mhLcpi4RjMauHinJBJjivMaAJ44s5y8Jy3S
GFIQZRLpIfgHxIsCbRzpe2Mau8bIziuf9wuVv1eHAdkkyrH3zzZhMFZ7W/xQ
TGdJkpzFLM8k4iEke7M0wu4zHWdoZoKbx+3PF5L7FSTrO9pPrbPB0WnaDjbH
TtpUYyojZiRWl51GtQYoguESy9BJgcUZzSMHs2hvQ8Smu+/QeStTYbtrsRsu
lmem8G/Z8whSNBL5dFZ3VBgBvwYxlP5TvDMZrNBSFZD2jcq4/QCtC27sSYhA
1QwK14xTqO+yMRGWJFqTbtk8vHnpfI1OM8kiwj4moBCwfBB2gz+fIoDTMIln
FiDHq9RnXJGGx2HvJgrb0H3IWsTTfe/0XstG8/Ai2Fy9kYremVAmllJ05ikW
L0Xb3PlxWYabKN9ocyP7toJtx9iYbfGbR9BrPrAzair/Bf+n/6OmhNbJokb5
NSaoybmZulFsPt69k9D8RdjVuQv3vYZGgGVYDId7UGutt4A5QpEYdkuMMV1b
dULxtW2JGc+3fnxxU5sQ8gIDhnoEmFghKOWN03r8e0JHpynssGF4zxBkEatN
yG5YhCQ/FnfsWjRzOJbkUWjSPFwVO5xwFQbgGOpgALoBo1IMrNbhGr9tfap2
07txeJZU2CfTU6UeLd0TuHQHdsB0ggWG2hAQ5iA43xF78DiZBEMcqwONezXY
Y5lKEZYfPLE9nz8DZWC/fxTm7S6/6EQjLQwfEYAVgXgvGc9OIwJFfSarS4vL
xhlZ1yigFjQp8uaPnwHeeNy+S0hIryFmi+Psqk1Eex+UFBwZs0oSWHnq8xwi
XOvg1D8jV5dnzpcs0sNM8Og/IvH3MdA6USIw3bIfTagQSsNdpcEAXKFEcKYj
137yPBdEjaj1UuIoOg0TGUbO42SJ17OIn4x86NTTYQOsbErs8QbVdeErl6f2
dSbVc3wDcmvs95BS0FkDVHapmJCS2KTU+8Xyt9Df7NLpK3ECQJvTfjQ5Gq6V
UlfEq5RnhG/+6Im5jjNeIOJcLTTtWi38kmV4jp/x3RwpGccbIjjNihx6kyol
dxBoQ3TzwyAxzvw2HYfYDRVOwaGNmnB7MpPv0M8abI1QJrjo3nud9PRc8e3m
YDYImkPyhci6ZaAr1sUONK4fsBclnfQ4ECazI2S+nZ9Deu0K7x0as3x8r6dO
iVDniwcSWhilua8B8v1uX4Bde7XgbDf3tksYP23ZICEqmX55mbbblYcsG4Og
DT5U92bN78ITl3tBF+P+AnL3JMGo/9A6FIPdhTTnt/Ka15oSoOJXY00Z6Lkq
ywXO59Micd09cuRoaRwkyRAGd8NbfqQGpmiyFOacH474K+W529noYN4SVHBU
F2a68zKfZT1KVRClvBspW4U9vMKbS74+rLJ7u+XD//fK6u8kW1qSyoeEw+z4
ryiA50yPnWVRPT+fdHRaCnU48/awZ/D30FZKi3UDynOYfCWPRuN1SxpDURYJ
lDyNUVhbCcULCygHRtyEh9E2dzgKAia73kCMgqU70q5MT+mGKTG8Qrwhhe3D
TP7docMZvJEw3ExXqrXh00H+MlzzJvVAEQw2jrr9LkjE1Nnv9rxirtVORUbv
KVpPVeAuUdTRGdHMDehNytt/Vv0pltry0UGsIM4pBgsg4G5rMow8LBrWbzR3
6O+x608WMMKBIM9d/kvm1GOiYAJxuAB0VxQvlG+6JGiTWZIrTe+ZetRCy74e
6tBT+EtavkdMNhkNpc7JlAU7MwKP8RMg/2PwXuVhshX8gCB0oE/pr+fzexov
/Q9QbfxCGXlvgMpMZ6lHZXZsRs1e8S8fhLCJ3NM+Dip1CYejUIdHNnW2Af0P
8Yq3imazzdPOon2xfYU5tPk1g9LgXYZsMew4RuobTSv/lCgs7jSYWeLEVfNm
AbbQ45oWpb6lMGv5CsF2EHLE9t/Wx2gT7PZ+XkltRzi8oKv2Gi5hCDoTE0mG
Eor8TYeFjEA78lAGTNrUbnflNdZKAoheTlwHgTq9eLkbwPwQ4t3rtOdr9aYO
VzdtBoF6d0HAEiqnT/U+7ji2sggpItLagyjcgJxm/O7MQUUJlUBPVn5Jzqbo
L1/82DhYubqWOysyb9iZs6lhRfzaiQejU6im4Zd+4vccMjO5kobtFpucsUQo
993vUiUGAL6HClPY+7JIgsb4F1wd16bVOheG2pQ4JHrRjFim6Fw5Ug4/Fv7a
01DOxUD0DAyNPXcT/RdbHEIKnHjm7coRx+RA3nxwwPUICSRL0xC8RDg3+NWn
2256T14tHg8ziSqk/8T+s0PfcGkbA5xLOv0tzI0mN7FQ75f/vLRKM+k3dYlZ
REjZWmrqM5Z4CPU2P5iLnFm7UN+DKbmqymXZ5X9jZVWagtcOBP1hSF2Ko42t
jHmgvoxGj0m0XCzNV4PwxHlAChkybMDfUG1vnby1VfLod/zmsmB7On/kyoIk
B2AiWeedyfmGje7MFQBW1wBSPl1K5YMyv31SFldBKC9vwUZi/5e1fcKWtf9I
qol1U244LvKyfRDhLmc9cuXgcHOwfNGrVvdux1HiK+MNIgPb79fV1+VXmm3p
iM2CLee3t+XruUriXqWx7rbicU1P6o0pIaXXJcv+SEeW1yimR/nAJCC8Mwsr
0vwSRIW7RRkr5FFwEwDpuYE8PxSXfn2tXlgXzCLlK4aEAUnT9hWMaCo29J+W
byvLI8K7UBXMUPBb5cZ5OoQNfNb5mA/8C4x6WLVh1Sx+aMqxUSDnaz6dPSq5
JG4gS65NYy1HHM0vp8txXF9/YTxX3I7lD1MTuEkcuBptdSiw3j988vXOyD2X
c1cZAleMsgcffSxf9kurEgtwDDZGaWBUKZ5ErjV1MDPD/2cdpecoKkbC2TKA
nGBP7ICA1VsiMQjB4JYWjDQKchDJhnKxQksF/ZwOTLdHjPCZ2drU2ek6P0yC
jMBO4mhhNSqABjHYKoMZ5Qw8rlq629IcG/5oUCQ9UbQBqxQ2pLQrSz/yGS6m
4IELy/jY9KRx0raqfHGOYILeBaSF+uhMRB+NyYfgejKNmTBDBJVQoZU/H8uZ
e6knlxBeyhK+TO40f2OxVmLrZJMcLI3QrJHXl4NynjymO6NmtA2z+i8weqgn
zC5PVTDf9xU+xI4TMcjTA4Ppp86lD5fVxEw7VtWTgxOs90oqUOn195Sr+R2c
7fC5mZL2IeUTAR/jKWWepcjIuKw7QmjhPQTYhYV2CZOGyMCRRxt6esRhAYy0
VE7e8yncmbcQw56xmXyf8S/DfggZNRsRSFt0RmwktoRFtT9oUxEs+ZFrU6rd
jVCEMs1V9bGM9Au+0tJWNKLfO5Ul2ixMyP4+J4afqcfIuz2Lx/2PJb7y9Fur
i3b08UbpWX+kMisy0vhSCN++8rBCCHE3kHocgs7MRIr1v8Jcv2mL9rQFLyAf
qb9GH7w1M/AIYKEzETQ+12I0oJPX4qzJml8RaC5+p8G9kEVL26RHKLCay7YV
L2fsG4zX3j6QN1OSrXjqw19F0ZWMD0nRQ9e36JwWiuYVB+ui25YJ89Ya2hTG
gnQ28v3fJz3EdbFcoCm6Bdyl+Q4APKPNgdZGhTZniJfkER06dCSvGuCQ5L76
9uaBrsDuFC53gAY3OlvmT0ptZRucp60qRyIJUo/BktWGD7btXU3XZAHxmO0s
JbowkOgOB10Os+U2U0WOXh5RrwjVrNnC96/3o8PKlTeDn0zpPuUgXsIZ5Qzx
JhxVN5sNEkX+d3LrxBtVj43N6eAsvpbjxpgB022lHmnX9d8FP1D7SnfcHuFi
0x45F2qyuOVQXCs1zxtjTNWRKK6TS6MqITlf4XHVBQXDEUwFNXNPo1r9zy7x
/Ar+twXk1aZxCacfiIVCxuEO9FpNMqk3bMg+Ng8pxF0udUJw4LU75sn2ZC54
iLSuzZlkw4K9Etfnn749VNG0gDAFgiuz2cbfGT+Z8NqwBUr8MNOnuIV45V5t
ybjiGl4/qnMtWkaD+ZAIOaDctzHOcgDspr9/KbyATYws4E9UetC/qXpvEhCt
H6wdfw5uaTEzcB0M1+XqsRKg/PalDkC6A2Sz1x0nurd85pePQlawfvSUZ383
a70zKKtOFleH6B6kc89FsRCsYazPeNfucfWGvpLWsRdtu+VFfbi3iNbpZ7Tr
sOwuDt8haTa8PffV9cGAM+vLIHQAk0SUnOQenf71O7knRD7rRqX7F1jrzoeK
k2i+gEHjGxb5Ihm1yluueId7o28MPUTDZni7SXhkfidHOpspTWJIglVHIKU3
JWBX1TdnXJIc5JiUOtTqv2L/ryXTu6ta8FRvZD0Lju3jekIyqorTqIqwIwSN
SMCNzai+RMnK7Ru6zuRA/ru3+/85jAfsBr8NVEFWONj6fuCWC0kFlp6g0Tml
b0+KQctVORwalxEfRTxFVzIUfmoKoRJ3SaXapTfUdJ4zDmV38wLNAIJ49VNz
lMdAQld9YpZl09eo01eOS+Jbn1Fo1Z7kmBV8bm6LN0HLKDmF845GKFQnKecJ
v4Ccrh/kHO58G9iBTDO+z/8rbc5d84SagqWuLInlXmcXTo2fuKIbtLfhekGu
w0wbaL0U2OH0huFCOKmuujlvFVf0ATjyc8QiTzHTzQPvnZmjW34uc1CL9dHr
ufMzzbk87T9KWR5Vm8fJ0YChiI996a0X3KEkHTUwkfOXt/n46Au2sSfaqQZS
1kZwRwRdHp5XWqSg4C0JU5ZUmwF4CbOjNNd+BBaJana0QNPkjg7iIRSJFWD5
GYjv9M1NEojCFx/4RxEmy5/GKndU2YIcH0mxTgNXHpvwXhg8N66IE+63e0/k
Jln1NYhue/zkgcCKOp9twFMjHjO/j60lygilMh0wOBWXGA7Gm8j+dX0ZANMe
OLlQXGnBsvBLdubQjewVh6fNlc2/TeBWvbUVECMtEO2wLWtqMkVc3LevjxMS
8jbKxqmRnkuJXWhwcBdmEY0G+VqAGKpAev1UnaCU4Q+SMyLwE8d/u/QHkFdo
tAeWY4GQQVHSKDcrhYRngd9b4z33rN2tcG+whjLkhc9BJkDyGj4oriVaPVib
loRYiwYyz0y7Hm7J6vKJLKcdt81TOaZGgTpEdUIPf2uq9r4BeFTJp1N27/zB
8ASrlyx1Pzn+F7K+W99XxiWwfmifXA3ENKfuspG2pjthU0gkVsYah4zj9euY
yviS2/rfi+5ak1fVngCTmUnfIIrZcCo8WcfuSKEUYMQG2L3lWrNO7ToG6MjI
pq1p4YdxmgGnu6mo4/W9Ya8/AhyhuHC65rA9kiw3loXlC++zXuc3yY5s86eo
OD/Js/G8CGZhou/6PDbhddan3ZphOb2KR1djcRs9pql+PUXhJvfhOrjVeVTg
3tJeQJkNgIocSEkwV/nW61OpMS0RgYGlKd2HykXiVf4FI3qd9xBurcw7uArs
F7V7ppUEtq0sFilYhhZY4CEZefM0ueZMJ1tKiu19iyeKx8e9Gxz1crMO4Vx/
YjgzHyOoQ5JIG+iMV6hMvgSfBsfa+d8z2KnoJCpTQX+VxAQIieoGk4ix9hBE
3PTI82YxMcW1NNakFJndAa69ChcmvI/vIvnhukrERXSA/VtiLgVmphT8hxp7
CahBONiWCTX2B1x4NA6SfPhxG1U1lFAQHYHDwhcxBTti0zTPKAh2iiaaHdCZ
31xQ1YHI29VtxD0F0220/JaLX8kHCNOzICd0+/Z4d0/tP1Ef84h35VV9UvQu
IkiIxDvQzGFUPyKnBCC3ACtLhUFNawQTfeXQlh8jE4Njs2un0tclqgDjmEtU
/rqpB4aCGRY9Us691wNmHZiE/4/YADuusEi1ryf14o9K8wcl43be5aUvfs/P
ahDIHARlyUJjIzzF5TPGiVze++Fv5tC0GJo3LI4VZg0Ew9KEbo8sJDY+Lh62
UvEbhuIW6xci0X6xPpfNXhg7TZfy3SNHMnxTcApmCFi2NcGclN7GCs+pPSMj
+YXNL8r2Zq1UJV1j8pXmqfPn+qmX0LYujchhhDVfEnt9ZMaht+rZjkmXPKU5
m0xtx88WodFdrZAnaLNLTa8KEZxSa4kQneHpXwGe0qpeZrKluDKsFittBRIU
KcMjtZ7WYDPavyH7ysqqdb+0L9AlZYTT2xPoriYfTR+iuabBk2Yoh3xjyWc/
xTf0m+cMERAXjtCGu2DHGl2SYk7Z5qxlD+jNRCdtC5be1dcuOABLOMnKtvxp
svglfFgJGs7Wk3iaccO1RfuHeFQDhZIZ3NKA4HW2MVHX0JuWKfsYEzwxwnBw
sVtsEivTTYl2xFcPiOI3IDA3v/OpDbwt9a4u9ASuyryXdtSojJssaE0wzTsb
K/wJi2QbUq9vUpn3SpcRhxX/4GlJJ888F9OwKR6bJ6iq2OGoIFj2WvRO+y3H
abDQP4q4iHkefMz7u59AMIBBKHFdgOhBp17kQiUEToDsReR63l+2SRV5whJt
vwYsyPMdZxs3uZVduVg1ZuDYp4S9lFe4LabInQgKXr6BcVYmiZBzVh3b7KjA
TLB+Y4m5iarppEv0pC7SIA3pARSkZ1icbqODmw1gf9OrS59w7OIg2rPcdVwK
7Vi0yxKCXxKjHYWwOGFSL1KLZ/Da5wg0VMuLbPe1xv22zQdljWTyShEu5OAK
BVPHTN+EzZc3CAFc2pYymESdr9DjEy6CTE5VLpdU7YdjyLeRdAbuRA6a2Zyk
3KJCpkHRixAfe4eBAdBIvXugks5vvTfq+l1+xWgDKIoNEVf1pMk/0rIJd2TS
hP8aTpFQNzhL/2wQgyHw2vJi4u2WYEYAlz8TOAGuoSxJI9QfQ7BQACBN5aI9
kgQ814h7Uge+3R305uD9Qmy9gDWdqkX+Y4NCWbx/4SgnaWVJd82v7+xfPRKu
R+xGc2JhIfMp7itHC+gwNWNo37ttLA9DL/ZD1mZZkjMCo675hLqgYSXdOFp1
WGqlK5+iwykCFOVB/zg9wrThtXk7WGbF4dbdNA1MyGtTyVetV7zJmShW9oh4
i3Z7I+cJnZzt/T/6nldF9gkXW3jaqFwqJoMsvqkExjKpRpHkvismH/Tdeg+Y
Rrl7DN3cgEGrB/F5ialZfhmK7IZ8cfLBFxgffkz7I0EKivrcVnuxkkonViK9
mmlKcLpTA6uu7sxN3r+6jpMMVCmOUIF3b9TX118KcuPC4OOBbkkRsWG/DFMf
5mq31eU0lzDUojkGWKmFbvoJZyUV6eRy+mDZuv0cQpUbfS40lFmDUiiKiPHt
9ZLdrNqYvXTwYLyyxymhqfA3I1PPsdhu45T6Vi8rHbg2YPh4kz61zKq+QHIV
q+2HOepyjPfIZX9nd9oZ6d+EAp4HuoZQ76aPqwu9WhXxzSERrk3741VrEw4m
OXfQJgumVPv6hrHA6sNabhz/+OyGc7KVedn45dF69ZwfZUMsWGeTz8wT8bB4
5Ua4csa8N/kl1jf3aNgQPA6RaUjpLV4/WwXQKO4NmbzgEKI1J60ESp863OKC
RmS29rmaiOgoqzmzfMWJBOaN6ato4AjKRctCgECcSLyC715rVUaTOkkjcr+E
gvQTv9PBE/X7Uf9iOdgwzKmLLllaBz2u0ihPAsjwONfonBPr7POZ06dDG5ZU
mR9S9cCVEnpcEhDhvAEQg8EMxWJ5c4cRG8dRDL/Pl3DJSiMbQKdOVNuJX1AJ
rAP6nGCileYMaCr2zDcvbONIXwWnvopO3agBAsoMbanmEHeQ0f21cdl0KDiu
0H9Ut7ncsqNGwneyKBhS3DJJ4QW8gYHkPWC1mzK958Gq7C4UHwLCAhKHA0tU
HQ+CQiO6M2OZpWIlK/xQdHUadLEBolBq1s5XrLto2jAhXBW+JH0JUhnj/woM
HaR4X/C/Z0J0R+9gWZtetNSsqD2O9P5n3oBzooWJJN0B8I8QGYJbOe1tyqDr
VejgHECAKs0PBWx6NaUBiV0CvmrisSCk8ZGZ9Zk/4tr/OBo/YHMAGiOF8QS2
BzSFwwyYL0NhvbjB04t9C265UQU97UBy5pa1qknrP13n9YRXRrU+B0veSI33
9+cY/Uf1gLyW/lroZrtjO+K8iohK+3v6qDJtYZGM63CYlQw4GhffB44NJd45
Qzhgo+K1jkuU4DLPBojLhaNTqDMgID7FSnFzN+1GgExc6Z1LAeji08WVpaPF
e4UV0geU2mmy34kSBsy6LajMD17uhXPSwNZywdT0pCt598Jc4TMwvXBQOH1A
ev+IZnHgxn7XcDhsWYAd7PKLsqQTwNF+TMgURZ/4ubZr9+3ZsYd5p1bbHUjj
8/v+NtXZfGh37CYgUHSdhzPVoFS9vBtKwUMYAvot5PRNJO97Z9ruGVF+jOwN
UgQOIXqVOMoDdMyb6fWNTK5sUU2aft6veuRpsCpQQw8zw+zdfU/5NN4Y5SpW
iUca3rOxvNt5V+JILWRnaH6JK/1BA+pyNojZ20f8G60WKJob7lSE1gwsBCaI
eki/XDY+7l+bIeFIVAWwiRaZQFk1WVubuYFE5nXJoRhkLqocVDKg8p/P6KHx
P6DKIyx+x9HfursBqddUDfSdu2lTCyc5tRt2ObKdnhNvFToPgt9h1fLjiq+P
QJn19k/w28AkznBG3uQor7QxspzeRU0FpmonVbbgWMI4M9KxTsFIxZgXLRe9
kLSpV87ORjE3F+fb/MPMktfpdmKnZ1atcguDfRs3pVfYK+mmp3lVSmtGJwl9
/HUrDyXJiORCgdrC0GkkyeSVl1kdLCbxafpz9ZyhZyPMi70gedz0BezVLeok
Q/72R/8ZWPo8BD/3R/EtjRVXgtDUGdMBOfKsa5tWmS48Y43dS6e+7l7S8krK
Ac4wNyZG7MQPjLDRQt6mOBh+uoTWuFwNG9E4xWjw8Cj6YElb2AzQ63HwAZ5R
mRuSVe2WlYWcWj3JuEkW3zFXdxgmpIVWwobBRkHCHXFzRUvgCHpQIkYoidK0
ci4bfJHNZa8E3qGGCSwEn/PYoYFwLDi9Ilbqc+7KqcUwWtLTB34skFYUJnW0
Yxe8kxeTWLcAi937tesgUZdEvYN+Ge8CciiUie8suskNUdkafrHn6PlN15zz
x4xvQiXctsiq/UaMXaB0RLXkgXXBmJN2cqDRGBI+FZeAt4TbFxSNtR6xmpIf
kjXyajfqn5/WJBnyqqB0fHCijAI6JMF+GXD0KIHuHBXx9PHFBeRzI89zDvW/
oHSygzOekl3tMjtiDOfRB9QyKp79S1F9tZ+4z3soyh/1Ai6kTGqnNY2Z3yqZ
8uj+KFhjcRoRAgrqITS+siOApHp7PXuqOd+/z69DUAlaq91IxWfcukeOgqzz
fCFMR99sNqZTXORciEKPeK3o09xElYvfSZLCx6heTxapV70gli+pEMbHOhfp
urjjtdPswnVfA40PTE9ShHEtKlFA9She0qzeiAZgZ9yWDL+sGkdgldOv8TFF
mpqILjufFtlcHIQLMORCwdRp7fndMB6PxOE77Dp2BrcI8+lx/cBHtqhQj6zu
3v0w6n3NNXgoTCi9YCQobrbgCRwzSkrYKSSuoNRufOoEpvJiWM6l93dZ3d5G
XJiIQGQ/F34N8iTG9a6oumoxDwaufNQUU9oRVrkc8Un6QhlBK3TZPec6bY83
NQNDyLK/1H0BuPQbU+tvdu8/4CI5d8WX9hDs3sqe6VLqs06E8/WRqiEze1ui
YV3to7PSf4y3ZNP7zGVw7U8meYkddCnqTAeuem9wxFPn4uSNfbk7VzSeti6O
C08owengZdBRjbK15F+9Eo+8mtkDaA+VkUkq18e5R/ELfDPdtOerZacHpQPU
9Rg2d0TPHxksHmaN7FIWF0QBr3NqJJaz6VSA/zogWQ4O3tSu7S6bzBuJ4tYF
WCRcRvwguHhDJkyWnyJDAL7ERhmNelcO8AEqap5Cwp0BGEdZmySZdpZsF/jb
tCrlc2Sxmhaf+XSs2YyhE87v6XRGz4wYnB48S+zhEfZ/eaPSdmjTlPyw0kzL
XjvHS2Iqv60+ew+OhfiFgK5NgjNbuAeJaWWKR7+L6zhYHjggxM7cfvp/OwGR
JxqSu0DHtkhJ0XWgszdFLwKqt9Ke1v2AXifeA4JxbIi2gKTSoqdJJZBzve04
c3HDCcem5rFlwyoZ1m5sK8MSLsdc1m4WoTOrq9vZljOZt+mNP+uCUxv1zsDg
ei6onk2qqE4Ddfhbb9C1f2blXuedsXkUALnfsiL53NUf0Z8GsLZgMNzo8Nl5
iEkgP8+YzmncNCyhdYsQgIrn3F3nsM95CzwCJDslXl7/JZsLOCkUCw6QsUs8
/ky8YoOTsWJVoKbsC6LfAkEcEJYe81sIvCQ4D9m1t5XCqxzCEAIpEiUdXUlD
ck4JjCaesZxTx8tGOdPaNVvdTebe04nu5HeyPiIvboy94kVMzZJBElqyWXYd
NzSkqtrO7PklHJ3WGev4QXqJvxmMYtDQCbuF4ZnjVrHZUQh2WtxDJur12GTV
IMz0+88NJaDn0BnYZXesIPtnvXVCmDziXIGslcAvP+ztD4F4+psEfaVAjA+B
Qho4PU2msYjeSqzEHbRBtFJPnuZJ83IAzy/xueqhvztwZQMahfVerXDdJ0oR
bFDD0YxB1SnHYZZ5tV+DLUrBKyLDDcxQfph/DzJvi7RVngebFGdpwzVHBqTR
Y4Em15TwGlYbaqgccqho54rKhoPcpv86a2eLATiHvsjnCUitmUsbhfxahj/W
ZyoZRZoy2MY2gAoZEu0054/oOZ4SFAanwXPpvyisWQp6EhqVOLQRcjQzr1FI
1ujKIKPrEet7AAfe7CvJThZRPTsDvotY7v4s2ld4yIlAi5XINOOcdPm3ByXd
985KPgFQxvFLVDnsSTjuPyrtzfpB4kHGfYd59xBtWh75yWyhpgaIwQrac1h7
aB37b3QA9in+krQdDBd21F2EQnwDzDhVyunv/XChfv169hwH2T7G2n3mLDyj
9VPrAv8IkqMBKODUK5SQOq8LC0F6xFpAg6SbS78EZtJnCR5RFDDfHSs+tUoG
2R14rHNsoEnqgTC60ra5Yo/iVmvUjJ1j7OlkmEZnUz1Zfg3WsTmu/F8HWtcp
t4IeQeEoCEUk3OmRfgnB2PH4oUCqYxbajI9KSOw0VVegLriX6ILXjCEVM/qs
JIqLOaMjU3OmUo2QkS13+f0QWJnWV1d8oxKqo7k0hNRezMVv6lFjaIl9xyEB
py5EVgfotu9tgN+EpKqV4ajrml7ORRlJ1OWGb8ho6wmbKYyMpZsiaWmcHCqV
/qnlMefCHFdot/kgsi3nHRa8IjzblxYlH82bPjQUWXcUbSv9gTJ47VLkUa4d
sgdKN0lq84DzmAmc8kUiWn8z0C6GqmIZSU3YiA9in+88v2MAhPc4kZc/cs4h
HsXJMXGFYBfMH52zd+mr4fWpY51FVTxk0ABlRUl5n/RufEKmgHidZOODO9Vg
P+q5pS76w5CgCNhC5+N9Chwdz6fvenAMfn/DTjmEXuHNWwtjbGxwqOGz4J61
Ntqqo602Raltta2tu9Y4OddJgKYYx17B8Y8NODf6+SRuei7VcIr52x7wNUFq
hYvVSqLBzTVXOPDVcKqgP4otlYU7nW7yLaX3c9mQ6FHtwK8MmKJdVdvlZbQV
5Oefj2nvN56YTKtg5AyKp5dzfh5BjH2q+9XALdYEGsKDGoAxu8OnQA5VL5X8
/89MbTiZhbHzZQJmx0NJRk5pThiz2K/1LucsAKXiO6HReXVtBGJTldAMRfKT
CDZScwhdu6GfT834Xh/GsD08uQN5odFeRDZPNDNgMxLUOgrd7WnAzOVl3wKG
na/XW+Mf8mnRRHuX4nGy+28kE4QZUB5YJv8IamoP+gxOl4p23eJJq4VJJeQu
xyFBlauc/LfMVOjrb8+QWGp1o7ZpRae61OzJaFL8d9A9i73jiQSzDD1eWfdz
mQYOFIUbUyUwUln6WNx6TC2gKJ39FGgwNIlPn8txZGnFwDv/YLMcjH0zl9sw
/Y01Q3lJD4Mm/sKGfh3ld+NIHa2DEQ+FOZzmMEgQFTC+5+GSXKPllgZVf2QD
88nT0izhDo7uqGJ5iP/KonhfQtreMUoq7wNDkIaOblIhaYM5saLvwEaIJioT
b9yXHMZY7QcxB+879leZQ5n9l/St71PeaYnt4IHRpJLkiEJCcnwSpt83a+i3
kAPFVl6cPNGIoIO3lFCfL8mOeQIUSauQV4ITPiVJN5XrxJ7PnPZzUN2bXtSn
vC++B689WhcdIVr+9/Pl0k4qiIPg+/W51l45Xr0dEQRLfeXP38TLEDcPGB50
RjfopOabU8CReIJMI7NUHrnIm6T6VmEuLyx7iXDFzyuul7a9C8O/LibIbm76
dkvCJz+NRYZAMw/76s64RU/i/0Is6S/Ft73d948XUjjT615qNma3FwD+3M9N
4f3pNhf35IGus0dyjnPIKdS7U9GIjmfFBTZu1TwPD93n/h/bvE7K9a+mtAHZ
j5r2LEMZOkJn0bBNjBdb7wpnBpZNbfPrtfnZltNyyV9YKVQIfqljVUosCLvW
Cq9rpnwONTW61fK5vYLKWzVFxnlHXRlWJ6/bQHdvTm3yfawjX118xJGuZFlJ
RxCQCe+HWxTYhw11f77A6xScAUcbtwIexSkV/W7gJWpPRNZsYvnYSGt9t93i
KlgAlsaOdrcTnabMQ4jqE/+5CvuQGRkcpDWIDSpcC3z5rbO04eU8fzME0s2U
+PbIiCCSdBdVfo2W9IFXWn0yZFqrH78bVFE2Q5q6HtQZEdYAB6rftme6a13+
BSMk+w4Xou9F9FKKyWi2BQQoXX4+mmb/NmEHX5myzlaEgzdEgVl82Aa2fls8
lkNudOIkUJYvd9rTeshtU13jW7TdRx/zuJbM6k4zjZjC+FJOf15+0UqRm+7O
TMcwffkz1Qmb6gBYlsPfXI17AkLxPWn2FfMtgwstO8Gr5WsOHYlnsEXmPM3l
LgTa7azoB/ayDEQeNo2Kp/DG9Ujjna/RC2QfZsnJmJxkt0ptPi7q77DLROh8
r/XlYAFYFtruVTMqXBulfPR6FgsqONebY3t61A5w46bM4j8iHVtV5C0MRYl+
NFNVPgCdAA3wU2CsGO6T5cleLivaPevYOhl4dj/cY8QR12gI040Cf70t4kWd
x2jk5Cpi7ssyqjE7ytoms73i2u4gMtXUhZCJk9AjzJs3ry+TqvPjWvPmQxqh
QK/j/4bD3wwq2izCZY1ytkzwL4pwa/JXOkG8TouC0mgG30gajwfw5yGwKmtl
fW/aNmLs/OtAZFRPE5PR/XyoAY2tsmvpudlYf5WXrpyid5siNv+pxvHJidcF
ZrvNJTTTho/aVKKPdMcPP2FNU/48xCqTqG5geH/HQlNKnVQbKsRr59kPfnVw
8f8Md8jJHS73IDaJaSIdw7O8L9LQTkmV48OacY820Ko8w3Cwgw1DtClgWfR8
pgKW2K9Q/REpY22feHYWyJrb1rIYHyAbkaHgqm0lOfH4XxaaeKaJw3IBBDWs
zzifhVjPGj5r0Jq9V2bpK/Wq7zMDcpHB7iesQQxHY7M/dx23R5yoArpQwHa7
XOJ9dWyQSPJVBJgdP75R6epkNIu4jk1ZWvQ2oFRXY9AyDPDJfH63GoNhrEgY
myk20/pebA78tRVo63xdOo0JU6LoOt53C26sK9LVXofVC2bNwHGaQXisu92/
65O5hiDFTGjS+EFc44n75XhXF7wOsbKivWa12yiXO0uKhJG6NT01DR4gLQl6
lWYjDqbA+ygM+VjZChmsp8dEzEPtXp3ZZJwaUARRDW4GhxK5+f+XnrEfe1Nt
DJ9oUJp78d2g9BMEVyaH3HLwclT+i/GUEOoHAv3QXP5R/3oXPSSdsdGNjE9V
+Kl9VvFCoHNB2phP3XWhKkGgJhzVX4lYKBE0BarxAfZdPlJfMeFVnMwFObrc
XUofHl54Ig74togPW/qbesai3wTUZBYZebKIU6cwfxK66VUxk8rp5j+BJVoW
YpDjE5MG3tyCmE8WHztT+NKYMWLZ4tY7/VneZg2EZnMgXQc/4DcRpmK1i64t
uKUrNcUJf6sDKDNV5TPPmSBZcU9mejAChVf6JwIBOJRg929NERqS/AsbJWGs
jCUDe3fjx3qp/6BJniB6jYi1gwqZzfq3iMbU8L+kOet/pewsPlQVvPHhCVdx
/1wQHySSKgd+7kJJ0462N8bU9M4P96LPHnxFWoov5SxwxkQlOcNfmjjJyRa2
ts5/+M2HMmUHKr+v3mjUY3hbK5iS+tHqet4fVVFSlVnccO7EO0Hi6TNNAItT
5NkrFK5dOwmnumPq+PUkz9iCkwPymgJNF3GkyCVt+opuUy3GfwoMf4BS/isi
LrQmh1TeMM5IdcQXvR9yxPSItP0iChoBmAJUCn+dA/ytNgiQk9qQJS8HyrBI
YdCZIKBeo0pC8lZRDyCi4CEj/VuD4dRx6ycmxJRA+QCGJ42dVPRM+29Vmz5r
Clhm1lJLumyVSvZs3RNpvNKBVe2unttLS96Av0/ihmxv0jAEYap8+s8jztB7
IxmrMMAJyhT0upj6+vUvIqOrrwAAKpTJMRssOxUJ5ILQlXU+Kju9F0MAtGsC
3J6rYctzucUoE6ueJFa7Kw7dgqu3TIjL6JjXXEM3Tq0Y3nl+jyXyhK4X1nZy
O9UpbZ+Xe0QvaGSH//9DVq5c53lX3x8AHVIT3fLVquUqFwmUMywSwdtS6RUN
r7Ck9iLomOB1Wu/DE8lo9v+hoDV6xSjsvZhTfy7nQt+m1NAvsjfn4Oh/2/e8
VroX+CumRZFzvAGz9HTGHTy4ekaCsD7oJJ1dA8ktO9V3L+eX/jCH9hBfSnl3
mk25NZw9zWHfwA4i3ho1ZMDlJpvUT1ITNWxgr/tADYDwBjyiXhFfSWFtkbfm
F93YnA/dhO3EZWsWEk/aWT7RaUC9ua201i9QRTnGh+fECK/qd/mBvrL8j4/j
EEre8IQGibAl91SRan0Z9GVOVAwpRi5dzgWi4Kj2Obe+otMDhfL0eP0r9cKh
OmugoUGsgEw4zN5HE1toSdoKXlMDwg4etu5DH3COKzEe9rnxRhywy8KtYiM4
wGB6t/XN1RRz94W/eKBgJR3kGQx6l57V2sO1KqLQrzImEKguZMxbVNlnQYvO
wTXfbm/ZrZOOiTyMK38keMZ1mPNuSriReDAtPdwpxsDmfoZK0kTE3t/rGn5x
JlultprBpRTLRbRdOUvNncCQHgd2ubcjbptVKK/75diMEUMsU51QeCIzH08u
1Sbk3fTJafwbxA9Ao6ru4l1VEnCP8dnO6oYnCAkDFjO7AT+CBTcK4pih04A/
Tt88mV1uxi8CJVDPCAdykfNAT28+szvO+5R8tfxIuaQdCEiq+1ZHRvfAkzB4
EwsFVt3qkqO7IiJT1HQtPITgw3f6k2SZikcIzItp8+73yYOgh4gxeCBMpglV
iEERmcJMOuyCZwYq+tUiw3PrLyr8fZKD3GnmDEIKV0WHjf4ltQfmyHo4lOpA
/kxMGMQY8vg3RvubGnqsqhc2RWIpIoPfsprEbNE2Pzi9YD0h+JN97LQXWU2t
wTD8p5AFKJ/6Aocc16bEJ2kJh467eEIEtJio6LWn+MA7aUaXOZ1eR+NroClT
oDgSJM2wNm52sjSiiIeAJ1yIVLUReARmhSGKnu1HywYnKvlcdh8JLKS9n0O6
oP5omy4yEPgvNakdc5cIDGTDwDF1NngywZvKeXoSPHdGilGfHahBlNjz+nm7
EkYylDeqYCI3HLBgDChDOfwL3kRFZo/OFcK4ViQlYH1ckSoYmFC7PaJJte4W
e/zwcSVMdahlxrxlqY+YU60wCuNufp5D3jayQ5UoP03st1+JcdZKq+yCM2FZ
GcFyFnBS1SzT9SHYEncv3HuwRLZJCck7DyjrMNsOgrXj4LJ8nqvhtuFKjX2a
ChRFIvzqRLdTjS1V5JP4oFt8SAwU8Y2CMwzosmZtiOf1t0Yv+k90ZEcU2o4H
027BH4Ko05+SGxtXEwPFTw+t6VDilYxBZ/Vg1zkAvS5ar4Rs2RCxx07hFolG
HDWY5jorcKuhrWP9HvoEP9BWFLSUg0nqR9sL0WLRWrMuCpV5UWm66cFAsjAr
B429RSA4CPzBWjJQ3rzXxe0ohyql0xpkdGl9+kSZfVtazAxkiBEGD34vyUwK
ej5ex+3dcKyJvx4qJxOZ3TZB8HJTiZEB/UYi7fgETxuMK3RcXwXWttUiRxcL
7PDbaykb1s9N0Jc8/kQAMIS0qj+2jucue/zbBk0LBa4FnlhDAr1/VtOiyXP5
uYtCx0Fr7Rn3OgQl589bmsnVTo0kRQynCVV4h+pmuYhOlcYn90vM7tRAn678
++ehrA9mffzQEDaU1G5IUDvmUbCQ1FYLi6o6unwtisfU9SjtzcXNAx76QrW7
cHrskvPq7n6I8Fj/gx+WVUdrS+71Dwa61SIcJCSUfeIbj6wHJgxWz1IEhdZ9
2ElsV4qiyaBspeKPCMA//sDFT1NW74sfyQSoL7foyyaJrv0mIffU7XH+cLzd
L5s1AFxWoqiLbpMkZFU4B5t3TiS0wb1KmIJSH2KL0HoCeXgefljbIcHSIQme
oxsPXsYFJ/xUqlu5v7RBLpL/WWZqZeY5WV4dWvIDCuSYeP3tvyJ2Dqhwn84v
IdVF3JyphVRXQXOzSN3seVCyLaSSemF5UpVEg7VZpcFJ0MMJ4gNgXx7wvXvB
iY0zU2R24YTzfu5HrdKcywQHY35yOF6sX7juW9ZoccYFrLBkg+5iukHbtpZn
HvDa/+s+BJSqK3mVGJGR34LcIVy42sfh8W+Rq11pC8hVBX4f+4/KDVjTfh7R
UZ62uw7TgPyFuvXBRBQFYKjiBpeoUOYN/K38PIrx9EESyxjW+ZuFd0kW/X1a
UMXG85X3lrSePgh5BLGPNoApsnJuTBwqDTm/NR6eZwoBnK3uRn/OmCNeYpXR
a2oF3z8lheGFnfEo+bskqmQdYn6p0/qc/oZ300cQQK5WlbGQaNwRXgWIxIOd
R03HYGM5XyZOmmaRXrDeQNN1FD6CCoJR+O02pHz5gb40miQ/fTUbKslKha+M
p6S0UuRHX9mmEU8I6II+0bHBk5gsw0xOBR5G/IIqkNA26fJE+TXbNg2kMi+G
r1NFYQuodLwzRW/jNlhd2R/V7seGMoojBlxmdXiO+wgI+unUiDGcbaAY+Usf
U7fCCe1vqaGAgriE5/NtEN3k6TTbmlYsUeCjs8/Ryt38szV67mvVaxiF8BxF
oLxXzZU330jWZNcatYZZSaDCaLZMqHuwRiaOqNg4bAQ+DlfBmFotwJgnenNt
imemb/t7yZ5n0XxDkirzZ1Rp9JfhRS/bKuaN3oDz2U1pg5IdaeoxHUUEUwgM
SPyBGK8qgfU/GOPX6I6FxkYdmO53e2oXuz+4FAyKxoLNJDXV2PH/7POiIIaf
qNmcDgnkfMmjHhYhm8CM2DJrzc8y2AVH8o2N3c6n7/bBOdg9J5I9FFePgk9z
ObQ0lMZ35BT7mhvKn2alW3fLLO13NLV6nrWUUZSn/NDw2s5tYqLeChZCf9ER
vXKF0pE0QXMqQBKlq43JSJcvZlqo96wYhNqk0+zI4lcuscbI4fErBHNjZGk2
zvKr4F2JbtrntHE4GwkD2Xifvrcd24dhuQE2OaAE4y1A8o6xoxeXjCYKXNT5
sU3p9HFoi8PvAcm6VNPBvoGgNGt4fYWC+/56bBvhw3d0ok9iUxSLZRXCpunV
Yb2Y2pFHlqaeDA8qp9l6Ior3Dnnng5zUZ+s7F3xEZtFghO2zJAjKUC/3Jc0O
jYaH9N0pz9gWj/mpLRb+sNAckLRGr6PCeZ2Cf9ExB6Oqi7eySvTs/AzNrSdT
Y2oC2juk8z7lXdh3rdaC72zmkJ5hDfNxn/QD9fldl5uI7dE1z14RhRh/a2q6
fNhpecQOzIHhdd2exabWdtFKg1+Bt1RujvekvpxslJTzh88WhSVnGlPzDwCB
nlf5yAs6V7gn+inB6gnbTbaQEBPJwV9kHdiv7Z6G17TCevDDk5Xiu3LiNn7q
sinS9H+B4O9oEoMXgGlTvB1xjtNV/L9lKL2IN7rT0pjXWbtRFxlfA+C+5pBr
oI/NXMJRU11cbZumpd3Q0JZ2M3RoaVo8eQTP2E6XzqA1lG+Z2m6fGJwiiIXp
7nCyDhF3LoudARK7XsmGD3TlDYV/xAGsQu1e7I9Qfjf3/JqQzXOcavAofR6H
5v7nBpUbgwM/6jfXA9jUmOap6kbt8umM07Eo0jtg0vzyatuUFcoKQUd3yTQ/
73QiTQuCKIrcaElrTvmnpQ9pYFaHgHHuECYdOkLg2PGbQVpDqmcYqCCBQE2m
aI/l6LqcPn7yfYwLM/H1G103t8zk+zvT/nl4YfHdlHuS0AuiCpkYzQ8MpRTg
RXQ1dZW4BYpdU68+VwUJaJvnoD6tPX1nylhrgsBgR+lmi1UtmI2ZSHoi8Kz3
DoH2oZRzk7sM/NptVgExQZ2Kvk6TVDJEICHrfyWQA46aFYlMoVf5kEMfAJ2z
VIB++35bLyD0ALyZiFZA+rmZnZDjpYZ4W6JBeIZ4URTrpf1h9ZNuXs5AI4UQ
7KL8dmI6KoVdkRZfR2ibjLH63ihnzwlb28MkzUcYekhtMU2hZIcARjuapjxI
zcEaS3PX6/cf/9oFrVSwBHekJpIoT4YRPOgP2OszGbjayyL+ox6ulKeKNeOG
Adjqslhf0qcbbZcNaBgW95bh9Xw2U6ALe1U/XbIfKHqOcBLWla0/w/DSa9/Q
gHugc9VT83w7pjGpDANR22WoW+IT6iFRxdrpw8zh553fLDzQ5D/3UDtbN6ZY
5jbTlTFDCuJVWi3Bgw3DHm4BIP6rBY8kUS91dC1XzzMmT/DV2M/JavroCxEM
ACotXlIU4Q+9GphP98k3/iob8XBDsKLe0DFXHt4uFrTQOFSaM9gcCq1/rxev
ufRo/HNOsEi1lfOuBqz52BpuzY19kugmoC//Z9m/iHnndaM6TyvQo44aFPQk
m/6U55higMjyZ0r6BD63P8rWEToU10h+r5OMnQE9R7yiBvAgCv1kf/rXzLsx
xqeyAM0mZGjwhghZOxi7XuvGD+aNBRvVd1QQmBAk6/2UBCusIVeb7ND4PaJD
9f8AXSH1dSSv71AzAXUAij7Z5JNnwTZ0WN2Q1HXGTGd/y+izu3oYTY1UOMmI
Iok0he5Ns9aoZfyE3cUjnABSmp0SIEpW886oyGZZQP9FcgmCvnDtyK1tBXZa
RihAINIu8pvo3O1PVsBcI7SLlKF8Sso5vvjtqmB7DZ29Evo7c7ILdiUp5NQN
qnMLr8c9t7a359uqR1VVuw+xfkfmILKQ1gl244+OQIQ7qct+TSVAQ4NS2Qk1
luQt6D6iRRJeM96H9Ur5nFCKFdTMwXcSsBbpNyfy30GmfZOULtvFQ7tVyE+Q
Q5x22vxR7EJCP3xxwK43NqspoZd54Z6+/cgWAV3NPGzPjHPc9Mj64iyBhDlN
xepngj+dxxDfQY9M1qsAPB2R6N0qH5NkGMQbW+O135a76vTIDK62VNRQ+mnx
+wMI8MHl5oET8Vrf1y3XlyBsQVWLrXOqO9q05TVq1mLnFlp+k3rKr4R2eJgo
cNmORJbRiPZ9Fbvh+wvAj/tsTovwCAyEtHoUiYSC3UCMXHAqg7RNV6biHga5
qw7BwrtXxPi/v6nGXlLVcxpLaV+K0TOxEWAVoX8RN4CDb/kL5uVzkjNgKobo
2pYhJuNdvu7IBZWq9UZpP7PRiH2g412+pVe+V7d6iZT5XrT/jt6QP25IYGBo
LhA4b9g9M+Rk/08KvZcCCZ9/6vgsVZVJYshydpq9bJF7ZQcvqXoVYgXttDV7
9SeSNiJZFrFFZrq5yCQQZN0UlfHXzjRIG5vvD2ze6bZTb5hreH4pgeCWao6M
9ji1mHc02IY9yBW16/CEiAKLWTrKTozPy6QHOdCwnoXKcGCL+k2pU+OkMuP5
e9PLqwBtywz98Yo/2gJHY5PTvQ3qPCy7Dx9cEtlttIi7xD+6azCyxmLkIvk0
SWFeJ4Ivr2guPiguaecRDwFtXbKHXt2rzQOdSTJU+eNVfpaxti2SJanQXoaJ
O5/T2ZN42Wl2CjKVrTKey74wfPQRwQhOySJlMK+7YUrfHmI1xprID8sWw/lH
yXKVEEZesjNHfBlZQEJlbEEQdq6Cvtqdt2QaE5AsJLx4uc3APJiaElaAKsW8
iU8Zs16F9bnOKnWMP3A+cLcLL4wSDmXO79AGj9mJ6UmxZCsYKbVFBdE1eXYq
/gsXtEH60Gb9I3OorTk6SDOb6xq1hRvx/oF2G2IDJ8fp9B9SQllkJVDrHrk7
nxKoXJnfKYqJ6VmUtg+b/MseDRRj+D8LKpH9QdR5QLIl0cLIMbcZiMS674Eb
/aPIeca56lh+FI7wL7PskolmbZOpd5MNqLpjGwuYbLw4ApD5f9yqzNCFubL7
p3hiCgCAW9oElsOnZHdzOnDsom0tHjBF3cCqDiQTtMJnaKlbUReiHdsiEAz1
PxzFNFQBVaDQtlVWO+Oz9jJMjkRlTVqMkJKr2DCkykTC/rVRvur+68zvzqmV
Av1vNZLOxU/ne83KT7ndaQ4pm/+iDWqqd/6j40AQa4fPtbtpz4L3AFaO79Wi
Q5QxltZjPq9Cw62bAa9YqJHJjQ51Ln4UlPABoxIZTJvLRDlkhc7uY+++E2Hs
oaN+hgtrIHo+QshN0XRj8I/M4ju0nnXrrEPZ+FsBUQyVK7jp+TeRAkx0anRU
w+ecxsMWAT4HB5YmcftsE+ZXYK1UYoMA8mGN82w0ZHfcBQUswfRf5h2Z7sjY
2U4bPAlS3gPJWCNnf/h7U7SQbufM0OiRK4lGZe2SMke2kiEYbCEOURvL4YzF
ZFPIH001xz03tR7IyEoSYmo00TkHi0FPFG8lyQoIlQHtfdkr6ByU+QSxf/jP
5HR1NbqOhBcVQbLCS3X36kDwoGyW6X/cS47ZXOU0376kcQPoPmAS74PJ2pa3
fDRq662bycjcAVKjaqthZQXbe5PaXwkOzhhY7mUFVB9IvaG0gD2g1saKITLo
2tw2wzyrr1sUqGVWq+zYbKI9mblGwoUisulramFzZj8eyt15LhNNSEIjY/J8
v2Qm5KdzbVlIbmv6wvwU0kP7j0KJMHo5xX6ayq7G8I19RowoQZHhqy3s+1OC
4pauq1zhOCUspxpY7kGWKAFWEq/Zs+u9bC0rP2vugsg0YhgbK1a1K5n3mTEj
5l3NccaPkWHar5G8D5pqSHkwW+cATIlLdvZa+8Cck2NAmunP48OSTuA/2iWH
S2YHpzsxmtrree9ro4mOPEgdSWpCUZRbmJkgtrILLDuE86EcnfwYwlLBcuxH
4JVT6KnvqKtqS7Hp/8AW0XUdrhU0yS+qFh4kf6i+0HXnOds8m7VB5sbi6c7h
T24Or6ATVYoKkjUJro7n90trDXDJPETwQGoTtGqHkRyP5kY+Pfltehq4k7ak
0OG6mVH6hr1MVeuZCoug+Z/0RccjsRCHbXNUjR2D0XA8uwKCV+XAtdX/rwJd
reCSpRfSNT1+ha2GgivYTt0HNSYfHaHN7IwqnwqvNNaGNRBm8xmoFi85GQND
3fQMVYC/o0XfHprP1lV/iO+1HJWykP0knrFptmoacDd9GfodzrgEwayVcTI0
GuEKrt4qkhYX7h8nkm67/SEllNQv4Ei/MZMswryMz6zvag7SjS3EbC0nWY7K
c4NDhb1Dzvlb/w9ivdAOJEm6BWYbVe38MSexWfY45D/vuWPVusKtuj2O3LZa
yLy57hWAw1Eh3v/C1CTq2qQL3Yf1knp1WVXC/jjWunr/+izP0t8WFYh8nrjI
iwF8vLSBurR75vFlBhl3H83ULqm8f0Yc6D81aczid6kY9Ckw1Xlcg9lZ4XaG
gHgXCBYYGwgKKkhOm8HnKF6GvEQtaVQVIk51ILwW4G/NytPvbYCDdMTL8u/O
SnKim/JaYOaos9RhazWvC0PdUHCci1UFdMkOG1JqPGH4VluJiYmYBXHr/whf
3BjrLahFugrd2hEj97Io7jO/gMRyodW/M2YW6ouX7RtNAgiNFPiPmMRSdV/b
m7AkqyLGyQ7CftCdXBVgmdacHaFGwqMcyXzXoBZWfN03cRbQw7CEvA3bkZOo
Vs/gf9NdXS6lX9Xdsjq73y9sky9IZaPleUZF0ZICwUzUdCNnKjwy9feskUia
pb2e+nxq99Kl56nKR6CQ7b/heHV4XUd9+QKKYNR6c/FYx8aJUPFNx2N/vi8i
n7kHyLbahRqjIJnr37ZSKaJiTr1ldhXMIHmUKG5XTIQwneDc286JTWpBKT9f
C5oxlVL8K08EJ3N+HdUNV3G3VxmWH0qBBoXyNrUhN7MlIbcJNV1QXl0GU6Dj
uipSl1wM5vOkIQ6KMlvElnHR/E4Soxq+j+Iu5KtBwxk8Iv+N/lg1xIXAMh8p
RF4q9b/4neSadClg0e7dR5UNg547NHzxHRcBUGy2I1T/Mb/+fqB64Iv+3tLw
xTKoGzHCQGAEgSxWKdliPE7ghZGsodYS9N2/fh9ZagSmU7tSd8gx2pwcjDOR
zTNiatsB/Ge6sGxnrkuH9km5CSJFre8DGkO2Ae4ZUccLo4tbbnP1WQtLZQXZ
wInH8Z+8OaovIkzvsfvtFWf2p8sv5AFJoXlkKCfES5UBHtvWnvQrktQmORud
IwQ0qlonhWvh3KNOkGnHq7Qn7Ef9Mt+QIM/gFa1a/8+GeK8+KSIM+h4vLCz2
IY9yp+Z7513M5K+xCc3/S1n0WrAsWoFTTnXG+UMhRVqG01VV26r/bqyjjng+
OklEe1lYXpu5I7ironciCgayODAmuYBjzqOwldiDFLHHn/jmqF098sqW8v9Z
b6UJtaJdGT64ABiHf1Fj93xkMrm3fZBwQMwa5LZRknP4HSQWlC5Y7cvxzsnh
7mEJb1IzH2Ejkcs4V++8iN9ZrxfMWJHA2Fxkb7Q2Ny4CVUqrD2rWD/kL5nQ0
sFU4vZ1zm1oPJOO/wHgBeil5d833KwC0Dv18fm6slZOa1zBHUvZ8qeL4UOQw
hRq80oYmZuZac0R3NyhiUGQj+vGdnwOhatma9ofgi9VAQgSKBMla8FQaHajs
OPcH8isMVsabcNYJbGH9MW5jiT1YkHMy/2RE/YewMhXbY4EjjTu4GXWWJT6p
oeEpsEZPl5Sz9eMw79TFTZxFuGpfhUwJbNkBPOuVGpfxTXV8kZrAd4VAayzK
z/hpHVRrKoVPoodykL0BdEhb7RcM3taFcfuVfg0Aj+9aEm6mZhGofrMrPDgE
FBzVuXSoylg+Y3z68YnmxQDLIW79+vT5SQGEF33OXV50OabofGhCwA/mzl4y
DzIMxj9ItKBla84MNHaYhQ8xjXSsUUKiLREn+TfZBBkCSVfgQx7yCiaexhCg
Ix+aktl23vmSuFN8TdHBzAEqsV2TQY/fjoNfIFeKVwpygdn6oomuz/cVH7bm
6CUVm8zqnnE+OaDSufnTD2Jnm2U7c2nnO4F0del0afEM0d8hv0e9PIsCnYBR
Efk469GfwAhSQRifDf30m5/KrmoPaai5hVHMTcbcE09r0+hKfyDIC4qqlIjI
Mpl93j+B8lRmyExQudjEQ2mq/c0Yp15U+OYCz6z86rK6foZjeQDhY9HnCCPw
+FRDzyrXMbCMADF5DIWo61sv31QlxeXDvIuitTI6wsPJvMtcm8fTS1czSSIS
/2DPZXwx7+hw2tIhXE4CEBm7SrgUObj1BzaVCeiqSATIE3/DLOuxcnYP1hM+
O4aJS4LMasS6ulqy3b7oMJpyGxFoUVijvv9L1UzNLvTvBuyZ2dAwqmPVSS7z
gHKDON/xUKRyGYGX5a4a4PbyS4Y4vYTZDiHH/tBUOF5ClNABYcAfSPdgyKla
b8wmxQamzXBfcVBjKwvzo8Cu4DHJSy5KoXYk6dBUBGvPv1T3bp6LCbIA6F2J
oX0oekgBZheKnu/WZ1VEUyJ9E6OkJrL+NLafeBqB42j7phX8ePMDLr/ZM/aE
eNgW206x9hBtjKcyRoeGBYRiEH84zd6cQHcyYvPXTv2VQmyyNreh9zr+u1wN
wb5Ia9IDy+iOqZL06+uybxTUjmfivlABERHC9jOqt1AwiH18/H4NLPrb3KDR
loFhjLQclnaEg3qoJRyoJItxQQ4+tEAWyu8zPMc+iNJQVaHjsxsCatvawGDn
tz6p3zDHgleQrD3W9sVpP3UzsfxC6yCM3Pm21Zn+BFBnRRpj2r9iBvPdF2x+
gdw43P4WcjRrdCdSiFyZBwYzb7wP/XKjbabS7Hy51o5Yl7WKzlvds3o9v2Of
XuTsr7OTEgVSvxbKuVDTRyo2Ev80Xea8e511cMdQuP1LjQ2foJAL5+T6abzg
7EM2S2Icp9POgbDBuobBDfxVMTohQPjieq6v5WFNWgbAuVTbp9me0zqnMHdx
PU16h2AfUXRdlCCXulzSWP7QD2QyGNK1obmo6M+xJ3VYJp+JLzLsqOd/boMO
2qElJ4rgLI2JSo2tPX6eGJIITlr5eIQ9ms/n/kkn26lYnykjcmeyNNaTgdZo
yiugY1SV7j8NKFE5A6R11173WEWkLKOGU/KpTfC9CXFl+epSh6FiXF0Rjgq8
2fHsMMkEbcLIWi9OG2qGXeZUp5XDCkYiUZKHzFvXkCcNmDp9opxgnWxUajyW
mneMT9MvaXVYKRgI9tCVO4SyxhlnRUxav/pFCw8KfHkTgxZ+vaxd03JssqH+
NzyKB9OLidie26u6aDb6hAqJHoX4wZer5mdPEACxXGUJ3yvmSoRRzgANu4bz
a+3Wrn5FPC+Ein5sysSszk0B9nXy1NjC9PWqsVwYyxfMTuSiN5tMn65a8Ip/
i6jVKBR8nGm5/hFaomVKCSpMR4kSDi/14NGVaY3pKe9tIHeBAjRTtxuzpUBa
aG20CbMzuiCajoaJBiniO1LHNneZcyCV4lBRjJwN1NXRXWf6uBg+r793RAol
jFWKIlq3IE6qMikxxjPuvU6zcAMocLBainzeZWVMBHFT4gZCx6DaNs8/Haq9
jQ4B6q1uM5zjWYVhWyDBacQlz7gTqZyIJhvTLZi+HU8lac+cU46htvhueXgh
/AWnAAMPY7YW2vMVF239YZmb/+VrkG4EB53oyYSahIRj6vNLSw7pv25aQclG
bbDkPmQZB4QpTbSnUyWaoCq6YCguoMqnZ6BT7/fS07fasVJSi9ralJUFDEfk
roLgRMzPt0HHuGXyMUBOiNc7LlUI5yuF+CdidhbbF59Z3rjGqW9KFldpiaIn
NQbhfoTKcrwX8OXIw+8QcKK0Kyxo3yorwWwsPMQ3aFh3HSGUreMnC9iRA+/9
u6BFHX8zwNlBafH+rHCJLFip1hsLeZZFhaR7gznjUlgJjhKjHxPibYNSSrcM
mvZGBBzRhIq95lWYLasInUwgfZDhNIl22OeHw3tZ+Glq9aDgwXFeuWVV8h2K
lJ6eaMrkBoRYlbvpnF9Z9z/28cvyITl+SQqmnzLz7vIoZKUNH4GX7PolTAGx
6NvBxvnswqmLEHfsZBatUAczTQo5Ew4iHoMqipfLC2xGuHYCNDBAJh5Fb9B1
rcKiVLE1Cos3ZGmfs8bf3yUDaGI+AgF7cxnDmzUC5WBdyUryBXy2WK61szUb
P1gQb61g74bGYzwbHjIl7P5kbtZ/rnhzakPmxHHvIhA9EA/KJ/OooOnt3wbt
LEKd3a190wZY62nI17YovBDgsgJ1IsYFlhKbG3P/4Jz5/QPeItfpv/ewD6Cq
UB1qVFVUO8SKSGECesZaDxnEIbctdXnObKg5THBj+XX/dIGH7O/enxCJdGWK
7qGKrA20ILr/SlyEt43wla3s3LbksRLTjbdCyuhA4+R/2JPrAsZE/4uvhltL
uaCDCoy8k0Iob8+E0hsDKK1K9sBORZWWf/dPi0VBiJfDczuNxlNAlH20jQzG
D4lQ6+sraIQHT85fk4LwjU4gwPFZBVRSNz1ZrV9H/qBuTr4P/OCVCRZhS4dQ
CfkIw7YbB02kDlanwCpRdWnQJ8PFHKCsRhs54kGFDZcuqKqKaWa14q1BwkTa
vQc4xiRhceo5DcQP5sH8OZeU8IMgpRdTmPP+0EW3J2NdfP9k23Ipu/eXCLDN
lB6JYtDFhlXWZinKRl5JBfG2QYohwHmgPumlTeFDhLYUXPndP5OwBgxlEuzY
n0QJXDIrWRyG5qigkWW0eed/olekRY7ZsRkPmMM+hYggG4nnKK3VQ81L8RDV
5Yzw4q/MT7jU9UsomuFzWsgTyx5Bqrg4sRDPragElQ/EQEs+EZtlSlW6u+V8
z/eL5MeMKP8ZqocYAA7fWBksDChQJWMcutVAVn6StqkYlRivBM5ipVaHgqvK
J62WnfYmx2vgU4GrQjldzN/5MBxUktwajReeKTcxUMP8V6FA38m3K5UcJD8W
zFrx/IPYNceIDcezCbnzsBVs+2o0hF1M8o1xu5Q1uXQ0J3Qg8cCu1wb8EPlQ
ZW6Zw3qTTZBC8TmeObuZe8JEo0boneZQnUXX49bGFr/UDARaME2RRwinwBNK
6ZnBxKmA1GqUA1o0EhESsernEpz0C5n7ZB6jJXI8bLYuVyeYCVLhxmPWSF6g
t2oh07zKE2HGvqOh9q3fMDYWK7lpiv47xMWuw3Bficjks12ae3ryHb51PHk+
I7IBR2eWcw0SYxTankEa7n12m/4AdoXLPcNUZ7pHTbv/W7458vW/bqh82uVI
H/SHp69UzQyJQUND+d7KOQVZm1O1pD1X8UfxIMWFO0YneO1ktwd5dPwSbCUt
Ma9ErdRDtSM5QaS77RVJL6IxdlqzSx8w7K9GR/XDxQTfiVUaBNfhAk1ffU8A
gjkT4NH3KWr9r2hnW/1dDiuzc67ibNWiuyfg7ReERspMcEbCgxn7hr2QA+ri
24TCcz8qFDf08Yv+0QKpY7YHqGsBSalpqyF52hWctrK62Gx3GH61cyFcqtZJ
s+D2L4NcFQjr5Z1HpYMPhtG3snwWqSa9p9Bxy8faFWNWyrJd153sRo/j+2uC
+yZgiL8QrVONo3ivyHLcRMx0rqF0O3RaM8UQVe897zQZ4/bGBMF5NjPD4TEa
un6f3hMMQg1qbh26nHglulEW58rcO8PZW1eqpJob2/wGd4/3Q3xlX8cuyP4M
9ck6ypZ83pmzferYx5WYAFmYSd2KBDm78vF4B3j+aEVXr0c+BxcGkNlPs7Pj
dcI+k7RwdCS5yXvGzhyiIV5+AchqNn1aK9f6/8ONjnCfeUru3X7+cLIjyUMB
4BL2qtj79mMb6GDl6GQbjPsxMsdfiMM6jr57MJEIBX/cQ8txc+0xpE5kkLzS
n+6P7BfB7l/sUbw/o4Bynf68adpAJUctJP2F8BcaVQDeEZr8LffvPFe0MEH1
E/C4qflOZdWOBeO5/nAsLNXa5pMxp9qLhoE/KZ/1PSL5KshPtGluA8axscM/
MkbE/8WvUJGKKOWtP+6qLLG21VevWKbJCnqAjwrsHS0a848ux8kwZUI3BwGp
4iGrj8TiS4JfJRkNGcB4HNiVUmkGoZhsdkHvy6Ss0wFphEyR+rNBjy/OjDPG
fAo2QBMhjZYX2wt2UFNciSbc+vpftQE+FO899PeS3nUb76700aKEGV2x30gc
lKXMbOUi6v2hWKkaCHebk35zvnVq5jhYNkpEYXX34/RQ8uhaw8I/L8wSCL99
EI1HrO7cR+2ksvPz3GTl/WN0UoEeEtp0FcitutmHjydWfUP/MrPojA65YPTO
eBvJ7/qKoBRQKdxiuIEXC2uSxa3P0svApu6mplI9hbH1W/Zz/xvM++VuGaro
2hGUeNJ7xE2jICtthRQ4aUi5fAtx+5/vkfyTc8LEbC24XXBhk7z4dlOv5NjH
nC+pFjkEo8gPJySUUsVi3UUTfUswRrTyZvFQOOx4zf2PQhu4fTohZ7SQlkx3
XsR0lkBudo5NDt3IZrJvrK69wAUJdyedWRr0GZKbnxqxcup+TdtQb/UH0cv9
p1u+ia+TNXtfg8WFL0SLHXeY6H+P9WML8n3TMdULmV63znZoqaEfRR5T9lF4
pEkXzIPlEYW8C0c5RedBVFRp6GaUkmCe3g186QCUSYfFd325eAbHUf/yxcj6
65+bEafOOFMjmwcRpEWn5bx8TfqYWzMvjTNuOE7k5T6oKEHplRmOMDIVDx2w
1yZsH5KGt/xqbCi0XFZkkn0qzYdx3fqAcPDuQqVemHFAq9Xz5rNvNKlWJDyx
AIZJ9n8LsYp2YnbP/lAvUZSBQUaN94cK6XdbE4XvtUZmX40s4Wk8yysFpumG
6VTlmeCQMsRs88GtKrgzrlgdbm0Fj2WfiAFgp5aLjFPFgl1FFwZBXTOg6KL3
cO5eu2zLhwXBtFKXiPoI8yR6Q4/vdfSZQ9oaX4xNy6NV5VqPsUMYKQIoCIsc
s1fbewX9mzQ+UxqKNp+JX+Ph9uRFCvOjnlTQ/5H8D7JQdh1AIKIi2I9fClbo
O6qI+Jcg6GqlcUwiLbRdrepU+u9o5UhCKekLewgTjcBZMYfNcTSp4qWx1ZD8
p063s1VQunpC40lFUSXsi1voHON3mT23b0XA9BqNU372uVgxzJMpOAiZGZpL
vh5ZxbHoNCCSytJA02ww6vcJHWwuesWhheZJ12bxnXrtBmE496zwWL0B0Fj2
oa/TlCbpbeQ1qgJmj4vPNk3KyJA2UUOKTbD/mEnleJaGrdS14UkHy3yNjrGk
lTbIlif7zL9FubSdXLVYQGnWXKgpGLHv137yogtrHqnSz9cz/THE8o8bOWij
xfttmlej6XpFGdmYTw5e1GFYb6IM2fhRgWA4HV42gUG/GP4CKM+CmsKJ2s48
sNDeh148b4aMKwlC5L9pOLqt/EnIAd2u4Nrz0BjlEm6qldEVb8zJB49LLfAH
eMTX/5cEmK1RJuo7av6C/fHLuTisIoXV9WcLatWxGj6p0fm8ZnJiRGyaysKf
dvZI3W00CDxVaN8aIVjwXarW7c6kMBT8bxlR80iL6W0oHlA+bXuS8P3O8JwK
Xyf9gQkqzT6aWtKkHIEOSMtv4wPn8T3ZW7TPSNjf+hdBANlZaYqKct1Cg7eA
Qg9Ex81OqjHZyfAZA68VJOWGd39NgtSuCOhyns25z/URerHCwWshXYCjHVd+
AOA6kfGr6j4tG22NXQIIsalrly0r4BWnVMpFxIgl3clL5kdfnN8mchF6t0D/
YXmJEUi0k148qbRWDFCsdwOfLym4zPP71WT9fZLk9jZwXr0aKdMn8fYK4aaz
X2IYkYGzYt52fCh6LdSUvXCxn0A5U01d5+QvK1WpoUP2QB2yYy+fG94kIY4J
Hq3peOt9EFcglyM6wV89iFYEKmttkRX13qmsP2Eb8fVV5zVbHEdgF9P65Ws3
sQ4HmTwJAPFULrp54N4U9OW6QlEtc3a+gPFga3zcCjk3WO/oEmYEfXOLAzuU
NNHlJNq9OFncEVx3OJ0dk86V67AyimKiprw2xYAkfZCEsK1KHlQGARpWTOHh
JYL9RFEFkH4Z5mCT/tSzLFRNkMxwk9uK5ur8d2Y8nFod9e04eKsyFTFohpRK
Q4xCIv4GuXH3L6fkXfbtZQVFUICHCnRQSobdQ1tlad/LkgkxJzS6Oo/7RtwF
IfK443qT9rqmk8NGkDYhezUOlN4byawRnYZ6aei9Bqx87HjFU8lbTypNjOmQ
DZwy6TN10XMOA6BtkoZwTP7dNMj2xQmX8D5Ovy9u/qIOdQp9ETvxw6WVXg/p
LH8Ndz6+ctM03j36gtFiCdxZOp0ddmvMubs6Rp3/qm9hpGWkx9esMYURUROo
7A+FzmTXEkS8x+qXarzRyZVCT7ThoeQPn6ZXUVwv115A4sc0vgJW+8V5tdCe
bR5L5LFN8w34eUJhxs2d4e+4rVuGChB1MuAsavRQ20/fL/Xe/Q6R/XsEyNop
SGuzMPHjs/lAncCTLWCTu6wrFe/wjQ8Do0CUFWX+PkvP91aKr2gNgfvqo26Z
Mm+eaoCxgyoJ32keSgiPB8zkK+DRX9h2hNyOkBKZ4fvopv9GJYxszaOO6eWz
rkX+c00Ifd2eY2lZGIfrXW0FX+oVwwD/Z/S0hplta51Uj80kNQVZGBDn4eX0
0cRFZm5BlYKK3ONjDKZONSxSPJqHVA2AlcrC1kh7+4nq6Uo2JUbHAEBkvz6R
DJImqEckciVH+n907mZzqW9FW8X5MlLI9n2vair/biVpKusAXTaxw7ghWUI5
iKUuAlw60r8zxWSIilu6lf7jfd8lUIPtL5r17jSfENvAvlySd/1zNbim8fRG
2QTGaBuw4VKeFpEiEOzFO759Dd4tY9J8PahYJ0/pZDY6h3RXqlPvkbhw2BJO
U5XCAteUsnwzdEowLi/jj0q6BAPN7xze6ufDdrk9qzEwMyGSWjB4t8LEZC5X
mBuTxOb9TUEfcQDEgr3qyQ5vwudbxWkv1KvOzxKXN/I0klRmGi6DWQMjyOid
hZ5fe80aZcnvXz2HsksBUjaJg7Y3qlTA3eiaYJjNgXegaZ0ii6UjhRUduCSp
+lC5g8BgFs3/r20uOXlnQIiVWeWtcqexBbfDVCKlkxZfJpX6kdqsgFiqXej6
skCZGK87HmzqoXJfcjgcZFMMP9k44ZhJfUibsjlr7z7c9RZOk+3cN/z59VKI
yYS2KLts/c09/vT7HI71d5qxbriY/7bhX/HUYiDFzFo5JG9QzZu88vkmlgds
KNXZHWILT9594JGP/HdnB53lct4ZJXlv3L4/oREw+0twuCe1ac2Lx25UccXK
Oc+0TQvyRx4g5dSNf/cTqAJ6FyZsyWQmEGwqsv9GLXiykLQn4SWG0fIzTRtR
UEyieyll457oCOoaFm7z9samEZzteMNZPfF8Pkc3fLesDfqQXfjOC4Y1YQEA
+orrLCdL3CnFnDXczECjxDf49aPWBQmrzJNNZ+AzfXvBWkNWHnNtk8leOdkV
iz4n4yoLosp3rH5Uqc6RgUh8pjUkopjlZpOZmXyP8r0zZjQDAknXCIn2y2RO
rLxL3rkQTMKzP80SXQLgbQoSIriVaP5ANYlPf8euX3mmz1Mn0g5wprvX4M7P
RRgncr+ArVUo1hHXNwt3gTwUpPtjQ3ilZF0gbc1iHy6/mojnCJIPrhngyi+w
ZkAJVmd7KCfBOk/pP1LbPcyUTQ1KNSNsgDQYKQsMBqdMv30apAg7H2hTnR79
ldKq77j21M8anpjOMKWabl6hpQ6PIwql50T2o+LpVBhqcTg2ad5oJUUem7kl
J5ZDsmwyLd7osjBemRrc57PDL14JCTGvAvJlhRCQ8DwQQBmC8osq2ZFT08RU
4qEEYhXFEvyFgH4p/jtTfL0EXitx9Ey+Y9T3p3WZ0KZgAgY/tB9UV4iJ1hra
uWFm3ycmUrIhCVWY5uvakEHg3GVaH028QLz7rySnW+tgRFN0ud0Z300GTHt4
ptIvGIQzeWg2rqFVLl7a208SpfI+DoQz3Zz9lW/cvq0F57QXHAwvyNZZvMiY
sMnyuCfRmRZHgzB3IlbKVK/dnsTiqHsqp0WbrQHHEcK6I1OEnnweYtzEpDGQ
tYw6T/ml7O1Rd5KD2A59ptuMo02NvCXhvJ/qS9RcHzKY8wVRAusoieZOczNZ
8Jo745g5GBdIxeRpOgIUbZiyZUUa3aWALpxwSGRx67P0XNtYXSB1rjoLe9IM
9IMKK347gf6ytyxTodKx2gx/TW9prOXd3eFxrcyu27uTpF7+LFMp3TChAb5k
Hhsy1Bf2xOTahdtt91RfXI6guIWso6J7NG/0dE4vTIfK21VDRK0OzAe4nTgz
efCv8BAe32zjdOHkR6l4O14bsmyNl78u//MS1VcNNxJ3iWtbMdok5zf1QAv9
GXfr8JWdT5MnI+nG00La91Ork+V0yIB/MqFla+mZ0iZ9xpSFLYJaH6dg873b
EVlpYxyFCOSisIToS2B9p2S4BOmVZ9EAq0BcaYPzDddex+Sf0csUs+4irtCz
WENZ2blcZ4/jaawiZq7xSo2A0Bxm6CAqgLDp8wGlRndz1D2GuPD4prqhUYp6
ds8FMIVNe47ud1vwFY1nB9wkd7wxC1tKbvv8lhH9TTVS+RzXKAn/ksU8GNkF
UcSfATYby0d0+UXCItUHppke/oO4x4SIhH+pFSLHhN+0OKeEQioZAOwYRz1+
ryfj/PQVWVnx6f9iD7ZXeV48zWPj4Cbd7SI5PKIJJGYhr3qrmxzAU4n//d9g
PINgTyHW15JoOKAipoiY8k+UbLS5lzZMiiRNWDsTzfD7OFpwtqfKJszMOV0B
2lFrvMFdljC3+lS0RVpdAxsCAGCiK+Lpbfiuq1DxDsyMZqphs7ngoaTh1hHh
Wfsfit/NDJutUHTe6hiaps40qwWKjeKGfdSQsAtFl40maIfrN4G9JODgZ/c9
MlcyqEWQtofZYxDzO1w8mqr5qD+e0Yp27yRD4yWcD6qqkYq8PSvGMmRt0OmN
7DNcgEsC7jlA0DGxSc3SbhnAJBofS+DqixlGvYWT1LYvavF2WNJIU8KjwlCN
DoSoHmZ1qlqK5D2a1JLCscgSyJubzYQah9m+eeo4MOAmGk3ZhNAz3iI9erOF
n9xcEZCyRdA+ZcQN0irZydz+ltYgqdIwTMgcFpuzeyMUS4WaYSWWMv9po2v3
p+gfv2uTR9P3dOyg86GMDVVs6TbRYqnj6h89jYA7TVI0hn2qxIVhF0vdTOoT
1LxGTQpGzFvK8nKJ2l3KVjd2UH2J4CWwxpOBAKXxoS7SBwJpMb8w/iw5Yw43
FYOpinNmsA5n3n58iAC/3Wx/pwwomkwa0Q2j2Mq7MPcqGte9pHc9y4Gl6CvX
Y/Csjmpxxg7Jn0cM9MslafstnnD2P2o6Z9c0C4SctrpvyszuB9UoNjkaPJaN
F8bCsBqMf2CFcle8CtfiGzJpcEIfA8dxG4tjxzAKlLd+Ehf8pw9K9F3/sHlL
rpwKPi0X9rPt8yu2/V/Zd8LSaSIsWSBJC2UvDCo/iIU/iawENTzsT7krJ8L3
y+irFWXOu8i9HdJC+1bP/ZcR/VpuYBQ7V8OJvOI5IzVBj3ub0FvywTS31Xa4
GnYkwAyWNcd4dfJhaw4HARZa6vUFblELMIKB8Cd/WL7d2Rpyw6AGtE/iIyiY
v0GoNKMs5fVz7cFnryMmOvyM7uujF8QDqRIh3qA2A+na26uVROlaxGlC5Qf+
QvQSb4zi7z+svAGDGhG5uzoJJ/nfXDE3tDWDkeWL2c0SI8HSg32ogs22ioHi
/9E8kB8cTuykTyoWqg+AIBlzEJn8/ygf02UlKpexmcgK2VbUw/gzoi1Xu0ir
7J+TgL6kTPJpKPMVGsP/WhAzBxFHRXDcSChDcyTt8p6oXFyJqGMX3/ypnFq4
eBvE0Apf50Eq146gj7ivJDgle5mK/8+xXaF/3qMC7eP1JvLpTOrSu+4SmQtb
m3R6E1E5uscbJfVPeTWej4NAP6RbvaIkEw7q8iuAmJHsD2E26zr2ty+AJ9SF
oCRL+lZzoedgi65gw6qw7LjnK+2B+quJQVKra07DeZJ0T6pjKFTJyQIYHXB5
4hswizXtRtoczraYpj3sInNrUHdVte+qIA0S5mQ2FsBSwyQNZ0EE+jnvDuce
iH10utm4y3Zrakyc0TE5YzpJmThX6gXH4HwNBXhHgDoWicurBHbuAgTWcY/L
wppj4kvGbt0Ui7te4Ur/8yGgGey/drGDu+JVy/E70s6l6qJrNTuitsk05qF+
Ga2cKZml4ts9gXwVKc6ibrkj4c+vJq3zDli7UUfXKF999N65/0lV92IIkqY0
gLe7n03MQTDd/96hyUlma2n9VONZW8WAmIhhM0Fen71CDrbFUOBdK4X2tWy2
ymJXZKfeBSZC4ffN7fubF6tSVeO8PFhRqxabb5jBzx8qd5WijvM9HK5X3y50
lkI/csTJEdH0BOI8YN56GNMohz65QFqoUz8ByjU0BCXZ0zgqbUV/k9RyKUb2
1GhutLX6QwLyOZ3y1FXSHbxXYOQK+/EKqsyyMnoR/Bzz6HwkpHWmXJyTI/+a
kIhSUOI3jjYQYFNT8DLwTqd+9gPzuFTun/saUzrBPWmZBg/CnDe6weaLbSI1
jFIYJ8DtxNcdUlMdEy/qkiLvN07rPI6zIS9whlwGFMCvw4YEYhJ6g21iugQp
hEEEP297bWeJYvuq/WBY6MC17iuJbThEN9c68NRpJs9/mlD9yBoPi2/0Fk3G
sdL96LO5pnm5eN3hLJM4+O0ucdxZO7Wi1fY8DuNng09SNRs64QGJl5hoAAEs
ZFPQoh5uzM5bSD4ltPjzIQ8/afgV4eFgyi3IHGA+gRBbfVGrEby8aE8cTu2t
G6aeYxS8mwtEn9102TzsVEiQ15eeotjaCi8QXJif/eb1b3S7UzCko/FYZ+Um
/OBR9u3hyJxDOFQmHxGiKQM/FgHmR9FAAr6TnoykC8QM4I0glaSed6yD8qx5
Edvo7n17INNa+ZXcSmfonYnsJlBmX1uaojsEznUmJlxj58YtTNIc4xeBNOZb
CWeChZ5AH0XnhfvONU2eUUzgi6hc5jxRtRJKhVup+GazIyj3HtF04wUd3Snq
D0Io9/mdPqHXJ7WPkO4knQQLE8sLQigFOedAOEObM1a7AXwnvVk9F84OkfJu
DOpOSXBN3q8hx2jeIfkR3jt69padcqQQk9ZhCB4igZgi/FLES3FLap/BoxH2
TQy1HUQ1locYiCWbfxGmPaQkW6HInxBwzyGxhjjxd69j4ChoGaJUoPr4Hok8
YH+2tL660PIeW1hTkubLGezhk24r2Bd7LWpkRV3XX94WJfFWDUUMQj2EdJSx
5hGoox3cDij9/5/C54IOyXTvEfCcYGJGhczJ9N3nV2xjpy/wE18fS9iBKQsD
skIYO26sbHMNm+nzPheoS1r+KHYOLtl4ykK2LWiYP65l4SatK4S6YB7QGl2z
F5YP2903BIHham6FJgu6mazWkRrz5dcvyLx7NFNwl7+ivAeAGGZy6/jIoYFm
spBEj5mcxsEP8yu/CGC7VuSs/0n/GT2+0YQem5NO+2OBUCAvxhMuSfKFCylx
D/wxpmmVhaDL5wqJlesuvET0hfmEm/+Ql61Dhiwr1/Q6dUbG88XN8A8tZOg5
4EagExRVv3Yi5HGoX6xHW+KusDweFXflAmxKzuk7x+v9zLmsh0ccrRjQSMaV
KcqNZADvLgPBzHxLi5v5KMN40uCpH5zn8D2Z2sPMFNWYJLC41NMM3wKX7DSI
ArNb38Jr1S1kbGlIPilFvJ5KYQwTKMle/6wCXeEBELJ7tkhmadI6M9L/fXeG
QilWkhbz0d7GVWev1KSGXZgQ/8c9Q/GukxojHUCAIRWvdO0rrhMQnWfwafvK
RO5EDVM7Z/3iUqavg9onGhnP6cS6kT65IMj4WaEqO3siYxI66nobdzg56BRT
glyGj4v8l7YWjAu/bcprZCX43XlsXKmCepYmcF6vGd5X8KL/eswxmgt9QGSI
wZVR9Dk/iirIPOdF6k9U7HZWuOyzz8V5xtfFQ7NH40cRJifH904AeHNeuYRR
2PVU8UFloiCfqjrMY+Idc58ab82tlFM+XvAYkay33BL7zOesQlYNMOWkvMxi
iYixTRQvSUigkqu4rqhg2JyVpx/F5SGy47pZhGEgVkfAsflLTfFwICbgACDn
i6gIBSb9Ozf7fRaDIfynPZ1Mb1GeijCyjrrCx3Z9/BNcUCcr+igPvT3x/A71
8AJG80DtteH6atRXB7cuE00/UFza5W5R4pUOjP6VMNFm5v22AhEp2FbEBX7Z
nvC04ACxynscmrv2XYI6W4K0XfVIFKAp65oYs+PxwSb3M9RrivIGB6ouxjb/
qbRMWWgwmrJDAYG+qhdFPqWjOZeYZ7XbSf4mADvf8p9GmT/9HYNLtjF3zLgc
G3UO9qX7AqoJ+TKew3M/W2pPoMwjOkum0zNfSoet32xSTvHrsxukG4NmnQCL
HRaAc9YTtT1dKMY+CK65yAAwCZYNRn5A0mMvVOdJIz9Qof4/gUX6OCFHvSSE
HMLQ9GDdKncWSZ+cBGjD1eHufI63w+nybDgTUcG6Y37AzJ4YxGRXzrkm5k3u
DozJWAqgVIyR5Kvd6mBQZeyV/obkgruY5bO7AWGejMuE8zaYVjNVxTX7zarw
iflBHdp2VOiUrxdADrkwjUv2No+Dq7/QcR6VBPZ0DzAQubhL2Hvd2RDZg9+T
42cjgTy1eSTgUlCBpcA883a0PG/zF+vIjnHJo/AErCULQSFGNOmYFWRVdIYe
vgmqRaoVLlMZdbsesKfQzuERr9aRgn9Z04+OyugcnZnFaLOd9Fmkd42icQ56
00oubX41BqFPCxiDVJRqcbealMRis374h9YV1FwzAoibENBsJBlK5QE/mHp/
jZnW+SiHwU6TPHElc7Rq/V6Nhdm2efTzfCkOVaqH/EODn67rgYi6c1plj4/C
/V/+P9a+5uQkv7dFRGK5aPWtLzePhqf8T6DFst+j7Bz04cagVpvHvdmBaC0i
asMctozD6fqKNF7qey7wsevh69oJVfVm5Iun/7uTNodbWi5itGOzC5f+tt12
mYX0KhiSoaqu+7c8aBXpkxwL5/RAyybDSbiABzz8ZTcJWCtC3SbVe/t8Iw0X
sYoVajDXFQVDFtkKt2GsaffEc7EB2FN5RMugDu2uVhcwNt9JIQUsAYccqqlD
3ZM3eutabaXL/MvfJ8TDRX2/0bzmBSe0Y1Dk48BfF1i0MpNZ+B43yR0eyuAG
vmI01ZNwbVtUHbtQyEOQnhdj8V+W+fNMlTLdJikyhtAc1VGCqfUwKJUqdCA4
1Z3lRvj9bNtFSwohzd/A/zWw9as+WzIgaFbV+BhLXSRq5bclQvK6kL1gahIu
B0LFcsoNcyIID0pTIwURWkrMbdR5vRwlzPNTMOMVoFgd8GczTvkYX7+AcNUY
C9Mf7W8lpR3hYAUwVaXlqbARmKbhzUIWONkkjBdgpy6xB4b0FHJQBBOsZfFX
UWlGd7fy4pB9vousMjU9Ux37mVKZBjVp6I22qngBwetS7TUWTI/t6rdXNmDb
iK81WXvL3gCLQ3NfucxVAMGfJxxGGcXou0Zcsoibkx85JO9zLR8W43n2JeNb
X79G61FEVdOmc7TbUxuXcuoVUf00W3N8G3qNkP05Pe7QVvMuqvWK3Z9nfIr7
qStqFia8SFP7JEZGZx1aUa8sVveIsmRqVUn2gcBFzqMEFcO+myeJ3z3DZFlo
Nn18XMen3qZPdXakAanigzsoMniLbricupuDTTpcmr6yXQ6O0c23WRFErSUC
/QHQst6k3GdgosMUHMoTW0cSkIvJ6PImmXvM8+7tp0S4x2CjHp2mQFvOzWXZ
Lypdz6kP0z+wWqLKB60LuUwRWGAw8flv4sR3TjFonqLpQcVxhIyPNfu2+KEK
88tC9UtGc5bBqUoV5co57rrLOBDWWOmBCgsc9sMXygEUMGQizttMekSf6hN8
w9xkeIrNvj+oLyl7mV0Bl9+MRBAoJWytAPnCg39yRzPKJDNWugkB0YrqVdPc
TSTaZU5MqwqCq3b+iBkJErZzH/cNUKZVJp0xVnjg1c4gv+VyG+wAfxxSK45V
4N4T0nepCDdHrXqEPjsGXdlZ8kMkf2Xm8CpAqJ59yIvm60ED+7Kcw1QpHQas
Vly7uLyjw23VZ25qdKAVbHgD4r2n1xAdpOVFP/LJchCiVtdaI493/aaS7Pfh
+p4CNTvr7EI7blhW2cDVtHOEYh8PFTDIb/ldQmSIHyXZF5SVvDQMo7ZVHgsw
g7CP6GkNb7vOar8LlYtw+VP2Z36TpSWVGwrPM5tDnJOpIodqPPdxVdqvlFb8
y7WlWg3saX2Im84h5NuuSxj4F83bEHCbdclSlfhb1NtiWHSjR5IcwrYL+0jO
4bEj+bEJ+zYchf76xvlpweoyJBuXYyXOTOMw24DGXsnAvIJdDL7e5cTX3uvr
ZdPL/Fo38d86HICQa8Htzn33lsdG8AtmRRVRUpe2MV+7DsrMbI5N7WubtCoE
+4LSmlsCcfKPbW5crZVEyqdwLyU4pkMc8VTrATNkyYHZHhKf369BVTc1I+H1
u+42Tkupw45CwtzhY6/zQfMyhsrcXKk25tF/Ms2lgIiA2qJ28eJq78ut18Kl
RJ9cEjxg7jA+UGQHBaw1VAOEsSE+/hYSKpCLQffAZ51OLee4NsAycOvDZ2pD
KUwaYprIVKvEQ4/eRYmpqXuy1adg6ISvNx9EAW6pFBEpq80vyzI2c3jjQEOL
L8lvyCHWA5BC0YelnWynLEflJsnd7wxNLg4fryPmV1I7x+0ikgDTE5L0QBot
oUHwRe0zyU7bOfBlclqIIJPNIp4HTsUqSYsxffKLSeJkmoARVXh2nQva0sYE
+qbXHD/y/uQvorbQysyGHj6Dh7DkudxjIIG0G8YK6z2chKwcexfeUc68Jm7c
9GOkjw1KFYTDG1Nk+dp3f6ehKKRTuc4x/K1Hz4T0eCtGjGMCTTgkaa/S3yPW
7FjWFkZqJciGhiJZIce7CJbHZAPyHiEg7yIqbhEp16hZLutdJOoN9K2ouYQO
tctW9ho+O5ngAaXbIL7vyNQySiFxnVQqLsyCoxh+i+qX0tmud6DdlcKNDMLY
mTkJtPzDJ9viZEy7SOo7nndc0CgtwadVMNZipoIZOs8G0QkiFuUzOAqNbcBn
x9SDi7dWEBUxfPcoQu/UxQZ+efD7w43e0pk9CC4hVu/fkqtZ8GjGPQYvDHuw
TkteSJ3msbtYaICUCpryICt/dvA4uIq7vbNT21YygBpPtpSStoLqAjiLeZWY
L8oUQCkdsn1yd0AcFie1PBKTMfVj8o4aaGT6sXwJPOdptXgYHN7NyAc+M8Uh
+rhnJxLRNtnEVUpo8h7GCiC0eWR08rRO/8IVjq95jb7+n9bThON7/ebn6RTz
wUhzaS5wUZj/Gljzjwj5TqlnfSbaqVfmr75Ah9QIG+llW7d7Gw8RmyRIxEGz
ie5CVXsFh9lQ3wVsJIcDR+xhxauTMjW+Pnxlrr3FeE7Ln3vX4lFsgFGFOjWC
Po9a5zSmSZ92jvgPoMRwparK4hPsdvrppOXzUBJA9bYewqqWnjCT6eBuyMW4
RZ8L9PobACHrW8L3AQUcs4b7NyMjXIzD5I5yGRMOfBagJRRjc/TtHiUL7j4s
DmkhUsWo7TA7xF4X4Kv9CimvNqW5moo2PDW04vRsUWV0zrAvClYGQC7CnN59
6c+IsbZiXJL4bfTMr1wuTrvT23pCJsYX08opTIEsWBdN571csz95l69apnnn
4yw5ZmZp+B5mpj4zUqBNBenpNTPL+x6qdekRGWfzO6JbqZuPBR0yHO5jpgKj
vpvu0xmJH8Km2xMnXmlXMnSwZRm9giQcAcijPlgLmcb5IHelw3XUyEgZuVNw
NAx13A9JJoyhanwr9WFqGGP9KaxanxjrpVwX3bT0zJJDSC9ZrjQOob6XM012
+Zi7eDtORv3zIBhKTeUIBflezkv3v0BM5CXEo75QOKV5RJmJdqSFGU2yJu/u
7V7/uY6tZ6TZFzeC+r82JHY702XsKS8I2HWBXlp8Bw4xwlW8fBrGUQ8adpCG
Wm9n5w+LcJA7d2ogccgRRzvfjaP/f4k+H91Qzy3xWBOYKNug1J8MtqdRafws
VluCMxMYWG5IFTZpMtW66zbdhoY3ILrzgskMCTrEbQe/L18rUH19AUuPk1Tn
UJ1inI07xwFDY5pPZc6A08blWfU0z4M0klghSwWCx3rRouZ+R+mdzYkkNQ+s
jBokL1D5KTeDDhW2CGD9teEP39bxRgC7jiRJHUOvlILqLbhqfr9vdQah/Tjg
pmjxNPQc5GhHty1NENSUwmjPdpFHeEnRPJ+U2pSKosEFpLvPa6tslAUk5Xce
klheFKFtr4Ovx3pKpAWzaklQy88DcDxpjg5vfyKjaT+2+QcgM+FtsZ87JhiW
fIXPxjqxQ4h001PAsqggE4c4nyJ+GBn5CJmf7HU4+j+T+6n2KZkNvjquy/7G
mxYylFkRMYRuZtDKTNLC0zNW/BneAVofhrS1FwBHPjQrvoJ7ZMH8xl2A7HU+
A3zRpCatdDe5ezMAu+fWFMlPk9w6lt/53pFjmdwYfSvSbOtNj0Jyd+HcbnS/
CbKNqNKjy+aqBCPi1dsorjhudgNLv+6bxZLR5erp9N+xJvFnbNYnzbCRG6jU
ONtNTQ6+2NzvYGX8GvLlG5DxfL50XllDkbFcl9kebe1vye4Q3IvS6tBPxUzz
kmx25+VcOPPLO6QXqkIAoPLEPux/cVwBq6ivm/K9l9NsJ7NYl5dqgd35coyA
/sS3HmCm8phrsK+bgwHnaQjBrWgT4/IwpgIvcU3JHmDqOsVO0/bsvMb04NT1
PmmT54VvnWCTD9KZxRJyG/JaJ2kQ6e2rcEZmpyfsOWQmeQOgtnt8S/LLnwXJ
waAPlQAUmWFzP179d2YX9AN9XUsGPyl+qGMYSeqqWSXmBjUYOUvwiZ60dtpH
d0IuB0O97EsI7zCZogsQdfgpwMjkjCvP/nUY1W2OAbuiYOlQiMJT84BAGYnE
OcRoBhklsX5NdxurGXJXLIwFLCegbXJk2i4twyuURbJu9/6Fi0P+oo4LCbga
tzcnzOqWfE5yMAnXF3jdnjaVuwaCpzJX9h8texkHb7UBfWCpHJ4lpvTQo4hZ
0PaDqL9asLFp2G4A2iN5uxOU9dQWQe4/zmJ9rFWCQ8yuy3UhA3NeCxw3RpRF
ED9wQdNJR2PyofOG96SOgI9r6JUBJpBYf6u+6pifC6kXfrlOfbrEMvDS6xNd
USi1iWCETwv+0hToaNNDhieGENO/HnCcJKIbZbOvrfFpCGoWvXgU++DAKBdi
IXGVCFgH4WnZgv1Kjdjwimbt+JpkPundXhWYwx6tuQ1JLgYfFxUgTB6sL0EC
HT0jPvvfwRgwyn95amTZ0fH3TdkxBB5OY+rRurTCRWz40iG8OROZpOeIQ1bm
OU96wE6PjDKKXYwhOesE9VP+pBzaI1h/f10jS3atpMX85hBl8fnwI+8ONapW
zASakvd7cM0vWLgegJWHraPCxWCbafIMf1W8xi0dOGcxkC3uJUpqJOnlvd/z
ZolFBr1Ji5I3ebaBVCQqQVo8xTjG+F7DYiSX7q8aIpSuXU29lsJd3r5wwLBG
8RoYcTPl/PMBldLLjt107ODkC6ew14WOviXL4R/EKClKC93LzWJMSlikeqTH
MLH5Nj9AEMpFvjeAkEQyWRriHQOAGfZYqF4VzUJFjxdF2CJaS/5epszOfce6
PwP/YhVvk12epcDf4M2lCy4bpWahFx3Av8fEz+7imoHof0RFWDLYyz020iIr
NmhA/N3xBca29oCKgzNaqA936UNXddHsjn+eVP5e5d+DwkE+eUTlmjrfDn9u
fYdQtUjucHTTLST7Xo2JUE0yILSXU0l4dY5A9RtpRvVDI7VeKIX4AZJQCBGf
17Ry1E0tgVOCbE0L1J56LL8apLWfZmQ9XtAhY1sQjuzXPkWKFGG2e1jFScvI
cORfskrQCXNPxmsF4eY7NNdfptoloxBGr5u5D+2CZpcp68li9KdJu+8s+AvL
5aGsSEb3NisGhOwUTuwilOX9WFTbBW2MtRqm0FRU0ZWDEfuz0nqM1Y930p9e
dKBlV8uycBD6fCXRjL1QFYhAIKcqbM0gLdErT5RYsI6t8SccJ3u4uYXY+UHY
SXFrV6iaiL5Q2EzItf45B3qrlAXOC/zh8X+KL1szK5qhfwgCu/CjD8KtsPDb
EHOsgFpW2+dvs4yn/i2yDXF/pypZm7K7li03NImU8JyOpz9EKVolYnYgfYTm
J6biOykj/gq7jtoaPB5vX0nQW+8+vKZ6DKGBvAqNBL2RCXs2r1s7Gs/PioV/
xErkfoifS8bz+hCdboPcakCAC7ZuHQF69eyEENZrlU/yHB2GpUFEHu4N0mnO
e3oeVQl1erNOL4eVgt+MbKQdMfM/Q/QhX5XXtPGqOtpHV7mvo9ZS0n/dslU3
UWjYVrXme1kke2iZjoY9ytCNc17U+gPLbhUnCG4BnX0G5JS1BkjUTtv710Mr
vP757XrNqpyM5ntkl0Qzsi9utdwhD4o0dfit9gZJ0zzod3MQ52s1li9Ho91d
keZO85CV0w4HT1776KUZbrgn6GysBdvFp/fREh4AMQ3d5BNYQeNjPFj3zmMO
oB/cgpxqVc3AivwPZV4bBJlQ1moyRqIvDXe4I+washCCMW6q1Dp0HmMU6AGW
HHAnNR93GDgqqBtvbQLi9bqRhfHSGJbVYUKJhyg32ns7HcAyO+rojdZVe1Is
1a1Y91oWwT4b1Kh2e270Ynw0lsrIzN7BfeXMaoTYz9JOXoGfeFVZbEsbqRsN
p604QKEytNZYPEI7Edv16JvfngCzQeHxczrVLKq04xgpzDp7O4ZJrpjEr5eH
z8Y+8n4GfOe2CW8jDAjvOuKOodhJesl0LOdP78YPUNmdsnaTYvJn+yBB5dE5
V5p9oH/cLyVKGKJVb3n+m9tJPBgT0yFbQeFxJlljHaqL1iQsKjmhQtPlKz2R
oaWtmHaPXqL2Bv4qv8pkEUVxDwoT2fNzW4pLmS/wq6zXwiz/Udz4+OgAOQcN
jf4IhAUfnGf1cgxEAxUKoRbN0ZH6xYMQ/joz3nbPmHN2GXpDZ/TblqsT+nTB
N8zZl7jnMlIfnyQn38xLP09CYIXiSLfcjxSP5iERfllmV22BbDdm/3Ik44cY
4b/hBYvij1KdX7VQTZXdBBCs9LaI8WofMhwH7/98l65jKLL72UMNegPewmyv
jLqStIaunzkQvD3zY6+gyveA+sDuJbn2P4OkhhAyvMMdMqVmw1q5clapyQL9
Siz2KftCvpKbIkpej4CYGoKSjlsP8VMXsYSnObgiOk8w9Y0rJTScNCqpRppu
XHsF60jwTu3pwrRATF/Yec1rDL1RjtIxS/aqn3jrJkt/RTIpSMjNUzfO18NY
HkoSSzrDWEtyOPGSmC71HTGjo5d9ZqemPrFB0B0K8X4vclDit45ZzEZiGRYS
Wh/3VP4q52zcUl+RzxcP8MFjUQqigQEuIOvYWih6Y+nx5xM0UHPoqdzI7Yyb
hr6zIIetMEk2CxU65EtkElqxAzdYz/wWpE26XOjlYROjnLZfDB1e72VzQUND
BBRq+GrflSpY3/4iSkjt8lafQ4pUtbRGuTCxUXOfNGSOrDQRMemrfZ3UBkYn
fEpGk0nmFZPKBFBqDhRvbVJWoVNdACD4b2d/4L6AbITZVIZSzPy5pijkB4En
uNrL1L472o4iN+YkOFlaVGaWQSx1whU5RcbgD7I4y3Zaepe8NOMiY7Nnc798
8kSakvIrRQQ65AiWxRKVyOxJpp/5S80uHMiJhACV/Y6QRmTqq6MOriuU+vrE
o7nNBkNzq72OoS/DRxJbF71mkkNGkq0b+YhU3zLnXRORNgWrVlHD6iasrqTo
YNyidbA0HZ0N4bXJuhQFT4hKcwwuyjWhd4u6c+nqV5LgaPXF3gVA8FS712p/
FnM0KzUbtGX1kQwM9+E6J+RNnb7nRCSy9FcriIiTaS769XrjA8S+WeY7WTPh
9DGBvcKLraHq45vPD47ahpAJvIJcW63oz9goMBVylFhEr3CYdkWjwRgvCw1h
G59PJ7LAqfoquqbNuUcH1khEbL1FoongVGX+WZSoSVEaywKMrlRzPzxrD142
WfSSKmqhQH70+cBnsrePr4M9nK/IvxdtCfMzYalf6eDZzZuw2QFH3Cnak54G
rxXwq73s8L3+yDgow7sjPR0vgbgsuLwlgXlz3uxaqHMoqQ7TcROFAY6ZHf8Y
JP+E+zT5h76oT6O4svfkiUOV9kDmIlf5AmuVy0Kl3SPeRkN5zzWyZMJW6ZUf
QBpXJlEjLrK6Oyq1J/6oo8yxN6FjftiILw3h8yRQNeA+uzuQeglf+RvJhxJZ
Qwr65DYZ1HAIn43r8lpZZ7nNQQTnNGPEir0ED392E2J5CMnxSnSqMM2gHp3/
m8iSGPPw2eYkXif/s+CanKEXi1bxshvPbAbb8SNc6sqOQc0RsuYG9CEi6eVa
4AL15od09pa2qwm1xwb7v6OBsABr6DCohjKGKqlhq9u1H9Mc5N+2BnTevf2v
EjLGkb1bMyNzntuofB8Gufv6Ik+7LoBnsy7+z05ZXilQlN17/XowHt24E2vg
khRUXfXczXDQwjitsiGsPOil8wk8/mKu5VgBK8ECg9fnguA0s9cAfiynoq34
N66WMIv144c5+uZYMgq07t83VksCfPtsrwGMNYy+WE1ncjo+IARDHz4jbtkf
jnY2pT37zKoS+t2VycETTrqs9O3dbjAWf2ztpOkCsL4+9LjeJo0CLieMdJCi
C1mtj76+iYjHPKJ6OuB5n9y2ssRzDgSafeFnk0qgCrpMYdG5PquOp4MWCq2D
2NTMkyKz/IbRG6fFwM/67W+o5xmfrirkuNU1aZPZ/nw40AzpiAuYu5G9iEMF
N78trz1c3GEjuSy7yCyl2nHfV91HXuZkctx0R6pDK5eiZv6lyUaRBz2N0dUk
6ZY518pkcjSHO7q2BYSunOnRVpp2J47wIh4oi25o6T7VBAlVMUwYLVmlEuE2
KmWiU5krxWN7PaTYwvb9D9jcxySRCFxZSk8Qy1F3iVxSJ3QO5rzFEE7+AjBJ
iWAU5Vaycf0yXNHi3VNrC8TQAl6FHL38Ez7GB54C9TwhJRRt+ABkMQmihAYn
3h9nUqus9ltX3f/+LR29uFrWXAOxlc+92u1qxiAfkz3js/o6OxZD79BGZ3HC
bu6IjZlEC6TwLRmLv/sZfJrczI0Re7CevmnxLF1JsSfJzMowEEqcQeqk9QNN
vs1lSTsik4ilj+uKtx1amCEpRLv/ox6FxJ9lhXs0zaXqSIZmWFwZxEzm4Op9
0MTiClGFXzzQAjoOFL/1y28PU3GfOU6EDNxRUbWjM5i8FZyUC+9nQ1p3T+Cl
bM0PbHF4y1VKOKuvFcKMfXyUGqS/xch7F8wVE4fAo6V1zVKtLWFx6N+tQU/v
4yI/Og9TVjIxZLaHEdSwOXseZwc51KA8SQ/GQ4cNQ3/cP6X2lTWJTTXH8yMM
V5HyY5Jr24z3lvYkW120LYkYYTFqODAYnQoYouloMFFA1vuBZxV5/I1fv0PY
jEgBHBxMMC2XXK8LB98rwPWjdjPCqPqQzto4kwwgTnBm9mi5aGDuavzkPMBW
ZSXkEa8To/P6BMo/PkSZ5nAfHbGA/GNO4AxN6mVBAa2rBsswP6n0ilIJhNVH
t3r6kDkxNIBK3jbSwPS6OS53DjBqs81wBuRke2+LyxC9yH6XKQOM3N+bG4c2
2reVV1kjvWKorzCSGxn5R97tNOQq/yJ5nwKqA2wANyugZ83q7CDvzY4QTJgI
X6WZBnslYTqyUIvVkRoUcpJaglTq7ZXZDKxd6cHlDJmurLEWgZwVztBXfN1U
mP1CbZ/YS9lidmeFm68ukpAOFkA4zKII/BGjoB/gB0+cZyjP0h/t1zCkZObA
IoddkGA42V4SvrrPkliIe2ljk9LNBUhvU069Ab8W3wa3RSaG5FNqk1/GZ3f9
7Sk9QpT1RWmEcQr1uCBYljDmyxX6/wWERefnOAWQHY6bsOy/dodwcUnCZfqM
MFuZAuDWczedg/E4zpQte52hoFqZAa8J2PyO6GmwGq3tL5HK3+Ai03XoJHiu
fDMxA0mLYB7Pl22PvlsBkJLT9GSqQWxi+TqGLGWrYnLhuZvWH2opNQqa4b6b
SdYubmTmDdUm4xQdoifzn13wRRFK2LfaIn5D3lsC2U1VCQG7PDElt+rBCikD
2VpySvWyEgcpqYBBdcYMxd9QdyeXg38vnZmCRUOORrl97/jPtVRa/fUmZ9ZH
GIwD55ABh2gIcrxVfk33XAXbFps5vH2A4YnpUN+vs7Mu3xMfkzk+h/qodgU2
92ZN/LOR6ZfofbU6U1yIbaE3AZR0ZhQHZ98tZLaiPD70M54FvHqJ2n7hrQ3q
BmDE6TDa6YlkjGOsFDJcluS2ZB51j7blv1y8c81r+ZmwUiLj0zLizyCeotqT
CDIJ8mE7Skq11YXiD7rK13aovZBKJ6wdwa9lTAI5yIqW4aQiL8Re1RUvyd3Q
5h+FJy0UXlcbHnVoRE2maLbjvRx7k/vMLpK1EZWmnUCLrfni9y1/IYa51eTQ
TbyeXTl/DDmuOaAA8jg0oRcarDOozfybGfhwLDQbtPDIaX4196Ut0xaxtbdP
pRrz4/IXK5sIfx8YHLQ0jmwQW9zbovHFptes+QmQaywceXzP59MMQOSLu/Ih
puePPlowpsQY7lWoZEleOEH2oQMPdOXJyEZ2Tb0p7IVw/kD5AyQCYTd+E92P
zQ+fSdbKrTaC8znW9ByK3Ke9CJySVANYXfHuI+PxRRyLFjOjSFoId5QCWrj4
NBs2PF/8ND4sZ6MBFfOevcuLWtbXWvKKfmkdichta1NUo9Yl4owOtSrnaLU5
voRGzn6/nPROgZtFNyOJpdTDvP3o3nYlpAKfswW/WsjU7/JGz7lQTQOqXKNF
oDY84RHmlSv5AJDL8pXLku2f0yLefOwMeV+iWphMJmqeuyfetHmELsBmcwVP
j4L/FmiYMhnkimPn64uIOTISYjmT7nk9duf5Bv6kfu9WYydRoq3Xb06uw6gL
YomyTgwIjytH6FlJF8xou+O5IYN+s+gcje25uUn0a7b4lXq3cPGpIg+wk94b
CsPPnbOE6MJVSD38boRXGbHa0jXnT5I2X/SsRLv6LQBgN3mFBLPsis+j7SI3
fj3js4/lS+CH9VZrfO8hkE8drqIXi57yKhXYY/5PrtqqBrhkDUKaiMPYoI7u
l1tWFpf4J/Jalnl8oL/7vToKjXt+tuWBR8JBBCDY62aXVr2/0Qo6ilenWF6k
cYm2qDZSs9T1OF8Vc9OsF48wO0ujk9KVOupue6qebW/giD1QUDRnD6YKVYrM
lKHRzci0Ee2tWg61jLxCYfdLcr6/uXlwzbrgEux3K5DwRjW7i0M35n+NHmDT
LxD+TsC0+XhVLUeTiOjn4XEr3+VYzBtfOPVHqLGCsd2veOX/MeT31X0qTKwC
Ap63pprr2Z2576sl0gOHdDSJW3iOyYI70XEPB6KW6hCdutyAD62DufCS7m6U
IlhIvWhTAbU4NoRKAEzaGXPWEcvFq5L9u/Z2yZbJ+XTRJWFRLIkM96bzZ1ob
XtEE3ikqSMOaUmOtyjh6JFvQnsazfT2UgkSv9OIYDYjOQxHdurBhlgJR+vF7
TD3tVb+ZHKHtnVem6ubbeyPuTKl2zBtv+Yb4zeB6+ZOyDW41FWnRKkQb1+V3
TrYIINFWkRNXcTgWD6EUkk/GicYJ/EpElJCp2i6FFwpsWXldhK3bksWDT3IS
iOt9lCWh9A/FPWcR8GxSXuK25CJhfiMuqbFUuvkDMDXGZqYno20FiT76ZXNW
3isQ5RjkB1lkvzyNQedMYiINjUvHHkurEp25P2tOPnVDSnzoNkKV8TJuO9ec
1JtuevlV8vgupcfwWcfputKvvvotJiHgIMKIWpVsJsuHfP7Ry/eFx5F3f9nF
C9mtgQasLw9namwWo/OND3+S9Ds06/Xaw/GoB0+3jZ7YA5lMRA/9VYo2/Uz2
idPJ7/Jdmrt7Iw2JQaA2K/vqABQf3nHlNUtlIy8MjDEwzpg2Fi6+jqPExUlC
H8z81TMgBlthIUlxf2ykcglBRmmN9ECq5aiWRS+gPR6a0Zk+rQ4cxfHt6fvV
cqqWWbhl6mC1JNOC3gLbWoKsCQejTixvFjst4NzxD06WgkFmhIOIvd45KBBo
DPDME+q9yXJpLuPgQ9H/k22nqcF4AE+L3Hb57HCo49Z26TdXfzHKjTjudRvI
sknm2+M58Xn9MXejyPB+dlkouq69L1CpOY4BYf6nl9BrwyJfJrBGv1XCAkz4
DF682GAxmyHWhu7sz1CIeQRyFpcwyArhADwTbHx8F5X0jWt/eEwAv6LoC9l0
ZP8nnOo2/nQ9yirR632GaoeTdYRmFDlNMuQ86/mWxvljJIBcSz5ZS78xLE7B
HppPU6IP2BWH3a8HOJBB2CsJ6z59XGiXzmS9VsPNmbg1L/KMAHZv10s9akFP
xPIBwGUMjPjYUaMsEg1hS4vOvw9UV0nju4QF3V8NNTlp0kMnH652C1KvV7ww
u+3BzKfyNAatu2degvxp82kos6WfBPiZluB6Ghh6+sE2RyrVoN/mQVyisPaO
mXfsOS+43ba/78DMfluY9CjWmX3Uxkd/gJPlGDzbsOpxL7Ofoe1bUJ4UvsB/
zpA4FUP5SXQholcoEdg0jZLStCeIMDGG7t45m8UhIWrMkSKcmu/f0rfj1Nyn
EIV6Vg29iecwzztjmmKpl56ObetaTRu+CfwidUU188j+tcYPqY5ey+rsANPu
Ys+7cMC1Y0vQXdY1N/GEew2l0glzStG9gDTdEWV0mmOHflmviYomJMHEYWXW
ZT6DpwZHsq2PYd8jIse+0N3Eo+PHMWcgrYxj/jUmm73UDJrNTlOarYpoEen9
o6IQ1OSx8nrFsRoixtkpUkZzFvvaBcd9qaPyR2Kjro6T1pBNFVHjbaxQFxp7
8+7jjy6a0zRNmMEFYp0nDgaIDILivTmkbRN64U+CUHRpoDPGtMVScoKWaXi1
CE8cAxctT4+l+TGV6QrgrqQon0x9XqoX33Oofi6PtBaHVbYmDXiMrkj3TqA2
102qllJxptmRretffwFIbq1RmD0gOnHYsgHC4DCfF5H0A19cQtk6icLQiv/H
+/EieE+3XoD03vXcWlfVfKS280zaqaAhLY7L0Il2XEMUO5ix/y/U9WPRXAf9
tahd6ZI2FE9tIvYiKKN5DXlu3tqAcTVniXfhYSay1IhDl45EwrQoUd4X0XI5
OzAzC0ECiSmdtUmkBqk/znUcAjueV0xaKtkG3l1LBjFq5HZZLt092U62mSQJ
gCagMr5nV3e/EBau2t7PkgTT40WD4O+nddEj+yc8ZQL5U1KRYPFWFpIKEiVE
13H8bwKrgUyl179zpmlanIWQa7s+go9xqrb2xjvTa+N0HZZj2qFQ36GrZ0sn
4qktsIPzDeYx53rxCzdmS4YyxWRbayxidyY+8G0AO4y5pK9Z9vCeufRQ5h2e
zbVHacWe31XrKSQksJ/EOX3y7KFcxg0GxY1mRURcqfWFsMXxCdA/bXmjrtdB
GhYbTG3GLUWlk3caFay74rsnvSuoPabHuEv2rmf/Luwhop4OeQFpc++FMhU6
5u0cQWNP722UxqwBMzUjlSQrJPvPEwlFvSJ/fSFBUgvDc96JlyvZ0P6WdvGa
b5SYolFz+ci1m1YWI5Tj5iUuZLrlL9w98fHB1wbe23ClEhL5prFtpqFgv2G+
v+RbsvnnDY3vstmvDjQxngLEL7/egNmTrlRXWznp5OT5keGBJlDhsA3D0fJN
AtFRxi6KP/TOnJd0fek5w6xONn57F6dgVkQnpQgcqfwbYPWCB4hYtEHpWeWQ
dIsojltIZ7e9PlEhJvDJRNsY9GgtjKK1foq5f12Yx5P7RtYNzIJ5iqxvKYp5
CifEtPRSzmJul+VSFChX0b8uGgrfEdKXjJg+NxBaAZtbnUSi5rUQgvjtWmEZ
loXrUAb/ZceRm8+DFkiYD3I8U1xBFP1JHz1F8TVx/QuNMBJuCv6xIRenDDp5
KyvByiLxNxZT0kgsihczAP4qNFkVsNe6UCatsYwuqytx7Gyg/AO4Stl+gbhD
tFU87nVOafldmRLcvDxbP/8gBGKWrGs4HF3yWOuKU0kJrpzgZPbPbxK5fTpS
++a4Y9R0SwXBn/qdf/rrWxrxml/7PS8S6InMOQx8i3eXNmezKv9KpI3o9z7z
H0XjjEHEBK9JpIiZH7HvxKR4oCbA62wFqWY0GLWbu1lF+m80HgwXyPBJZsgm
vYaVqMXH7oGumv1tdcY3CyFPfIW23awuoM25HUw/hLJrRvk+IhBIW+7E9BMT
6D32Gp3RlqhONEgc5nRjJRDzgXLH3E8wWBytU6q3V0NefJFnH9GQyBGjX36S
4wPoGupVH/nHUtWkqGF3kal8M0+NmFBuGmPX9dXbMiUuGwcDtoNgbXd39xgy
vhcEbmtJzt1eC02YXOVtZIPTOA9HHFVK8Ucdh6bfjba/7Tz8VvqzChzdkFKM
jxdKKaPjaEevFXMzw5XQaWEq1fKNDCJrlKp0vuU7Sfu2eiGpT6peTt0dX/Jf
YebCHqnZBZ82OCzSKHxKg2jcv+fXXYRForZWDQ66OhnUQ2WHnCekFOuQ45q9
A2QHLMno4U2sLNyvZPmUsnHIjZqppwdZlV77CB7GPLBCGo9sVJh8raAmuuVC
lrA+UPA1jbm8IQbX2WaqkZNX9u5lnQQC97SPlD1m4ii8CYlGnKWBMDDj/KK9
7NAYxn7Z2bETQbrS/fLM8BKrXWarKuWjL9DGCnxYSWmsyLNs0lZhwhnIvud5
MDWauI71uGhlFpAglwW9vPU61VZlpOD8tpXI1IrvsaXj/421AeegYg2Q0mZc
zqcvI1LbbQAN/TNLyNo4tdwhwsLwDXwzHw9uOMWACKQ5dONoqBWwHphZuj22
O9ywB7XzSOxbp95uGDtuj1D9n/sjMbZpkZNVZgAdkhJXeJdJZ+80vBNMnCNG
jYH1vH4hwWMOvYfFBixNNdem73RtYwxpFaMymnWQNBKcYpHZdXLOsVkhuzgR
PU9372wxl3xp43yF/tdd2ULmbpvVLhRDBSI2K1/r+AFVv5+jl/dqJ+RxmPrt
bdqF4eLsOdL7/B5Qgq5PYc8KEtd2V9isJgsnn2UfbAs+OTc5cdbg750d+f8e
0tSjEPNmmFvho/ayl7BTE2lIMaFGCiYKt4ENPMnhbjxVtxl1fZ3P4OH0Zyl+
hKrlFqS1NvXr+8ILWAfNnUwqv0QX3Ypzp3Gmfp5zbEJlbpGdLLzmN8sYC7qW
FPhQbuxuyLqxbfkuHQ6TzD1WYS30/EgZRGVxRcV2JxnA99aMTx17XQlv5n1z
1q5SqLoDDZLW4+lWrMwJtI0UAkZ3j1ToEJ06EpLzBPdO67u/YXT80nk3+R9d
4WN08Yhqx9JjN8k0NA58TTRYF2FA6iFixWNexpNt3VYeh6P+MoclCl06HXnn
YVnNdA1/es+Y2eba/2R5gcFM9U57gybfn0vhiYPF2UB4JBhQDrcBoHBZH9DS
WO4hvJIo1w/HgcvI7OHi8v30Svx5Nmz/lqG/OS/3f/4jLUmwEg17BVKjDN0k
avbUmdQiVw/d9de0rlgARY6lD92h7lwxVNO8Jm6Fk6QFHtTwoB3RyEQgbL/6
RHffKnWsZCg3XTeY3E49yDxG5v6xC0pREm8wml/Azs1HiX6ZL4YGAZ6HIRr2
iHH6jpXejnvuSk3jsxLAb/LU4L7Bs8Mydcd5WTRhZJ0YZ75ENguXybhP4bG6
+Mpt0YXiJhDpZvd0fYIenBvqGkwK2brFZcKHD8N5PNS8zg6XWhNmKLrgW5cv
+aYiMN109y0y5+Mjv8Gsquu1lh+W/EX+bxwjLtCztdRlIFkqlj4VHgIxH2cQ
SsQTOj4GarqHq7ny4iOarZTALazfJoop/3tW+mJmwratUJYgnt6UlglAbcvw
uj4XinJWMBnLT6OGxsqkT8vaha4jBpOCI7Fw07BpIq3EczV860xCN2HBvyNz
+rMJTslBMdkOHoqFrP44dUNdfatYGy/UV3114d7ZE31UeB1wRSBxBeS2wIis
yT1XBQyCFHzUa1qpMCswnEtwJ1uY6B/pijyz+A43+HDV3RC1rBV7fjb93UeW
LfEDcrwKmHsdJDlh6fzURyaSiASwDDz40NbXBvspNrspUesB4PiNOOfweYby
Jj4AI3epMSXuoBwWjbEX821vswgENzWayR3JlfFN8bOkGg1QwPvPlyglprPe
eKZWZuZxmv7ID3LcQ4WXK0K0YptZ1+3aT136GyABXoEuwYRNVDMMMzdyJWtF
4biTBEZZGph5N94agvhBWC9VrciQKhPueY4Ye/Wkrwhbh9rEoLRLEyGP19zk
flmRhSiW7YYQLKckLgESgMpLl9qdq8MCr05GotcAqSQcu8jQ4T4PJi/htLQc
oCioyFBeNb1h3Y6XHQn1BTk5EyvAz3f1hhtPLfA2WTs413leruZAVJNqCZOC
m/XsOOMO1FdaXSsbbcrMslhp9jJhzWvLyBk8zsc3cQkeeVseLcRWPuChiPZ3
GfP8F/q90v/wagUGyAg/8zi5BdI73rnxOLCZ8G62zRHkT0fY2KYy0mLsP7N7
6n7YLUGtGscCjVcdDwWXSkqkfaWS9Ox3+XkJdjwVh0tgBhdzlltPLdBNWFfF
2O1DV6Ui6jOjo+K9fT/lvhsco2gbMFkE2Lp9nnBCLSEbk66MglVlp9XkQ+r3
G4DYII/iRUrZVdnTThiSWaLBNYkxou4dCOQYUnWVKlyJ3EdTt1nBAPfUDjOc
E6xnsqq/1c7qUZRi7xOXgf1OfB+T1+CyQ+aZulVy6wuG+4xA8aO/S3I0Kzqw
/FgK0dRG1QHU5OvyqHX7whnqk0fm+JHPYCQ6enhYvZV/jfDSgqsUr2xsg55z
npBCwlWJ/PoHY77NxN4zrLQeKNshq8i1Kg/Dq6SVaIEFbc3hjCIbjiZvLZeV
E/NJx5Sl/A5AkYyDNCAw/4YS3xbMr6zFwd45TlMp0gqun4xHeOZE+SIhhCl0
DmbT3QUgb3ogmJoY1G8tpytZcJiSusTKtScbdLSWuug536DVe8ZmpNJWyVbJ
U8lb43XAfKr7rrSSTO5aM2DEuMAqM4E8+CdBm3vCCBLmKlXjYqaLH2RMJHLE
OI3o1KqGZ9qys5cUi0bhMsvvbvMRV4T5ogbaVaeVjfH+7BbB9HvkWxFfoU5u
OFSYGbcGpOM9SL5Srcn/kNRFf1iMlIVRdAe1bgGL1sh1J1teWTqnrjuKlYop
lSc0++KiCh0l10rA0mC/cqWoBMmXF9Hq4hekGptG/2GGls/e/0brbdvz98BS
H71cMstyzys3/GtuWziGvOI9b0c+YlfO7vxC9fnLgn1GqN7iLmWBWCI8mVav
D8p2cc/RloBAbFAAhx3tvC3EqvSKaT8QToeSI8Pcm58tmX4y9/ZXPMxMFGPm
ebUnOamE1OqGOUZML1/FHd7gjcH/ZYOzwe8iEXkI7baSDmO5ZFq8b1Cabp0T
jq6dAV4DWFTsc7FS1/TROzELeCnYzMSFuTzGR5rDF6TgXAfvGPfuwA5i+Yoh
Er+UJXmNpx7o8lafzHMsg07a9oEPSGibaLZvIzype3Zdqll1Vnmg6mKEqD5B
ZfGspaz1KVQIyIM3L+QNSKeZjmdNmcrzaPz2319UzlY3ggO0lJSY/mrdPsVB
4ek1sYu7upCykXfVaoEQqQ9NPZEOPeGbBOB+CNKTs+yBNfNEa95RAEaV+tTD
QDxC/5KwnL4ZG9Nor3fCkc69Tk4NStnCQkNvsNyflXImwDpw3lCPYK/+OYFy
H8y/EUtAOCYooZXUPq82p9dYWwe1P5Q+gkIuKZsqjNKMSCb5T15Tk6hR2t6Y
og3pxQfGNjuHxDbQ4LvKOi4ASUlL3Kz4vj+5k+auUovhLXrEAH2/zbzp8LDt
RFAhnfx3ZuRr+qErKNZoJeMWdZInhMFBQQKy1tCDhglHiwdItkcRHVEvL+pq
qFWBRzdxcNAlvP2UHPt4+2iUKLV8traA7BuLLCl1uZP9Yy1MnJdav3OR/YLL
LbMyRGvqtZ1/eMirM6y2CxGEY13daDQ2epzLUYQWvzjikML8HQODzB0gH/Lt
1jSjcsV6IdoYSAR0JDFQap/J04hTHyMPz3UCnzKKQeou2aVJnTeYrRWSaL6m
/Yq+341hgFtiuG6Ced8d5XlOpxacr85e3c7byR+Z3c5lS7XFQR5DbUAOMrSG
cQFVqo5sXam780BKsxCfJbGnY0qmzoO/5X6ImTIkzq++H5ChTjk4Iu84uVaC
B5J+kSVqsh4i6gvFYi+FCJIqpBGGCTj6aj7cToVkorCzL1zLHKuvo1W5ZW3M
Vhc+1kVODS9PVGsiPvUMKCCnPjU9dG6DGZ69DtA3yJDGGhJY/Vh/55NCu8DM
H8IGM3iOPUPBIwehlVGX5ZS5+EuYCmKpw3+jjmPFxCBq4qqx2lKqzl/zkzbP
gHfy3TFaiQGvHm9zSZsB3CJYHOZcoGfWg16tzjbIoA4V5SC14nckYaaOatBQ
5N8OJHjOBLgVU6uDnFQ3qiKa6L2DVBbxYewnWfimfulPBTaFWuCQgFg3HfDp
f5w7ZrMktD/uUaba1bpzQ/s8dngGGUldpOKOZ4A0QBR+1XDoOTGAcx2qYuYS
iKXsMBGFBghVYAXt9HPtxkccKxhE3bd6TvXt1eFWjN0k8X95VHanhY3jcDU+
Se6PFuLDh1BF/TfHcOHRPlGlJHJuqx31eNyyVj/MAfh8dSutpICLSWL60Ja4
ox/vJUjRdrPLtmyLHCLw8A4mc3xkyicKv3RE9Xbwcz8t4be5CzG/jQdIP376
6wq6LYZB3Hv+EjLdIWXlsz90qbr5M949o09hbZZQDGq9O+63w6e3bpouvzmf
WrAVy1v4QzfoEED6hoHm08WM9WaVIa17z/YTfJDW05V3Mu4k3UTVhESVcyJz
xVGBF7c/9Ff/X06ngwufmRpj5azFJRhtVw04dzcazHxHQDBJxaPWvc6yTeC3
nWCP9JSEA7rbkxOq2t7UW/Nmmg6StcGXla+iVy3wsY8sHLQH2y0bT410bDY0
zz5aHPO8qH6DJ9pcRSURriqaOxqjLN9aJhZ1QVHbWSrE+08ymOo0FkvVNYW9
PhtwX57Z1W1Jl/aSA1AmuyAzu5q/ArVvDZVeT0eujhWU9N//6IwCOXkcZC+G
nIFIpPccq4k+C9caogt4kayKB/dqTh8iNyqhfaaKCVdnVKd54FdkeBiUKm7Y
o67mDMEDnhBDizDj0Dr3s+2JTyHVvD88iFr4FcH6zSPd4JQVQb8wVqUbiQPg
ZbRpkgdr4S5WlOWoQaZUjnktKCG9Rf+HfvOWU4xm/N8v8cpKpTGWNPbynrU0
vrEiV0/bU31I9OHQfs6S7qgf+lcWV13ExSm9/XeYyMpG77U6DXaIzURtQpaH
EYE2jE1kEeDdhrVws95JZD40LYOufEbClBmKYtm7xXMEjLSQzXt6ihgQ2El4
Z9CCqdlkIFLF326ojfrq9Y4YY1hqiS9+TGfAjnNWn0RlmaqXrLX0SCMLXCQX
3r8fmGDtUCyfmrAgiANRF2R/52jrjTS0PiQAxA7YjN21eUXgowHGQNp+966h
1gXqujaRJ0A0urNL8Ho8YDTF9wY8lHOWGJIU2R/wWxUnxz4odovPzBfhfV6C
CX02lOt67BCMcfu8dPoc0ZA3yvnOUBVGm6sgJxP4NjtiM1SUfDmV0YRDVadJ
MUL2t8jFcWjrSDf3M770U2qzOxLf4d/Yf4Uxcnfh27Yzcf65rVFok8n19eO3
yH9EzNEYfw5uNgIypK7F51yYNS/MotguY04Efc8KIPTq9kCNAOqw9l9oU28d
LAm5Mwm7vthRW6Y0MXB32Ui7an/ka6dGgfu5t0WsglJ1qhclIFABV537GBr7
SEd5dNH+dvqpYxrqBO9PfJUp8/SFCOPLJBOKS9MF09EnSUyS388V3wPa16E0
rzkdNLNFZ/NlFe/0jmF6CkRd/0isYl+yzQ3bBXsw9cq+VW1vy7qkLHSSttXO
yJrc+dFT15vkYNBkghuWvQ4+tLQcd7w/UYX99EWeMM59DSOEj9l+KgKW+Gts
eE1zKmcAeEVgZKRs8l/+LzI7tgcPo1n7NatqTbzbDsP0e4Ua0OkHGgd+MDmz
5rUPl9pt8SXRi4mXomPxaY472yfxzYFLYeQ6BpOUroH82c0+rvPLOMrc6Hid
UZCkQqCUtEZQ++ZSh15NjhrYo20/YK55JTHHhdTpwCmnm5Pyye4Hq65H3BD5
m1jz5AnXVYPdtzGRjNNeW7IjYglIZIh5KOUJcHUEm7j16hilO5/gSnDn6QLB
DRgJ0dZe5wXJRLzFYnS0Rg/jAZSO/gkzNgIOLoUSJiFx7Fr4ZsEhRMNLzxK2
G9dZw1BxNF/TBl4EJZZj/gD0DjenpuRYhFfOdcaNqTTro0+/3Gbd3pg5BPnr
+rKf84Id08nvEK9AxpXyoSnHtmA74Piwo/7I3RORCpQnvnUGlsmFO1knn1C6
5xLKLgTP6WS84C1mKnw+aUzEwIV1TYDVSh8YKD9WcS0ktnC7/tWnMKhysN+k
EJVoM0oMZdeHLW5bUWRowT2NhIElri+3307PvSUHvS5rpg3Rj6x6C5hUbfAS
CCL3gSXhvqeN65vyB7CYeCv5Iu1/Lgvl031ur2yHXX4zMvxawqeFem7PF69b
vOSRoTaNwzimqFbwU1rfA+lFmIV5BwhhdTT/SC5Txr43V2tR2qQ3W7iv0Ajp
Aq7xy3cXzNdlHdGPxOjdqgj7jjbRlOn7v5do4RHPIHQ4U9u+w8YxXBUUnqfk
MAohpM6GpRCy2FxPb/Txkelr+n5iepf//DmcDHP3aLnFeMHmuDKxgvXcCHTf
KQoPFmqaZG50sgr9uu4309izcq17G8Q6Ye/UOxsu7qV6M5w+VcSgAlYkfVf3
REIu9xIyeL8mXpt6sKv5c+BC6GUJhrL4+D4BMNIKTrkEMKWmHFNAaH7jA4dh
yOhHGRXYVNpOlrOaFBCrqD+fMZlPNAf68Jo9G+6gmT2RLF2SnnuaTOFfpnYK
E6OqNC7IDXbzt7ks/AOCSNCapsGBYpCSDR6h5+j/6A7ZkpUbzCkQNCLSZotz
cm9Gluh29KMFunuFrplnEuYN3atXE1N7BOVvrmbcLvkCZuKp9TsfSv/jvh9r
20MudWcWTADNm8xdM54WLYNo2OEEyrLwWFuz2Zmapv/7TzPXwlPHqrFdnp03
NfRWxI5FvDBV7yeG0E8WfO4x18r6TVML95Y0GDN/s8EfLIW7LGuFUQMfLbqo
mrirbd4TrrnCsBEAR6qCZGO+O2VL8OzLiX3Rigdtf25PwKxZaWTIa/RwVnM5
eqoWVzzvBm1oBlqhdp2myIskfpZPWGz6kGFI5Igt6a57PmwC2tUxeqwPfURx
dWiwxnFbk0Qvc4OFpTQhy3abhkcqpgmMFKFIyhA+woOY8Z3fVsQvT2Ri7xuO
hzyowuAQGG+E7+QDP62t7y8btHqBKfzzhfLsPJBqgRhOhuB1fmu4QAReTIop
i00d+bVbY2ZIy4hRA286JttwtuHFLph50qUxK86Xn4e2i7k/uRqgYF20QnPE
5yCe2GriCJBltOSFm7TAwCgoSVluTQNcrGfTPNluO/VsoFtkYA9g8ZP/+4rf
B65PE2YULXHLrH3nH+ooISZiTZyCLnx6301oy7qsjWLp+x33kZKoE5YuGI87
KNh6BP2cFvo7GsOOjMf37ia6l8X8Uztol8RXREeq7p8fktx2bpzEz9b00kZD
+PNiX+UyqYj090o5vh+Z5f9+np40rdrsyNvND50+pDqMQ1jDPaL3bp/6pDNH
hw9LRdWi9pnXuzsAQw6u8fja+jCRb/zonSGecEWL4oOwdGm2aKx8fuOlbp64
CRTDlssVUYHmtUwIKCZCS+9Udadz63fAzM/2cpP4Fh+h2EzJa7XPmzN22Put
xmXjsHDc2VEwiag2YCRWO939zPjEiKnlHXgYmvpWBHtj7XHpmSPRY6VvvqlE
Y3yGXhAA6qJChiHrTc3jgbMaG8Glvet+2zwEjKbcqdOb9D4e2P4ng1u461GS
JczuCq16GqP8NWht7gCOYXYlRbIbw1wbNdEs6uViGntveEw1tbXEtDWCPRc8
7h5tTLTuXF0W2ZB1yY6agWjT7oFSqYz/KNVE495brpk25bFAGHrmQAnXKJFY
QqU3xHGtHo1XVcolo7B8/20UTVloQTOPDiPwhFLuSXkwUcqvfVH5qy9K45E1
xMgL/u3Ia2vkbTWj8oR/e3OVN5mqez6RY5E2JlmNCMoVczVNGRNFD3q4Jit7
8D/UfXk/Ku3T/oO2LkrD4vYpNbzorIyPss2jcSVa5cKg/H5sZYk1v9O5LLRl
HxMOG5Ts5fGVNc2mgxfmw2UkoHDPg+UXbEnN0RE0Igq29vv6Zwa9cOmAnh/H
XLYTww+OUU5v1zucpiO861oQevAMHDQwHs0wsMLvDx27/0G13gZpM3x3uWVM
RmBpmRNPhBMM0Ru45uNZMtP/sq9zFaZsGmneRKyl5eFAUXxH638Sz32E1EzY
wH6Gp1CdDMbym9UbLq6pe62ALU5y8yVxqMLHX+08UirSg1r1PaYFacUJhgxR
Y0EInEFeKQgD6FPRtfrEP32aQmgiQGp3p86+iJYiiqc36iqTzjFIR9Ao2SFT
YM5PZO60hyebjeWVlPllxKLX0DMfwimU7D+yCzVFxir8BZRKLvH0p//tC6ME
fELHFPmm4bLU1qaYepB5VA6KKosG3NRzlqgcoripvt5Vvh8G22xaqUys+tc9
xYm+l/2xlQeQ7ruA3b+XiYofPAdwmoeEdozGQA3UJd/dTKuv4IPkfGUl0ux9
8NtmA2m0KC+ekLSuu7alqoYvoYZr15qt6pNVquKOb1E2GJpqBWrLHr0dXw31
6icIYmMOa/TArXF7CxsQLXIWInh+d5EmlOWVcjSrLFpgWyQ+x4D6KSKqXMGV
cBizrYJhvy8Mc+fjCBU5HQEqTP7EFbYGIQSzduALFG6odDQgC4R5XrkhIdAw
Ns7IJPxR/HMRQktcVNHscBEvhHQBPZDFYxpKhICxaTi5IHbRLRJVivc3H5mM
kfEwS0QEIzrap5QqPupyQb5vmBjdkcReMWBDP0gW94wrwA0UA5j0KWOelKok
ZZpjvk763rYfhy7mf10FiNjk/fAFEIZbtO8acxRkR2hbKbe4vrwSkvrtxjBD
6RF2BemozfeLxXWSYeRCMO3gqO1wq/nkxqtk8OnCfFwO/EaTtT/vQ2Yvhki5
LckVH3cYBxNPTp98MVlod2aAk+KfGRERI/ZOb28JHbLxZmXKqD3YrydFSL6/
pTeJT8mX8l/J4/9nr0D2e9PtCvQioyFUum2JrRrE1obOU/wI+BaoQ4yuafEK
rLozpeEGH5/4YMdEVxKRoOKc+HpP9qMoXFKS0kBEJrRe8YCfkgsymzedhx1a
zDkEM9q4U+tIBEPubK9XSuf/MLeBWAqPadCUBNrb//uftRxoyoWeUqZkSnzI
nJVAIgBvUz77m3MB6aKEtLUhwkxmdY8HKCDP9vpvwATWy08sas65nBkCSFVv
BDfLo94dvDYCW6oD4aYu4bqd0/YTTw/1PTR/uBqoIYVcks8QvNMTz6mbObM0
0MEBqUKfUHT17v4QuT6HmtkZz2+5Wn4iPbgh1Ozfr3k5PKElUrLnZ2k3sCEa
8vS+DYf/7HDEgIc2Usba6f0KY2dJySHqrguvEp2D6j8hzO0j/h1li6tC6XhN
7xwb1whsE2G3OT+Fze/XvYdDVB27dU/Ie3K7JVyW99BxP4tH7niT/h4seTW0
/mkVWkp+aJXWX51m1kjTXPicYdZ3c/lrE6BdgtQ45u4TYHdBWCJyilXvXzc+
KiEhBCFNDOVaBkueG7M0GtyC0EMRyt6+x8GDJjWynDoo6Xja4imLOKF2ktA4
FXQ4+QLnqdINJHZr2F+9Fpw42Xhf8G9zSb7UHZpTr/wykfhx/V9ddpA0ocpb
IpmONyYcm/yn0dXhlBQ10CFC7xxUi3Rvg5OOSr/mU/lpr9gG88JbV0dNVF2v
Fbdwy8LCtgPYIgQWuWw6EaE+Hi7ee73MUEOGnVTLTpwyzWxG0GPr/ik+IQ+9
Wq+Ukl+ef2491yoCFC5NVfud6mne2kKzjf25DKA9S0M12keAgKH1rtKctnaB
3nW56yRLjfVKZR8xOs3Z0aB3D+JzS9Z0dT049vk3wfBlz+4vdd1ENoIaVfZc
9PGKtcoBZ/FhxWXGIcyKJDhTQLW/Vt8tjPHzHWRnMc363ERIzM036sf22c1x
H6tO2wppiosgBNz2RGvFf53nSiXhZp3JTg6mw9D5eZoWuMg7asos8IpzvuKN
YT6oZ2rA1pY8uloj1py3Zg9GdqY6wdoyh0uvmLZyIymUF+1e/ajDihPx49K+
0OKdXZK4QSuBV5LFcLL5PYJWv5QtHsgRCgeS+RLmES1BNgYDhz4josgT7BIU
/84t+Kz7RHp+1cgAiuY0p+3wWBRIa+/FYJ3E+rmVaOd+6dpCl3ZzHAg3Lx/B
N+pUB2Fs85IzTLo8j4lJRejMowEE0N0hJtCOblgFKcIVSK6Enqon5KuaE9bS
FRIu8GZGD4HWebjaNkArM/N1bgDOjMUsaHhyt4FeU3Txnz0pw0ZCDl9OOb9i
EXByZ1Gw3orLFurO8Xkm892qNQUkwtfTdewKHl4FgQrUOVpmkGafPfCcXGcq
oQwJ9wPY1SfuF4+97qafZDGbTzAh/YG7oIsCdegZZ5YMJa+GJh+frZKvUhnp
wtZfVyFExg08FsoLcJ/P3Bdee9dpd/whrjydikPHg/3Tl39dh2XiB74afdrr
YPBZjArUEkb5RYZpABEwFXWtClreDXmR31q2T7GHni6Hzk/YU/kMFX3HXFuB
nNw9dJjvYtnhIpRaM3v9mzAp2DkPiYpEAxF9D/H3XfiyAj63YgHj5dFw09p1
EmHE+EKlqT1ay2Pb8rzqPb2AiYmpbU4YRQyP1WlrS0MrffBHGlSOCwDuCngC
GR7eiyf1FCRWvr0CjH8SFy35eRUwkWilIpzwolHeo2rVfRhzQNyO8L6oByiO
VomAmYJStkaylnjus1T0+pyENaodYyFZPd1nmHgh4O8j2f8AfKQDXcOwTsvV
jkL1fCseHsDPlHyJPf946ALWjpiXSxAMdOPQSvP8gk8toMs56bH7EIrMZRxb
X0ovnaNiMMVWYNNOeOBcsQPW8dj2+G+hHL0r1h2Tz6Ag/MYIDf/fPFf2iXLm
5y8jEJrnhv3Lq8lG3/Cd24mG4ocy44NJstbSVLKRXtu/tFwpcb/LI5zNA+B9
HLQx7L1kJSpPa4PQNS5sZtVN5/JbWgHGcoh8E9iQ54FxeoHy+dwjBo5EPvfY
w11h+t0YgAzhs7ZELRS//TduUGlwv5892kTxegPzxWEcP2Al04I2XAdtUk+L
9Dh7h8Ii61PfmdGQWhu2Ep68y/o5ArzhFRXl/+B7xxbfpIWKuySPcJyTgR0h
xInZg74GGrzTDG1BfSIZ7xUKcM6EESWnlEtF05QSzwU7k93KkTQ+/rEn14Ba
aWkNmPzFcsk4pEQplIl9/1GiAF4DQIXdwyuCvJEdVtfWbsBarGZ9Nf1/Mry+
caOglsMKU7QyeZzPXke8dKe3zX3dAMgkABJVD9KL39TBU7k+CxtPfYSCLfP+
vCZMa8Ld0L0oKl8IOISFEKsfn8TYHYGwq0muixITtlH/cgrh7Kqd10IRk1lc
sHUmnzWkmbBJ0CjRtuhy8sN8hJBgLkM/2Mu0fnLYhg2vNTyvONszr7ywn67c
zH+mOF9d2/M+QFTQNjR2sZS+Xs20e91sOab0t59YgzPU4Sf8nDk9YKgKYNa5
KKKmIHvYqSyToWcMpeunZ+7SIT/tH5kBpWZHpbZw1Niz2rLRURJ4eCnOFdVt
5eHrCXHLe2uliVOG7Iq3Bo7qmSv+wNQIpEZ3r01E/KBxtQQLCSN3voB5L3XG
4rs/XTuAKr5A0Wgge1nLg3v0HAIAQ0bKKqKRLj6IzaCmSySuPH/o9U1+cKFd
Gr2YxjGJQwCnkpUBUpBdwPcW/RoUgCxd7yMqx1dTYBxpPH71T9SmyxgIAEhs
bdtHpg72ZqDB+zFWcEuUWz/ah1i4/yEY3nXCXautZNEE0WJ6278GdpjFS9ai
X0PZPt6r3ZJ0FSBSCH8GdA3S9567ZaaB15gklrJvadLir0H1mKJvniVcGdu4
RYT3CW3YvEIy0HodUd5rPXq5a1cK7U/4TlyZDCWl6+Z2BWRQAIz88fEbVcJO
KyfJmoznl43mnvHN0djnXZMchkz9mqr+Ku31MOtLta69sXn9eDi8G1A6+gwl
G6HXfmHwMce7kIbCBSKSXKve16IvT7WgBWCCKLYqd3QyVdCYhbge+WjdYRwY
DT5DTvy4t1UccYqYkSj9Pn8V+lBDd/IBJQCaOPrZLN6o0rMlFElW0SVDUFn3
l+8JghSgh7YV8/ggWxuJh/oWJIh93mX7IQobLfixTatKlglgT5vMhkVzr+nE
LzZxXVV2Vtu6lq8kfYPenCFNgWP46nFtzRIO+0zueMopdIWhaF9FhfUXCDfa
Ypr6btVA/O+f5RLqsffEK+5NV6Sg1WA+XvLRT3vgvkAnC2B6Giz+LUe6N3sH
Hcxyq5e/hnb2kXnAaiAxG5iOQqnKzjR95VjbAwGjzUZoCbi7A/tZ8QbDD95O
gahk58L6z8AgGRb0IMTwZAmDl05soRD2PFf17c/g0WH7TwuOyhSVfvvJOGsu
1ZrLUeA1vSZKpSeOklWT7oiiaEsxjYMw4jUcmUcvioBIp5Sp+v7Lp1Gdd2lo
AABqf2jfXtmbYHvhkXWeYD7FFQhohJJqIRd3FKzDqdFlHOINvfM9aT4XnGQ4
UoLczhj9bHMu3sYkLCaPjuhbGE95LyZz8DErPkUFMqPrl3lygXw/1/rDk3kM
p84BlDYiOhoZ0ltdtpIjDeB0GOMmozkmzFHZ1Cs7LKUEmxTY3pIWa37nh6/n
PjeLeu1EhpScuo/JPHl8lD+zsRs/D5ORe1H98j9Af8bU4AS+jyMdwGfu82GZ
ndhV1/tZ2w2si/g8+Nx6TZhIhcgKKUxPxirh4aH4IyC1GZ2AYiPhFCo/TVKn
thAn2pIdT6Mvm/nlVRaqjpx8MRgk34kGPjIFysyLgnh0MbmaKq2vfspu8Euv
nHfdJs9fzyCkb+USSDA7uR5K2Yyl3aHTaCXxLUrvGtugmTu+TAR3dyAPQPnk
WtNf2yiAadMuVN8k6kb24gVenScEh3M+74oRwI1Xr5RJQJBBQAVe3+EVfucj
sWmC5ErZSjw259innn1qfA7Ch9aU8NCKhzx5WSJFS9fCzK391rtOcBUwshzF
T71avwamJAgyKibwW0eY14G714vQmBsJyULcU7Jsbk07yuaUU9raObqCF2CZ
VkWibH4Iw+iwboL6zCrtVKb+7JK4xjjTFeGkoc5zToUkaeZyUsS+8KJLAGER
TZ/ZmykEwM9jM1qL5MlN3Sxo+uyuSkUbzUN+HsrHPJIRWBYqJrvMBEyTU0Mt
CvC9By0JiL4OS/HNfgOsXRs4nhdDNNhGWsQnF1PWnwLiPBT2asU0brcz7Qf1
VGx5BOy/9myPLcyv/6bmrb5CytKFlonHj5CsM5lUw3F4rPiQ/5CpR1ArUaet
AHGZWKblF787N62LyZdG+3fQqNAdRxL0wu+SLUD/G+oRjQrMF2tjbgdYN5nm
wUkNPLIAuPBVRGr964p0uWvn8GtcJ/KMqHy4HCPr64j6joxztXM3usR49OR/
2F/q7K9U34ZOqublUEZ+8ggpP2RkN8VdaOPKovH/de5lOhYZnnTIKjOB5thj
eUGO6zwPEvWKw2h0Vve0Ynk+uoOaJt+0TDzA1iwKNurSLoJ9oDuWsw/jOZBU
yOQJQ9jP3bJAUPmvBJcu+3790Kg0YU39affhMccoKhy3KcE9ZFpdPO7ay20b
3LOVSB088XZgLEkMu/NFlqBvjod+4dsQO82a1P5dNuqh05s7lyrB2NDdHOSg
SGpadQrRh9g/Wk95iGleCIsXRrm73XvTCILYKq/dwHUGNAoYUYC2Byx9MrX+
y9a40x+Q3wuUzVgBD+nYJOMlbNAKnY8PuwTMbGGl/xIu86xGKFEhMkwOi1J9
n56MXz4RSZdrzd/4TyUcdBz0UYbZru5dlLBx1OYYmXpAWfxenXkgy1estqhS
cxf06eDLdCIbXf8OgUJKXGykrQGXOmrr1jg/BUcR7BvAnjehNfq7LETvTuP+
nksLOOKnXFW+rp9gwZzwbMFo8CRTszuOmuSawnE9B48r1EzdvhcOskMcMmIO
i/BziP8jesau47v1ZccynUaXAjMgSnJERicRmTprv9RvgKzfI3uuKnXjl/MB
2GJVJ131QJF1UftQGW+oKsVY2Np6/yJ1YdlYXnPPBwS+vE9oXkoN7YGKajWA
TpWB8bJ3l/keAjW4qm73Vi+5RltN19+xcPaOE31YKaAIVXTq2EI9SL2Syrze
o8Et0PpNf/HYJT1ay5+qbEewG6/PKQhCiU23dmJeM67JnI2D50Cp3sFfwvnb
68dRdZ/WXzHao5rO1TFEfEhJLwt81CJwB+JAqt5BQRXc3U8R9lY54h3avc1g
NmHg5NhbtZB6/a5VSP72xftZlXtzLv4DqSy5ef0XEJDY/Lh1OyqrwUFNpJwZ
mSVjheX4Jetl6jubUe3igEZRNeM3xRX4DWtDeDzhjGtkYG0eR8+2+7wEHPcH
9EMK6Hqu2hMAzjVO20M5N0sTF855jC6Cw1D/S6lgQxYsu6ncmjeoIO3t4Vt7
UQ6YgsguLGtMrh3tjvhFkmU1UZvRgf5d4nYwHedS1gfoQ2USp8489Fm4Wh68
4GJWypOJeUmtAuvMfxsEqhgMbsxkf1fThQG4uCOKa4b0GC2u/lnWG2+PZ6Oz
6yham/xgBASlFBDWr5r1IzNB1jOqBOZ2gaLS10gllWM9pw5SA1wKoqwOD5dl
J/9Iof+eBFyEjmWgyTsCGK9F/FXHniqumDSx22k82nXzl3yKxBZGZBYOloZw
KOt3TXt/sIpYNo7XTA7h3nC7dU40aufH39MqBMkyDNgGRfFwWbV/zXdraMaF
QW1MwboOurei/rnnwCe7Idw6d0YtFcvaDLLejFIVAFwrbEChlKJjDFITclhc
7HAwFPLRAJmQbJfv74alNLaXNgdXn+bRcn5loQJivT4QNFrHfon+MIJexdod
JW6+XzFyxBQVaTq9VRZ13nuVk4m3XfVTbYiVt/MrViIinD3nbtGBOPB6dN8r
c2NH8Fn6rnZe7I3ok1yrr5tI2QUqefbq3TwHPUq4hoYe7lwF1//s12QCKqLv
QtnuoVX6iGA7SPTjcHJqKgyIzZn0r3ZLhTNHJXIDJbBhM+SYGNroPs5YOgq1
U4WiQYjhnSjUfo/ld5zC9a1oZBPqWjPrCvpijIHBlH9GDnlDz1LlK2h2GPFE
VlPMphfA/7ac38ISHxedaKbDfpokUUQ2u2MhXeJGvj7c7j+eSbqDmaSC+SUp
9FIaXQtZ/u+bb1Y7hOywdNmNMHVj/4WsunKoatUe0hbkNYbwG6zyc0dMYLye
yN9cYWCQN6HUbBGNQe53XFcxMzuBDELkJOtb0gvPfKEu3FywzebwOnViw53x
hHOdDJuQ1NC5fZtFZPwuYhOwicEuf+g/uiJrnCg3KZPSj9qzEDmDjY7QQqhl
zd16WTzbZ5bkh1PucWznzwi87wnSezrmt0IkOYKvlDXafIwkTUrmlE/40TA4
UdI7APB0AGS4wkeUquDM5QMC18E5GhmSCAL1tBzTwbuOEzC/pbsmTf9Mj48R
L7oWSvuAuWPC8XP7PH4fKVHfJSdq59PpmF0oev8ITqGtEk5GcOOs1R6/JRpE
h2Yfey/yyJeKju7hUHNR53JcjukxEDu70m8rwWZIhIjVQyPGDKAnCn/YL6Mm
SI739riNQnvhQeAF7/U/kzLbBHXAFdilVK5eYGAZksYJwZ9Ks21CxuEu9CL5
6ps4wUJqkZ6iaeRX/RK4jjnznU0IDQhjOOK3DL3uoli+sp7KwyKSaOw6Cl/K
GSM+pn6IVfAM5ceI1BeApD18qGVq0eSsqEHB+VZ17vTgt5DPH9Naa/BqOH+s
sm05IhCpsdLiVWynUHeTPCW9HI+8OXOQ/MRPC/ZWv3+Ny4WJmwK4rNlafgdb
/SMo0Bbkul7X8XpD1sdEhEqB92KRudMR9LoKgAGFiobWoqESLcfO8fiMah6G
W48v7BwwKZ0oXjWaw3cIci00f6N+ZEUV71xRZWUNESnbnn+7KvZodolwlKKQ
LbjBBYLdiOwBuoOkwrU33imYndTGV95cyMNPLNZvwEH24/vX4HLoYkcB3uI2
yEdZxGRJOZZeWZBnlz92pjoufLks8UjgARW80NzSl5YAdSpzjEDOCUnOtVLl
GeRbUaCTpylIfMxg2W7bZfI2fN9x9S/PcIKab1KTpD8ljhkMGI830Czpf6Px
kolRnaIAW+CIOrEoJBd18rLrwSDony1zlstyGF6o2lNDh6s65hz5XaqiHIQL
jFBSY8d718/B3hdJ6XGvc4+k3dQflK32o60RWu39ku+85lZpQ6rPjjbp9BAU
b3fV5meDAZY4rhb3I0AInMXyxdF5eF8yaZKkIUIyOmcmAX9y4LdhOSOcDR4J
p8r3oNEekLrhf5SpRQzSLes7PMP547irZ/RVvX4f0Kw9EP3pVPIh+YQ1o1tG
EDKrqq5juDjfyny+ifLMr4OFFJO6hAirG50bVxmIJoxhLJwS2xdYxvXOlcRH
BIOswFjpK+v//DVQxf7PMogng+jzJk/PgCnZ4Td1A1QnvUxT4cYgOe6axQQz
fWEjf7Z2Os6Tb38NdMywsq4L2TzNh6lhjN/FKh8yRItsvDE+FFajzRSrhRgb
enqAzk6nq2PM3yKMjH1M+YPPYIv534oQOewZi+KKfVyVdGb28DUWo1h9lh8d
QfSqidL9BoFRG2hQeEHJfzZnUDiHGMI4TaRmY/vkkkTsLLwJUH/PLisHL+By
nUW/ZN+MuY5iSSHDx/wF/BNPaPR6BdydjTuF1P4BpFE65GPheARX5aJj/Hsy
iufrYIx99ws7pb3w2/3PGMYrQHg/941nPgPzKUZ+Mp7QGDh+3K0Emh6xtbw2
EV/HhXf9SalEpKd6ssN9pAKt4q9W8b8bUD2LY7+ozPP0eLj7lxRPn+Ejan+s
yFRcEialI8xULx3KrX+uZF9VVGYPz3EB6TtX5B6mbqvLhbO8UkWSasw60DGS
AzGZ8abRdzVpVQCjvtgksMMXIOrRIAITCBoP6M+iq9CknpI2vOKcVCZcLtxq
SsuKlSQtbnQARCKLuPmSzJj91SeuWem4PMyPUKdQPXGgvpn7GDzEyz4lyqdN
ZDQxvJJSl02nNHab+bwGzOvxtgE+Yf4okyVzmAZOSVh2K1pT276p9zVVT384
hiKiyD43bNEs/4CmHMHy+DRMN8ONeInqJmFFdyopLmjqDXoEJbBQfeX+Fi+u
qiASrBn+rqDNq6SmJKjYttJbFMkzRCO4yI7BxPpnEeRwl+fhhTIhEkyC1Xhu
aFXorJbPsEa8iYEoQlvIN3Vl/8wdlbzLRjkhhdbvXW2z1zE1MRxp16sahbAB
ekKW609NeRhHb6GkPR8jW4gXXNjnTpvnqVgj9pwMIvTo58n9BHwpyw/925se
eqIYIBeYtgPoTcBJqiETlC6XAGNOCRicLqdvn/kec8Tx3LaB0VepJ0M/AvY/
nQKtZjNOFxVAbHgXbFZ9mCignwwvA/efAzlxfE2OdvVS4KwtcF4MuDl82w3K
8Xpq0mWKw4N531c9+n/jJNiQaVrsFjLCaJxl4CAisi3zj2HEhMaEbeFah7Sx
nFUs5Q6mQfnFJQKxEUpLTNkzO9DKI15knEqAP8CsIYo8/AkZLiNFIfbEOzJm
sq2khMhAheZXLlT7g6+lVdtaRRouM06q3dNbTP13wkLsqgKwxLdG3JW5Sxyd
j9TqjxQFRL317whbvpK6IKwMM1DmCr22+P2unqWJx1cVgJQ1fRZM85IMcJp7
hgwa5hZSDf38gI6LW7HAaTxfIhQIYocjVxhNBHoDMBaA8JoKl84nrsbi9YNw
blyJ5NAqxIaCYKHILkAlobBR3KffUwEl96w37jgHIdYatqIcL1sDJ06hgjML
1cEMYmu1ujeAo1v2Q7UN3CGxMBqbss/fyWOEolIc6tZawTjjiGMhjCIlsapw
qlOHHaRJCOpmPQiacEm8X7PWvkNer1xziZB9FxDS0kODWzUtAQDlapHE1D4Z
iJX2N6mIg/0YiPasafEKBF+SgyRDcjYaZpfwoiYFtVq2EEkcp2ibQ77sCbit
DKuSq/IxOy/1LkxTlVvTXrXjaEGWrlEzX9IkbHYorG6hV+z/DAK3cOMKNELw
uSYFj4kbrVrId9DvdS/KO9yijRlNAeiNodOC7ayCDjE5b7Tje9xkx4r7x0UQ
dPyxa3QGQpM3mk+okv7V7VD9i0IyZ5fLrC5vhWShfi+yiUWBj79MlrskVLTl
KK1G3WISnGgL8s8uJZvQYALeaFmxt13Y2kmra6GnB3AhBXdSdnaNWS1ROZ0k
vS3AKkBe7LF/kdUoQPo3+kYuucfgI/HUOMfWqP4mNzEcv9PnyPllUrzMusHK
l5j58ggouGkpjjAz4DCKWJRPaWHgeW3PxM7Rjb0k1h4dKWEdAXii3SNMUxM7
IC/trF/zGAzuMgJ2xNTb0e8c7k/goRnxPM9Fy1n0izxLiJNUPuc7E8j//XHM
5jLoK2k2M90iBKl+NNkg2N2KdfSrxngLOCkkR8HVW678Vl0k/CpdqRIIJ/fG
1MAIdmRMcCE8Y2+qPWlRj3aG5wkfzxgBPTbvn0V8a+AEPid2hbJADVNez8HN
Dp74RF8AFpQ1DJR8Eaztt7q+D5v39DQ3ZEbIOTEewGgA1lcbPcAEbZJVsjGQ
pABDokqcguXqsUWRIZchnvWH8/OxmB9dxN1yQFAR0BQHpmyRFdPow41/4q7J
sv8MGObeXfq8pOTc6MBQm1vYXEF0hczn9UP/cw8WPgg4E9zewYn16Kbc9I6M
MzVNmFMjwFTJjCEM8BFdHTTa+JMHuyT3wmQsO82Po5aqK7hs73DNUZ1PNxK2
rpF9fjN3ZhMyMHbauTeHkH5pBrL5dPJ2NAIg1uIVsS+9Mu5IiQYOjpWdEBxe
utmNz2rO0c1LF/UDXGjRfdYtWZYpafEmVdvadV5fka3x1G8YoHYfTmWvA9WH
jKKzOCsfULJqSK8yaluclSE9ryK4EKGYGw1Abgov+egq2NDh/f2oAK91aaNr
ejoqoAhyEK/iQxIsqRdFxHHg6HvgZKiZwbqAD9p6jVxz7u8dwe9xJtdVu0rn
/B/UVFdqH/1f4Gjey3xnAuHI0RazCzwcL+KCzwTkJiCgVUFTLf0zNrFzZ+qX
YdgWHfsQWtYBrIDVjvXYx1ahx33lYVkATwyqhwW8ioq/qbeaYo0dfHC/oZku
YMMPhVWZ3ShTORXxbhBrPdRJxlwwG53eUpkZy4Z/QTolZvRH2SbXX8uoRizW
pzPpnk/cb+/ZdQ6JAQtWhHh+jJdyRuRUIpGKu6FJ/EobbSG00wrv52tKBpVc
Nx6Kct55Zbvm+nGuGRHNSKMtg9men96DpxRx/vzqZiXnDQME30LF6UXwcbKF
W/0Revk+pXLo2pRYW+Oc0LJQZujF+XFMFLM/DeZ7xeCjzwQSSxsSGj3Hk/Ma
OKdjsxXNOfreKGd3oVQNoPLIxKtUqaQYh6ZQcufdxiuX0kUc306sVruNgukl
b7zKdpM4rdyYZ7fAHCoO8GlGSyPyFhHTTbfjx3wdpY+MRm5OgDRmI4kHzNaD
s2yqqHEiZGH74ka4Aak9QKL+OLR/cVJLIbjF1ZHBjYjUPJZYXTe66hRZ5Q7M
ew4Jr0fqkiE+fit6A3+qzQL1vc4CALDSxHltW3R2a4+IipCZL6tF4V+s0QUg
LzmUju7tc1AIFNHDMYbpFnwm5gvCUnC37wFw3yQy3SiHJ9t/c0GcZt/KNYD/
Mbzpj3PoXiKE2SGY7uspTMZNHbs20zEZ7O9GKqUt6708Z0ObqoTiTBqX77Uc
6D17uh9/nrgvoTpT8krNiA0MT7k9bAQzq6xGoFyp9fatXr9oNZ3xhwbR6VtR
QIuHTSuR1R4RMhmCmc7zsWvH4110AC9CKyurxr0YHwnw6vzX1TG5Bb62uYaE
GE0B5HpU1oEPlmOHN7xbNdM52Epdh/vgPu+hrk8WcSfRAg/DqTyfNse0nOIT
opYA6spBzKfEdoV15AeDgr1F7o1J7bYkfyVhQOZAJuYktYeFBGZDyEvV2sfj
tAWji5Ae1u3Gz7T5EoBB3DT0qyyjbH1905jmUytzBlazk8CHLuuao6ByGDxX
m3UZHe+1bqyf53GKQQ1lJ1nz844c6IMsQPHWVW5hTDGqS82bHEUkWVXOn2CA
OnyqizCSBPpvD0Z2gxMPZl8T4nCXeS0dbjhL1lqjsIah4zIDk4/ZfsBgSvHb
OJkUmHDHK7GAJzjsdhnOaF5GCN4uhsAhciIyb2GC6TTZISicMbYyZQK8cY4s
0naGXsHnaqK8Zr9khrY9AjDBAMDjFCaIIdGtpdsUrHPWX/3xcySrGtCksCqm
Nd8ecBBYtKsW2znkSP08sNZF5NLhyFqDg9lCDKLFI25je+tqzCWGkbPKr8Hk
7Mty6bOmx1BGYzA3n8V7A1aOIe/DowQXum6eYuKim9QZhS/7ErO0W4QBEsTy
Pztk6t/8wLre1H16o2ksNIZvkTyq07C5OQf9r4AD+ruQwubinLHy8ONoXHxo
DjVeBjchY1qv5imLLcJD2b1+Tx87FXvHDJ88vSS0ezf+7S/OndFZcLvAGDlA
ipc9ISzSBPOvauCca5dIqPgewkRf0wuwTYMvfu0W4HKvssR+N7o54JRH3BXi
IN8j6l0gNdsxagoAyjADn06XNC6gVzimuSXqLQ1f+Qidg+u860MduTlK002q
gafrFb2hrTxOiUIlZkjqjNcQull555acDi4/jamIzQsiaF54+j2JyTZRr8E+
SooSW99Ze9WfIaslpI4FGHMPg4uaqVjIbR4vt1fl6Z7XTIq4hU21omd+4dkA
DD0ikasFzdRd2t5NgzDEP0oNBZGQUgDTdC+Neqh2oInBuyaI+n37r/Kj70qc
KVLJzl1clg4wlTC4oBhLVSZGjeTptlHU0lQeObyOf351HNI4p5gP4L9z0y11
oa9v6zrbNITrkqDNKheaScoP/XlG3eecaLni0lzz1fz3j9+pmgtCjzOZFK4W
5Yd9uEBwlnMxDuotWXPSlUcm4zIlnTUlKSo0QV4E/YTTokzTAus06x+SiONZ
Xjq4a/M42ySwDrKP/GpMrqiiSvXayZxnF96b/6+4aEPewjk0StPomJj1yT4e
0kRemwEiMkeLsHlmBZWImrPalBMsVzf9ZGv/a0mzwTWj9gFamouU/VBfP0QI
bqTQqpuuX+LmT8HZVJ0gpJdpUF0kQY/WPmczqe6CmKc+zzpWo1HurBhaxTt2
m80Blg2mndTf6Asq9JwWyoOQ518RybspL2yZgXnLM5vpq8iEZur5o40wa0Ob
8SMAenNxqktR+lbE+pl7xJlBUSI1DvlREJlZfJfEJpKoS0dmPQ/4EP3p7i/u
ZfcnE/5gtRxGtJo0AIwJDgOVnPFBMTUd71K51Yj8O+mC0molfIx1A+/5y9wU
iBIbkNXeIqUz6GldMDRdcIsrV7blbJsva/bn+EcBgbkU6zogpI8qTT/qtBAZ
habsuxSUw67uPa4OC/+q7b9vPNMDOBgsaHUzjGx/mzES3oXfjJd8k+eAh3UR
SUtQV2SJBjroNlBfed8WaL3gglwjutve3hAiPgORHgGIrKx4BOvjIaUNH4UZ
PjQF6ir4ZpUqwAk0DhS+U2TYiYgffskyjeOd/qrhmVPR/MXELgTB0hLC9O3Y
xM+dyYMnCMLvd9UGb17HNAdpXjMp+az56a39qP7wa3d00OVcU57yz7uVq/wD
08ZEjrnfdvsi4Pj1bDkhJb6E9bmeaiqklxqEjIi6XavpwQpuMMVS1XQPPU0H
5aWQ1JRBd2tFCBB5mzoqGH4i+KHSHzLZiSzEIN/ZKsomOO/SJ7MZ37aIPMAt
seP6Uw+LkFozLsRBD5nu36RNPXwV9jLWGqgsyHShFATA+U7if+5wU2cc8l+D
jsMy9/1RSBNCfzmQhwlnE/ZHGfg3PbWsnjRRxW0Eg+ABn/F+uSNyHQKWP7Ck
XsrfxWUa29xYJZiR+ThqovFFPAxoc1BL/fz3HK7/GLwu9siMEBQNL6ugAY3f
MMkSHSgBKW2YPCMani2pWBH1jH/0i0VKaGKpWjWqBXG8JMPqSW74VoN+ckhx
0LsyZfX4mUmvymQqT31olC64xWJlkf2aiP1n1FG/eEW7cyQxq1fCp1gme5IM
vomVMDokbS72refFQzeCxF8VhvYgc+2qxclIb7XILuSiTfLXKkm9Nddk9dwu
dHjsrQjorG7P/OzY6A4A+bo5YGIyifAMICWkBAxM/9xpvHDBut8lVDp5C+1H
h4zxHb1z7e8dHKAj42V+bEe6FYrmQmzVprnuBoWrJxgSa8bLnVaDHb2Xcq8l
49qpOuWihFANm/T7j51O+ZjxrNmJJin8yu2afq9VhnCvhw5v4B5Z7GYVopnv
cq3mS0PJYb9rljvrnyQVEuLfize1AEu0DG5q3Emll+iXdR8+pEeKM+9WexOk
ZtPBjEVRIR/5yrUSBpLT8zaI9o5yIQFd+eeaOWN25XoJqhAQA7HBLFCwPHab
J5iVH3JBBiA4cSi7eumzgro4qJNwl9x/Cfqrbt2ItzctGd1K6rUgmju5Ko2u
1HP2yFIKSvguBJCs00tTadzSrK9/68pCFTslAwwl0ZcyVN9oxIfXp58ZGd6w
xsQc9xTckom5hk1s42N4N7TK96yT5+c+16ohne2SGWWiyNOIJkMRFMUMdiAb
UKKdgTL8y9vdlgpq8A5DZxmmVQlbvuWLISG0O+anmXg3xVJ2kLIFxSS4aU9m
HIV1HgYATIsakOArB/g04N9Cf6iEGTAyqTNuYbh6d0JChHUB9XkbkwZwD1Xv
d0Xkam6/WiOBm6R3TIjhN+JEJCHJVQXM0LrpQBEibCev+bx/3pP+eKg2zZ0k
iCN0RiokIccQHOQeIcq4J4XGI3xQQnFDAoXstys7lyavV8vpottWxhZQ1C/9
jOgyYf3C2lRWQrtCoenRCiJBTnri7jCbwi03qFdAgH/T0rTkhO3LRm2bLvUo
srAVmMlqp3be0sWORGtEkp6Nb6RU541eAxyk6QhxhQjCtmlWuDGVqSRhaui1
Q/NfM7O+ij3vbB/AmH9QDeQOWBeVruT4sX7fXV5Of/uyxu1MEqmDVwgzkfpt
N1twrZaIXErw4xrssnekYAxPaFHqu/1HEhgEbZxnRFzcbAxiW6JsMCytiPo7
SK4nkooudn8MHDl/plQqmbnMHgNUIrnf8HEoaMDUFNkyXlRpH5eZESsly3+T
xzdl6jcOwTBuYJmnntWTSx1gCTeMkyx/MGhuUtv6GVYw4uNAxyjnTk5gWv42
W2yHyvFmqSkdDq/SQ7HWTxWjsKdCEB49MmO+iKx3fSNtvGssBsDD+NV6iGWM
5hx+niEtxsNHOawfu6WsAghjrSSri/p2OCwD90w8b/ydiAcZmECv0zUu/azr
6fEbcOQi7D+zn8fXcBQHXx1x8Gh7wL8XASnOY0ScOcepxfxvrYF+E9/fmg9p
YI499XFsOaKWboXj2hcQ3VHeH+A+wtvuLlyGc2ljpPyFHbpQ3h0ncwKrGut2
C58/LYzFP/l8OOpw7+gpPjq+wbDAAanobUnV48yOhBr4G7bfQ1xqzTaxI7On
HTfRnl9QSTNEMb9mS0BSitAAtl9Iik2HKjDK5dnb6lTRrMw2txAebZRtQPZf
jXGIFva2NeaUwseUvMx4npRAqefeJP/BK2j/bHKYAQXGv+OFSSGnVtrYpzNe
E3NgzPfyDcuM8Ga6H2NSwYWrbvMPyMZ1sLNdkJ7JQS4mRzIcBkMe4CSYnTx+
KZ5S1kR1qPb/7Zya1O2ZrNrdRFmcDH+Wh8U+VYNhRHh6ExFBtafT6GREw0+e
tqmqPnJQk6zHYn9QH4YZ6WXtNkyt0/NpyeGMZ5aCuUJujtCECKxbgj3mY6+/
MCHlxq6fZnlvQtybpQdCV00Vgdiv+4OCIFaF0paMRrpuarb0vDBRzKxF7/Dt
YVJD/Ly5qBNC/PVz1e8JMvmieg0q23dv4fCe6J1LRAirZi9xgL+QP+NtS4qM
cUpXoqWk1ClAKQA3DTZys61jhybypIaG+hbSDZkKyhiNyDn1x4g/teIZ9Wq8
FLFjBGICwaMG/M608SDPRQcUUalFITmgBoeMbKim2IYthew4UbQuy1u90a/r
BhVgHcRQZLtiAmcK56Qkh48bGuzqeF5AivJtcdheQiznOL4XJazl7HZM/2pI
Csldlom6UkAFYordygYpln9kOLMXyCPq34AzrUenDKpsc8KKil45pNVJCvWq
oP/VsSBpuVvuErdCuL7eAV4ZMfQT11CV+cKf/Ec9oFkNwZL7jpp474N2/TP5
zpU5QPqhGCQ48PY+5Om9FiWs5oxnLFEiymBxjauPNRf9ilDj8ptPJDwO3nkv
IuVGImGdhUWx0D6ptAttfW0G0U1a+s9ozURxFJCoRIu9OSOzNQwR//0zc91j
ZoFEjhWDKK0APc4W3MLOTK8J+Ek7YSUjdl11dyVOxeSlP63A5apKfBLCjLEU
ZtLiLwOrIUgZQChmQ5BR6lRYzzbvlEDxBR8mLWZd3AlEa+XS1+KozOCEA9M8
CfzPEUEMoiCtECqCDUZTGrio8wUVKegzIdFOeV20jkHQ0i1eesA52UVZFljt
K4+tdMfjdH8t63GtcnVaNoUg59onXlW6ff/BMMOFVlKXw2YWPkNteG3pTJpp
V/6DMQfeMEKTSUYxQoXW106t8JaB69mgqXBSLeqMtO/Igj2P9La+3hjpQk3L
UbND8yHpSMuzVtNmPvO1SMIc0IoEglqrd8rks+vWtQA8GQpBbZFI4ty6sI0x
DDZ9w/q5IgrHe86LnEy68qWJ3zNePMViPsY7FFn95aVrW/JnLZNj7pZM/Gtu
DWj03OgCOCW34WPFyUbeGP8/i+XT1JhZe4xkCm0aud+EaBRCVi3zbo5vOm2w
1za/al9FdSUtKuzRx5OQG6XWOs6hmodmL2idBlTxoYFWRb+/SXfnmLyM2Tgz
n+O26HTqa+ENZDnUS6osI4WTHfhKj+Qf40sknqCWBpjrMVWhuUNZWuH5b6X7
dv7INaboIJRrt6uqh5jvEBfSEbxhcPmODsZrw6wovnxjl0ASV3pooUpSlBMp
sE4fMI8c3l+fRL16OT/Pi41SvQdAWg0Ni6Zsu0bJmFMaa6yaOmiXmG1cP6UK
cgbFTFTkY4B4GJZjXirfeFt6oTTSLkQMLhyoYXib0o7MQwKxtIxIvNpv3Chh
fZrJgcUGYJUdUvorSx0egiWjYOQRhQeaORrhayN8w0jLOebomcPudJLO25X9
+jmTd4rNUWBV2OKM9I/wUk2WboLYwa+He/MzvaG8LGa+gOzZU530N2DR/XNT
9zZebdVvOglpRiHdilSNoWRG9n2OlJEuTvST/W+2UWaRIbX6hyEPY4+ROtbS
vPrqse7ivcYZmSt7SP3ixDHYsGaGjbvyWvOGlqyJJrELMXYCBe+OiFykYye/
41HN1D7IsA9DpA9ogt2jFgRstMFUJmE0juD8+wwE55G99iit1DUGQEByrnIw
8WV688IIUODIYBsWi+Qtcwr5XOgb/Bbmbd9F3uKeH1zH6Ux4ChyR0RwetKVH
2cfTtBVOFw8YiQnI7a8oPlfTIK9b9FSySQYXMFk1yck3w3jcIEfDIsAZSij1
/lPyqqXFSK6rXoJvC5ka8At0CbfoO25PNvxnMIb9R4OZN38id5WumWDY+Nbk
9UNr9VzhjCAgo0W4j7sx9BOWORiSCz+kjI6hvn402Cu0xvnILZlwvuFLpqoc
W+a1Pl1pf0wfMyg9qINS1JB5G7N2laxRr6bHJshQSQUmstxR/uQhyb7mmsV9
6zx9Xs5P0g5Zbg+qeYgznv2ujPPAtCB3tGY9iAyf/1SgUQMIF73Yk200WiPf
ICKCjRZpgCUEsaoVq30Nz8JDHTMmpJx/7LYUUpWofAlAj3kunoUEJeUQ8rAV
eC3jGyT/3iu0bFKrNoziNSuHw/Hr2u5D/0BEbBDNCaLWs1PZbRBRQkvawMIr
75fErZR6KO09WxpKQhBzcncX4uPnCrfPtmZ1ixzQ4/Cs+LtptVoOKtjLH5y/
hTbuQXBBo5kY7qUSblIC58m4hAdaFoTSeI6jxSzm/qLwtfmzqPvwuHTXjsba
xi6DW6R8JBmM8FSbP1ZGksACK4NwmghDo9XrqXFWFqvpDGVrpZEhYOXBsG9n
ErBifD+Vc+Q1MxE2WQ1qw8ww1/7bCNSSsH6ch2stNjSscSCxtqtfPmcVJex8
2vcltA9nQ0BCAxsWT6rgO+Pw9Yljti+90xg35yqkZ1Hmzy9DT1WTZcffif0X
u3lzsU1Q48WtwuBaXBigrvUDTMVsls6qrjmY+2Wx0yR4P4ixSioH9C2Xp6Kj
zTrq1wBvSiYkA95z5UXrFuYNTekbLczYSuBoE1iiKGTv+9PlcGh+KaVZNlvl
fEMWnf41dFk+MA4UKHPuJ0HbUrl3v3ChkBENIn0hfIa20J7qwmMNbaS7Z2Yv
dwFVHLk0w6yYehAKtpJFYhOJsintMeBAVCvgXfc48NhE4HMlY6RiHCZDMuE1
rGxgsxVgtujg56zPzpXLXaikuWVSJh616IwWfHCEAvYd93KQYonOlRI/kAmb
b8yUehh25y5SnHFEhvonInLURqMkoLaHiuxNDlPMl5EQaecEZdoRsWydyOem
THTVcAnWQ9LttgzZjTHM5JjW5cOg0C/k0js62o4mTYkm9LfexS8Dbd/MG4Kt
DJRmUid8qbllnKbWLGKDjIMxjqSxsc694ffvxkyL3vzGR8Mp4vLli5Xnjm18
C6hjOjFpClgJCE1zQur6l4rljnU3FtBbDgZIb5+hU21Joieb96mAQ640gqpQ
I0oRS6drdhFIO23Uw1hQ0ZUAz3bDp7N72GJhxS6HhpP/bEkQpFhRfgvLQpSp
cXuV5/YSLRSI6pgsUINJmD1GynQ7GtssIk0451cHw3Kv9tijtAynzokXZryH
OMlww2qad6ar4CLfM3lO3PX7oLwxeAifGdCruey6hGJdOLVa5Xqngi6do6aw
t+msTxPAdDayQ3QzAAhgEj6JFfUSy7pS6RDCDsG1QciK1PvOcshXfOLxXK5j
toK7sZLc0W+TBo8pEPrJae+jx1iOj5wydzMB3KFXZsbw8LqQGksk5ECY/CRn
+ZudU/nnszGw+LFhmRbxV75MsJ5F+dtr3NGAoSeJq+Ec7+k6lvqwJ4o/JFjR
CiHtxAxgn5bpwjYdOrav5R3DEBPv7CWvXdAuq9U9bOoaCcK83MNzPc5h04qu
D0QDWfzdnCOyiWJxQoEQDl1ANzNXPSLTFirYjX9cNhqQYMObiTw0FYY7gOG0
7GYx+6wBHjjl1VzbGsRZMaep3Z5ukXfuwnVYQNLIZyUUiZN05U7HZ8W+gwdJ
M50e2bq7UTf53bLHaIbVxABR9GRbtxjKi/3t2npMAS9u4k72+nTFyvnBmsuT
M55xW2f9j/2lBm7tdXvOg1E6wyligwWkbe2c+y8jvWSc6Vnvw1JbH5W4vHe8
rMv+F3hyjXoFBIhJPDJd/neyCn7mJ5mZau6lo177Bg6WVkcni7+OkzCciFkl
7G5+SCeAQaGbcMdJomJFpsoCdrEZWQ27FWndInJRX7AU5STvZr9FAL0or/si
P39jST7E73CDjjbhDv3YM4oyjV6uSCyMZ4Dkbye03DWoE61T5/8tnj+keQQk
FPa0zc32T5E2S7eqfPsV3IEYnnfNbWwTD0I6b9FsmIjvTHvbhzL1suJcsymO
FkiHnAHG131OS1D7j9AWl4bRtD1qWqHphV7+uDO1PNEvXWMy24tg6zaf4T+c
iTaf6wDTVRKGCppWFoUcRWy23h5APLlAon1Acqxogeui+tDzjjKXmmpIpiaJ
hawEF+bsJ94OpZpuiLcQACWPWjB9XKQDjLm9bCnYwG1DJU5/KT+roYdRKdCZ
UESOA142mNuKYjVvVA6Da6rv4uJo+Sr1I+/Y4Lqmfz/qKF55fvgXUc4nDaVt
qjGR0rNdkUdzE6ODGojKV1O+SPss1olBOC4HrJiTltoyT60YMcnxrLPUQzNx
Whl2E36RL2OM+vyhm/0OOG6DOEqMcPdcm+lO/fYzAjkIWFlG65ug8T0UVSBp
h7pej+3IqpLinMyIWSi/WRGY31FvSA+7H/qW+P/R2WfVshwmzImmG7YfIgLL
cPuFr3R63EHVy/i29N/prRHz/Glu2pb/+Fhkn4XDm6A9nOJxvLXeAucpcKJm
IcyvIzdUskUxRvvRIcGk7CKYiUt7yh8l5yVEdlOxJ+f6nNlHy5eQv9Qo0WiZ
mXNP9KahT+/Ov3x6H/OZrp0zECBgBBWRuzX1BnqDG78abAN5crvX+xl7K7wg
J7bggopWWwZT4oh1pljKJo2Z8lMlSVmik3NbM6CNslEuHqi1lqWHm8ziqaeC
KEnexPTlMhqsEG+jvGy1P6xXXYDw2SzXkJlBIAKsKFXpU8ZhpxbcdjDnelG8
QSIL5+ppQgtBeXpUWuAf/LeYfhsvaBbvNa2Sm5oJmG9oN0uWnHg0p5H0wvt1
hipI1lV0e39d6ohfyROjYgHrcl8kE41izWyKzWmzT8TdumN03sQK+Izi5P/+
ZuKDgRmimIemSyaxgrrOoAarrd0Hv1scXdXYmWKDseF0dQrXSB7kWro4mGyY
VAaIxinhC3X88RVWvXRbIOeMFQa+vYtMvp+LHQzD1cx7vB0shzjPkQRob1Zk
pXxju3ssB5n8o0NRIgjBhyuzfqJw/5RKdVnZ9cJdnPT2JDaWC1JvNjVHoQyf
D9hn9+qTsjheorZoMwBxfvP5NParMsKdCbyTihx78OLn7Iu9Scx3G8LbviOw
GIjeoJ1w4tWtr5PTety+IY+ZORMuudn2Lb5WVukSIVaaHI/xJFqyXVoJkDau
6RJReNdCGEuKBzusoZDVC98LWp/5uXnKUgpY+IFiMLZiBAQZzI1INj+uG+hy
/TYFdNYCNmg3u9sF7V9xNADIWKgyO0VeJ16unrg+rbaBzgM4R7O9BwJvkvks
UXdfab2YG+6e1rBXWVs7SjpKq6DuhhmuE327V/tqGJ9u8DtbrSKxZBngBJJx
287dVy1E26NIR0vK8/AC20AcAmNLLd1ivOHMnuLZLJFvbW2ZXeL6oRihR9ri
8Bwv6gAtsoKYhOwP/G8BUR/ejld77RDrcEwN4+73wDb86a9IOJd42BwuPo8E
6TsI0FTx7GZs068/9RZ6oAdBtEpU904FbYr+JARaZx5UxcXbLaQviZPQjCqG
+4pIa23VNCidyXvfel97F2Fplf/cBrtv8+EE2YlVWlV1Cm2RAG0RZQ7gRleO
FT3jxopw7DTAQeHTpKlSIoUblPoOb2brwGREv4U4xaOVMzkrBLR8OnWqHVaY
ZA2NQF1BjM+AsVr0gQsNhsW8cT4mutWwDsvdDklO4jxZi6xiejnmf+Je5jaf
fxSbhsXbzfbz/DMVFcl3DioQ18d4WjCCej118qamAJ4EpLA8TlvZWsqSkpwq
N+xvChuh6VPJIORTHhbrNOFDfBuzuMIuCxAJgxYv1ZvqIu04dT0rqCtwSxGQ
d2Ndj7EWU4z9c0CIfwch9FsMSguYQ09jgynRswDjw7edMLG5QplCo4CWIhys
Su6KPHd2VFzXPoHQn4IhZts7PPptdLs5Z2e3qLX/f+RibgxhdKxZYG4PacD7
lYHKOCFh3dmyD0Xnp8ItrTokzV3qZdVeHqq+CPuG8LABEDApOgxyjWTLWKWy
APRKiyGmiiUFHEc6tAFV1epZi7DZUpppsitsd+8grOSO4Zx6Pnhn4hY132DR
SPrEIiill8lFJ6E49/+4X9OoAWaVqh60OlLpgJmgdGkV0wi/bGjoDbq5ymFV
k3RnUnLEAjTlyYV8wbnPsN3yCoGYK5i5cN+RNLq1xtiRRPNNIy2vnmwXRwi1
kxxt+q0QgQ5PZEryuJjLPwULxCqB66FJQRKI8j9pLfbkpOqXmLMxdBuhtLIZ
8Gw1SIeeFA/6OCHhhv8YnfYFZhvxl+RV3EjtS7Atbu2zYDYY4dXPAy3trHX8
icqxzo4ObZ4OwCBv33Kv3nYaAkn7He9mc8JWvky13+41t0FXz2CHvZ+l/SKz
Afx/YLPxI3hkL+7AkLAp6M2hwBiRtICeQxB8nGqkV7zwHeUJGAknDWVOEMUY
BKoEBhERCRTjt4ZWX2mt7sWX3vItZnPtRp9yKpHInkR+qdQb6JSdfY+PP9nY
uo+kEEOjs3i/fgMcqeMimONWxsP6hw26zb6+DapB9LjfiAK7yO5Skek54JbK
B+2FB3pVGtl0GVugw1BsSbG9WU71ToW3ylH+lmpqFcX9b7asZ8lZIBWpT385
U1UXROw4O+kKXoGdVG71F2/VeByKlXdAfmYFNBrSdRgP+0XftF8wZwmy9sIH
yWpjqsyeq/H2rFKUA2gGpA6KNUQxu7QOBnsdOyKJawz0XBDgzsajJfjegm4e
Xj7DxtFD22UbMVkFaR4S7Fp3ZKg1U1IF8WDOdzDPYvMTN1+/xHO92i8U7SOa
RXn/NsmvfyIoUD4O0bNPvW/9qndJ530Fi6Pcj49XBzXU2tNZoLQiiRMHLgxt
7f0TljbAYmekK52sPn6BgwHJbfFykQ48q+DR6gUEg3G23u/eBW6sUhOpeUpi
BfVWyM0sUpcjgZFwmrhtZ0+a+Yyn/ADuEF5n+LJ8KSp+FsibfqnVxjldDbQs
AunYZt3GVW9P6pNVG/MP1fQ1u2ZvSLdn783w/4du03Cbo73jXKfUs+JFCGxZ
eydb1WJ81p16nomdhUJ7O63z57tvlgv/q1bdcTvYdEXrMZw7gSbuGQ/J3SaJ
OkTrxnEc962lQ0/419MyMlThCIs90SH5HlZP4ylJCQqQgoHTgcouO+s2A5oK
G9j4BS29irYS8VfVlxYxoMhRIpqCL0m1ppSUHZCvvnicHw2BIk3G3j9eTZK2
tbKjo/4WbMSCnmwNObMNR5++MLG68Vjc5wlW2NiQDQgqwH704RchqLldT9xa
Tiac0RowXGzfUk55LeDqRDam3jP7EiO80eiCkKOLsB9gnwGGSh8dvvBPpvK3
fSFkUNoMsIG+GWjxNZvsS4BWzOdGG3JqOjjJ797lTMh1Y1kEcuUiAs51e8Xn
NnKPu+WbdENEQvZkw79PULIW9ieeQPCB70bWlVcbwGxB38zeXvzZIkwARqvp
Qby1LMnJm5QP/fT383C41LRx4W7jgdDRbOtcepM9PHjZhYtbrDBvQa58WSR3
7unO5btDMa2av4zeK1+eUcPMEiEaJ7ypphXwviclFJt+nGwTosMMm1jwMHD1
QvEgHpJoYb7daOdKOgcpjMEwpVK76air+ed6hCMR/89/hpvh9MhiG/gSQCHE
U91/1Umn6tMOEZjjtNyY4kxi+BLuxs/0BIwmhCnSeScf/slxJvJmNlFW4EqN
nEm/mB4KqGgl45ZQ9YlZqXMFWc5a7X3t2EqbFI5+AnKXbPfoYSlYlrYZshGi
Zn/Z+qY9z5KPq91Yh9xO7r7Q34jNqMntGq5E2htnkwE73w11a7oiD8Zr2M2R
ugKbcKy5/tlIfleQe+GlGfxfs47xSpWGvNJgoqM6r37VzJ1gLGBQD4/qVd7L
QGn5D+20fuH5B5lK/AHnxAKtlPwI7g3lOSOatWi2345Dts3LGfHNEAPLCcVW
h6Cs7izutnc5me+IRaAew3uI8PLN5Jja2g0dh9wUAUVzo1PM3fS8HJ1TZmnf
KDiMb5WDQLWoJlUPJGrJEKJg6q/Wd+CJlkRd1cVvfx1HhiELUnqGwKFy+BCV
JMRN65CsUUX9z56JfWbFQ9QCgM4rz03CoaQ2Lp0hyq7S0+Kc2l3XslYV+x4p
bd+Pzz7MOkZvRp+dUz75XXQwtxIZLn9LfpJZZRyxIRWmgNvbBVsdRr48ew5G
4qdUD0oJ+hUKJHXmMLYaPXoxqQmJZMUCnmt3zSgI4vB6GSitH/ARiY40Ml98
STywsUjSBr4TjrnOdRB4VhqWUkit2rhJPCinIdjIeQGIsN+0ZpEZ6S5TtprF
ca6bslMQOYTgwtnXit5u2GWWZl7ADCqOJFX5YMnvHuPTRJ9QEOzesucIKWfc
PkdLaANG2ftPTE9ddoQPyfnqpB766Uc1qedpe5Hge6Y9TarDAPf4mvgcJbXm
f/oIaI7EDP07VSnAveCY90XIwmqJmClIdDi/a63J4s++x9COy8ntEyWxDam/
uTksPl60wPsKA0touPBV+YOCTYHl3WhkA+QEPkj1At/iZFdiFb18ANdiWIRj
W11rGLfKXCjhjFDI0arSQLfBF7hd7ucLYT0Fy0RpB6mOLjOlGcArcmIwxmhG
feB3C2R4QiGoLdTOerF1LNvs+9VOUcjDVeERJroRepAJS+eVJtDEfN5RriYQ
5zUtTEt5N+8j5xxuMWZ8WCqgrgcFZnGynZ7x0PsfiDQH4XPslkv60QA9vjEB
O7YWuNf6wY7PkvLBFCQzOPCzVNk9VkT+u2oivXCRhzsSWxHuVIZn4kVp1PGO
uwBBBihe+oMu0AXkgpA2n+EQHgrwM91v5q/AqRw2r16LNeDdXRLqvFmR/2eo
+y5o6vdBk8knLfQLnXGzQqFpyqvrn7fqjuHnmaG1jNH7w4jV0sey+SSrlawF
p9hF9OpAHmeKMwaAZlhRo8rrJfX8+VHDyq/F3m+YHFmw1Ag8KiYK+bhWGJ+6
BX8dp1YcEj6zy1NVZbAvIiJkDsS1yIJ+ZNb0yjmqEFg8v2ELfKGNlDnlApXd
3swcwDlDFdN2jmYsnLPGsEs/Xyk2wpR9kJmL8RdUzhpOt7lj0pR3tS6jwv++
SYpDGmwRogM4oxorpL4kzLBOJdKRIeG1SCUWhsYdT+kQLF8yEqz24sUB63m4
/V0RSkVuiB+o1xYXotlWKoiTfogmuGvF3LGY1G8zR/KhEfJ27QdKgoWxCV1I
vVboUeeM+ZXTzsZ/s2se47zOIliaNVwytzdk1CDGZhA8CJWEtW8jt8/ffyDZ
DuZRkhOPpMtuCj19rFKpHgsDT2IU4u6RMTfCfcMevzlihjuaNSVtWAtKwzbM
lIAyA7/o3IiSyLRCTKtO/Rv2Wo2nspTRtjRdMmVbUXCZoEzlfr6aWTIAlyBA
ILHL3nMvA65XcBShMCxhdVtdk+25ECc6uakQPBP9C6bnahGOfnFzswDqXAeW
nWGOgvEUamgAOHkXTH3QoRfA2yHBE+Crnmxo6sKeRganlmSrFgJ2gSWFifMK
0IrKlXpVvxFpM3hmjBYryLepcqKtsM9+IA56FlHlwkZSdVBgyPq06BvdYies
eGVlenhIt5oy+zRKTU98QqOzxZBM/HPsjtC5VNwh7tBpqzxa/s06NNUegjS6
m/m/n0Z6u56UL+6iuTDcF2WIDdZJ3gHyDy/qnMzBg23KgxJEAXRB2L0SvLPS
doN8l3FEHNWFuZVK1/cFF2qeXcHPX1T6AgvaJizQjhG5dJnaAQEsNeyFY0/1
5rZ3N8OXg1ZZ4/DKNAL/3gBbOIjrACOvYae0/Rsg447xWM12r3+WO/k6+J+N
2q4hgjIm0INOAgyWxo70YYP8P+ejXWLhLMLBISQa6FYIsDrNr3hUsET6YOul
UneCG5LJTxAC/jvSfIvnlL9wqRcDdop3gzJTEfj4f13e0diTnb4lPIsYkYPa
42PlkqQNQR+pFK7f2Q+C8Rf0OtfO7sZrH3OKO6rKJ1pOnJo2GG7R8IuNFsh2
6W6stCC+NtUCn9BAl45k2GAVJuAA/4XOrNOu7IgRloW/ZIi8hBoGPz1aSxPz
J83305gtT/3dhhjlvjav6S/tAzlrBeyAD/Ri3StwrgPozUY+WULeYHah85YR
KviYMZh0MG/GuoT7VngeCZAcCK5eF6qnnFEFjSqCHKX2wbxsqHyW/t5xtLw9
b0CpJe8UpI3nvyU0v+bAnxsk9B+zr9s0gd6YalELLNfS5cj5ciPWD+j4a9je
5pB7ixuK7ZM6DFPLzYoJdBMOhHOTtave8vDyyTQj0cCDJWknbZYZNaxw2/2o
YSEF69uTEnI5aQz0i9cj1ompUL5PKCKoH7+DrihI3ZuwuH84MA9o4tVjJRbQ
Hp8qd+nkrqr09pZiLop9yMX+bdt8ICnc36G3bX3BFucz+s6jK5KcEm1/Nprn
TKRyLNlhEHgm088SKC0mRsbxS+GONajz1akndp4c9U9NCqXgZ4F7oBrVT++b
cRBcpHn+e1bdKssg8AARSt+QlmIO7o8gQHd3bT9pNet/UidlFawn55W+ZM2t
Ubtm6Of+WNHfJTR2zFd3Y0bI5MChJlA8DDys7O6ATTvup9dcRlPGBvQOK2iI
hzgACIGZVi3mvTSolY998MI2ZO8Zr2zZsyO9of+1Hk7ufnai6OcnhLADWFKo
pvMW1818Y0MRi+pMYFLlt1cc21l1/8BY8z6qsTsFI/iuygYgWryOL/0Jvp/z
0e2DH30iGjvOAhPPVK80x5AKtrWu43izyXSs0spuUsy6I5Tn+U6spqivyAjo
oFaO6Fmfo47DSqau7wNArAId+/O223WGuaio72bVb8Ei3U+sCcGwcPR5K1Ii
QT8KiAjYUWoV+YcXH9n3oxi/TG9rF7HDNar+b0SBeC1xPr236Ry+FwaXSLPz
6vybO7MWDxBlhSEZTr9ANTuNuM07kVCNhbDZRke+JvN2DWLzXD4Yo4cbt5R6
MmbHyBUrrKP93f0lZYTJV2Fd6yHxfbdnsKllytf+FlE2+GmnPn8Tq5rGvHBW
mQF69UzkYguu3udWQ3hiMvvNfg9kCiLv/Ov405Rw11D3/kePJ87+V6iRC1BM
fI7ptz37+Jy1Tr49HZInYQzPpFJI//L7BdV02J33RzlIHqXtxUZTzT3907Ww
Xionb8mNVzNbhgLP0J/RpaZcaRsVzppUKfe2Zz6iIzsvajHXhQEDgA6A9c3d
lTy1R6gJUk0cePvfrbcsPs2Vq3h8rvzs/cbmOFQlGeuQlE4R/qk4xmfG1Kul
M5ETdPfcEir+uWn1C4WGqhuBgUwxxS/AXgnnJ6by8oWJrP5yC1gEYeUuDjIj
qLnl8itg57j2FbDm39SEMv6+h75WGk6q6smH9YpJMvlRpZcSuZZsEMB4eURp
NvCPvhmIUdL8QETpialyErXbpxivAVaJvIKwqM/uxPbHdPizwhcqH4MtM7XS
cqZC64+ljjGfRqex0s44iOrqmuMn/8QPN3CrX0ladHJRKU7X9gh45HUwDPaw
26C7qp4ZgNDASzYPxHCdmxVnYn6qwTX0nfd+5s6SzQR7q4WlaWRR5qH16a0h
7qa/rxcQ07vtZGOIEygJifd/AdLt9sIBzRRpmMGWIDcb/CyUtCDC/ijJOkIl
X7jPACrMPq1F7tiO5OVB5SYL1NP2U8kFDMQhUMgUC17OdMWwDkDj+L9TX5tY
c5FapTP0OW1ziUDbZCX7kNHKttGKeJ40+Oqyl5UrLsBn71AxbgZBsKX8OXle
ESNXJG3wlV+Apl1cmvIoHKogRWBghkwPYbXqaTlYGEaCuWlkWyFO/ancF4qN
CDTvyPXp4ujQwRju7fA31QnOt1UsSqq4ZU7uYzn1Q/f25PREoD6k0n+wSGCN
v7KzMnc7iYScXOIVVht18mQY4BLd1g68OKwNCp+SvQ1ICYypzE7dc/V/2qMJ
dpmD2ROGyfDmmbwVLCOnLxnoAQXGtSWE3p1/Jc7opcOQQOwkRGuwPL4eavCd
m//rRZWX3EWvPRkMadHkugVj+dg4DqCvhr9QgK+UeRoyTZiLZMVsOC4HEmpf
GEEZifHKMA4rSvUQ6BSymvFkPQE/WIwyZJ5u/aGmnDVBcDAExTf9mUGrevq/
m9wRv0SOnpxfYPy5pywf9sGJ8sgM4ytS1bEue0mtP4Osj/XRJDubPl7bXE6d
nhYt2h193dRa8F+XQfjj1xj+9CRCZ7sRGts1JHvdw/dby+Xg5EB8wxQ4FnxR
6/NaYmyHJR9HuMS6deWFc/miH8nZI101BUS5xTrrp3Zh9+8vXM67CNOcATem
3S2azvDpTbgOyUnxX4tpVwTnaBAJgx97lbYRaaGo09VY175XBVor8DB7IUWq
ykWVOy9ChQxSqzSh8Cq7A9F9Io66YgWNNqOaDSWCs2KOaGPnEp7Kx2Yskmmr
j33qNRX0zy4+i4Yt6DVZphpoqdyGO57w3hBhPVbbm05/yrXAR+GcpIXBLpZ/
bQXzhJv6KTV/+9WQOQbLJ4KKzLtXNV48V79litejH4Y5hqzPiuWe0BaA1hzP
mmjj20hv5EF9WIcIaH2LLbqN7eZx396YA2So/NzyPbv/hiELFqPpreZtc3Qy
u+HMJQlWX68lwY+dcv//WRl3qY3jaarP70ltPrLQaaG1NUMMoQNndndcKrYn
v96DihtJuDVRHlQh5FtjB7eCLgCUivv7v6Lk9R+V1Il4VNAxGfHS7oFWRU3B
S9zFToUW2JtqI82o8nYqyQUWvldw/SMK4R/OBYeZLs8t6rYqn2M0Z7KLPKzx
kcHrW1dk7+IBaHMoZR3lw2IXerEAAJ8VOFqYqMMPot96vAKMA8NCJ7bfkbIR
YWTq4Icq90zj0KYUl8t2bFiZGf22uXmmb3aiVRsvNTwunruKXQ8Z6PqDwLv4
DiqBqyzl1zehzm7iRLIO6f7OqdiZ+9ZagHoIFqKhZigY+oVh+1kQkQpyTWS4
Nex9yYlmuzxtmEH+N9tWrm9Y2iMtpcrxOnQlmp8hjG8EkAwR1nWF4TZAmazt
VeAU4RoZtwB3ci3DHZ0m5XqgB/a9JSIeDOcSdYg5c1/R8Zsc2ANFPsSdHYl+
r5ITLZ1mzL2brN46SzCxHq/N0Ai7/sQM96a5nL1YwGare2LRa9eNT/jbXVEn
o8GCiscxBE5vNDPFSm+tFIr4QqpYLTKRebSM2Qc6pcUcHxhuIFvhbvcBJaT2
2t3UXb5wPXc+RrRF7KiPpd6bjWXHwIXESzATVRx3q7SgS4e4db41Re6oK3WV
euKeFKxyxv/hajIKXHE4D+JSZJzCU934qZEdpze5AObsIusQTzfhQmI95zrt
XWpFmL2OkUtAyzAdkKc/naJzdjwA6o2qx+9JEWDAT9HcyDhP7g4ujO/dacLF
XqkyVd0N7TdqknN+OGyD2cxWTgccdkO7IohpV2C6A1qJW/Z0pbctz2bihAuk
JZQ6iGR945J/4016kletzkgx30q0ATigJZWOp1c6PH/jhMDFaHtGM+L502nI
reS41CqZDiojrmWU6F6eqENwWFt4wCb4vfrx14L7/JChQdyFKRwZ154gH+HI
cJ8fSOfrMMsknMjRLo2g4CINN72b7IrQDtQZVcwGPBL0udbwKr57KBp9ayWL
oldRVnG0PRBgG7dlKt8eXzzubdY+L0PNZ8zo6KT4xIfVRZYtnujeEfgp3R3Z
hiOdHMdxEEPXFzV3WBNzoHdrnlY8CC93hi9EIRKr/4IBobCR/z9ZZ/S/izRn
0qRoj3iEUzvFlpAIhC1HaqBaZwgYQB224ZY6lgDMZmkbtpLWi6ofDrh46Zjj
jdOaaqtsJiE9VJyIX0wajKr8PZC5HZBvLJstdhrSRpV9MsMHRPxjqz91C9k3
T/DEr1AkuMlpJWuJ0CEy1+rCoemkpcJ84IZQIQpGtcsNZP2RMXwwdiJgIPZ5
2TTh19fYHfbhfAF8FSEWpcLdi91ixJCZeMcq/G6pXr6d9E/tGrTixNz91ofa
tgzLP8yuxgdSLCKNY0Cxgh8iAFMf6jRbDUqz7TZpk2EHRkArsRm1Lt9UqV0s
1hfvdkIc9zyjh/qjG8jQ9EkzZYSTQ/W2DAQJZVpnFOP9oEIMgs4F2C9u2Evh
M3TPM51H3ZDhDJOedCHfH6++1b5DjWadgXEAVcS52avxCj70YU171p33O9Yn
8oVQb5YUpgAoDiRrlVIjFu/eNBjGkGTnEmcccd1VmHnf8Hmw7NCwy1vZl97U
CEGvUSSo5eaW/t46RETcaeNw1/tiwkrIttzGOaiAXgmanKa6vEwqWnc1YAbX
E4Dogxzh0erh/LDwIiXUGFMppXUOSsRnqm7Aq+xyY9nKIWJF0YQSKxs/2TXC
eWB2xMOoV9rRK2RwcjnstksYX9S7xSz7rNICeh2V15Ir1c7xMQraq3qU4Wde
L3cbkElDffelap4nGW1hohmEw933OohTZGrD4QFaKpE8wYO2NJUZ7JvTuBIb
I/Gy7m/LY9yQurtfbuRY5y3QPQMJTVJejnok+pSNoYqksRGF2nMrd5oVenOm
Ituz8x6LQ3if30hxHiUoCblR4nHep4VLK2Isf85GouvMYzSD5C/JXqmAQ85/
Dla+uO1jQvVa1WMQlX8aKu+7gYd0Jh18Vn05gfDVIKxW14q7WViRY0jvaupw
JKm2WWZc6r4j45+NHvI9C4KPCb4QxmB8lPs7FlXirFq2COCsB6ziuQePjWsu
zrTKRPPu4ZP7ZZOLLErgo2OoS/tzimvUHZ9e+CoHLN0DcN+OaSyslNhsVISg
GXcdZD7K2s8vdOSGXbtti5uXR4ao2tg2Muj1OnUbLnlVzSUZBT2eS09hUNQ0
ntvOxXhHzShjDtVmgY0DgNM3K2FfeQQairY+39iEJk8asbDoTvliN2H6H3ca
in7NCcW415rO2quYbpND+AeeaD9dX4vWq4DAxSYcZb5kMUrMdVlgciDIjetQ
mNJ8YGdX/dNzvzbka6NCoAK2L0UUiTDA0mSiDcFEjjx3CSQG+OLX5gHSRmA9
GvygrM6vhjQpmuCzs8Utk/be3fZLJ4fB3AjUK34Bdyiir/aq7Mip0Q1+8vjY
RnItcv6hfwQOLdHWrYbWW8660b36semnOiVkmCjRqBSgQD6m9UQGpchLw+Dq
mn3n0BPcTHKFNvhj+ss2ZKecBYybMZ/2wopeBnNA0ongr009ITXEFmyYfoD3
yshUC8TCACcd18sxCB6e3v/JjYRAnnjW1F7Ha3QvX73eRPW6NbnXFkZOJTRf
j7AilaFf6cK3o0ateJNFC14FCybWLPxME3HKmNU1NfjvD6W1q6QCw/+pzn4b
P+HuHCsjhaKa0j1SQE3+SRznZw1vh0LWt/WS7V+HZvhH/zH14IryqY8wSwtF
0cI+NHJn9/yFEaTuU1/uCXI4Sc0H9t3cnztMfA9qDxGeHUc/WAtduk1Czjx5
wOp6Lw/2iTdNiQ0nDT1fJ2Xu5cf4YTeuVtpe8PcKj8epyroKY4/yKJn2cZGG
dGYdxWRaqUvtk+HFDsFqDTxNFP9H37elaJ0fEcGlqOKjQ76bmJ0YRfcIdKnv
tOzsRldMbbe8v78KN1woYXf8jGxD2DTd3ZPYcJ90bmQ+aGMXeEL4QrVjRaa7
0pSk17zeWXeZ8i9rFh08+UvqpgYf02lBsHJjilpCxp3VBOlh6knu3/IeVkfs
Q8NYFVYPMnDaSEQZ4+r7/mAhqeIgXPwlc6WRW1/8Oxy2d4nAMS+LzNX3n0cd
jfMVIg69imRXVtGwGkj7WWsbdnq9Ry0AL8nfaL/S5zhcULUGaRJ/d2gJ5PWs
hsPuMjYfVOL4lgf+zo++eD9NswPXexNVN2e0gCVmZv2BTOYRD3SZfH6RM/+m
ePLY6qrkJfebVzJjfTPUlZZFoPbtE9Bv9XDbQAFUP1MxiIb110QgwT2wu4Bp
ID/oXVdxYLQYUeeUI1pQY8jfd8H0NI85Z1trQD+OZYBYfJyBwNEdVl1ywdaR
8zzRYjbcNMqq2YLT2lSD4CZfwjQkrOtHlkJQ+O17N4DOqGY5m4i39Bn2aMvK
NyldJidTnz+Xl47Si3L597fu2qz7f6fNQqCv53BFO4aHXpnNbrjQbkhNAJYf
++uiA+ywDBuWQCT/eXoq8yMcb+7YXc4DTghb7yjEkerxukxRhRk4gCcT6E7F
ArQn+kPB17JzgGSskfXEUOHOMOw6flxp63zAHsnwl9oiWMqUAR/eVeXxO5CJ
J2rqCR0Hqi4WSthG4TsvjLtgskzRIDTI0kJuZWau+PVrmeVb8KcXAGXec3co
32b0FEjv0g/ty02JbpARBDKjosCr2WbsUQ5pgCPyBoFsNRCWBi1UaVHweSTy
fkaSG+te980cm9SItTlgZTnFpNd1mGgHdFXfEo2hgsOTl+TWiqw4cdSzamfx
tNK9bQenkFpcyOCJFkLhM9mweAmm+eBSFkL+tq1wsFJIMRI4JrLc8QO1L0+r
o1th9UoT3IuTg3YEcBqVNzsovWWiCuG8+mN4Hvzr9z41Ur5G8u1jwtfEw8wE
J7JKZKuxvp7psMAsAqGafs2ihJmNc7co4KNlf1KdXZPomErUhyHHvSjuJwd9
CfFpdSIcOuLYnA8UwzH0KR96y+14bnTQVcEh6nassR5cQeW6lN+dhhd2dDvF
pEbUatZs45UoqsACl2fNv+X9wV7Ka13IujacMCog3NJ7m+x+rQdSvZwZN0W0
mDYi5u6sW5bx/MCGBW2Qc4DfYAyxzkaa2iYXS2DrYQn9PTcsrrfU5AFb0qIz
lUVuw1pT05exlOucIm8B0l8K1jz4t2QGcHz2CMkA/auOh2C5Q5JKnYAjbi1Z
UPIV1oIaUmPOdna6oZS002YIxlOwwEZl+uFrsdVOwybr5jzY2LfahP0SSnoa
Txq518gNHfOiMwyZ7hsH7LQJ9wAMBrfKBqIuQh76AeFvIwuIjEHBgpK8Cz3W
JnxdQDRtA1zLgvusQcKclisXWo3Boq8QoP6EfyKDs50KItZqjFbQ3Fe5m5PO
keJt5NQEMHyYrFYE8nkLPmjWNrXTlkhtPIwRp6uXtbXvv4N5Na29uXgeSfed
WOeVPsXCzz7e5+B4MQn9T2j8w9ALa9uWJa33RrCyCfTJod6i7dQLi3edUjIO
+DAZ/J5CpnbLgR4GppOdXmfpghk4tJXuW9EiOQhMyTCjq3kykXnVp/MV7wi2
XPXjUOU92TZUTtOvqqD5B7kmE/z/QvxbK1isYj/Nu2ksRSbSFOAwQODtYQ59
W8ESIwpsrXa5uToq33LntDNDyVv7Nv1F3nmG4lxlsS4SCQKYqfRNkxuTXweS
ofgAGAfoLCVzvN3dUt/p5+638kWvurSa6ag8h+gSN4fwI9bFOuX2bCqFy4dl
z24l+Ag9r95dhyF4Ub6a4tyeXSyVzYohaU7/vKY1E/VVP5UHRSQiNnxXJU5D
Lq2IFf2ubsybMVtOC4sj5CBYiwvgGf4fCZVfsN7NrAJwS1hMlwRTGguD+M6Q
LJDkYX2We+EnhLrVmizLlVVBjoBTlp2+6O7iVX4yVoXj7asPhfWAHqb8vpIJ
0ZHfTGx7OTKASBi3HQLfkswqSHpY+ogpq1Y2XC6ye/MgeiC+2GY9duAH80sM
Wx3kgzYi1uZeJECDZQgSTu4L/RwIoVkSYCwqCABS10cy/syQuuSp9REwLZnZ
4b8dzRirVXIqC2ZF71m0m7gIRq+L4zVbG+MYqIFfZHSqlvRcByy6kxkOOVPt
BV1CrRHKFw1lmOCjiEZZFki+J0nNLrFLZlKiFaz6WSiT4W5iJaH3rtCyWVZ+
BGV9IhuVZk9X7MXIPN4PsYdCEnc2Ff/IqhESBtjiJyNR2OsPEKnf9SiQZ4cb
/Dc+rZEo+JVpjx2wdtIda/LDZlWcMe4C1fZHc4XYQx6yMIfWl66lMGHgBCGF
C6hGJ3gRp/5RJVzm8gOM3pKRrpl8d4rhUJPseks9VEV/Hp+ejxTyv8LJ6RLm
MGsTOkcOsm6zKadl38PiRF3gf83tku310aPm5mTravwQ1gjpIrQVSfX7A3SJ
frxsQHZ8BcD0Vn4HKTSPoVWorO9EhSU8okkZRssRsqfLOyWF0x+YwcHio6NK
dvF6GA0H/iSMkEpKpA5nddNi+jKN2PH+SK/kvy9yzrbdkH7zX58fZxwqpq7q
DOUPkkKO20KBs2nVtnRT4bh8mx+rFH/nXY4bZypb0wRtmEanIwBGbWzhz/Mf
AFyIV9GqYv/FdL5IYVMhtVY7kgU7TUyzyQ4XPQiEyx23Uh9ZhNFnjNdaHo4B
UNsiYlGufdMhjP+AbCh8CdOVvwqEkk8ZVVaxU/z7/ePMEQAD2ffBKOIC/0TQ
6G7sPl8p4KbqMx9jKzsqToBItOF8bIXDbJpZczP8sqWM4v8IMe+puuyHaMF9
bk6fpjHgQM9MKiwcbZh0ElauJqxxf0DhL/+9z2VTcZ/9Nitfcgy4FY4pRwdx
6sRg4pyHoJUcAK7ISMBuRtDBAXyxpfaOonKWN7YD3Eg5EoU1CQfL7BUkmtEF
Fb8CLaXuxFsCz1zM56SIa3/o8A3MKgWEQgFVjCkS0YOmGdnlCxeHNoaj1tNv
UEChyOguQd4cA5niZ9JcEiF618SeQe2TN+iLuC42U8Hq9AlcVQwCQJzA/aHn
IYQqgLXmRRFNPzkTuayK5eVhviU9Kppco15js9mvoavDRuqdCqhCmlwWKU+O
bDfLTUwWNGRLmP+HjE5bbJI0/2sOfz7mwQm2R1YsrsoSR0++J7fD10v2FXfi
J0i1LBlbrtDdhJIBGBIgJttJuRUIAsW59RQZLHfoLigtjrNG1pYCFcybCrzw
l+90zyvD8YCpY0FLbZQOHNmEXcmsrD9WEoxBXo99augeAooM3p5WBTPN+Nmm
mpkC52K4mjvypWyPkJV1qZpU6ZPzkD2LbpyDzlIeuZPdKSORC8TZdpmnjm/b
ba/IXyoCOYmIy1ocWOI48PseOQWELeOVeoKZJaoOa1JGkQaeD5hqn/RZCdL+
u1c/3vmX4PrpIi2/L5QXUDMzc/D3wi4z/FpQV2IxZ/amuNZr8ABqGn/Qa17N
P/cj8MNyGN+Q/zuVvehwxeJv7Bh6usKLZHQuy8WF2p9UU6n2jMpQlbEnlQE8
hEZA1zQWPyAKkfRqxa4exQxQwe2h0ZHIaQQ5GWUoGwA4+MX5G+JEPZvBbdVb
eeauxoW4hKtxwFI9ZGI602OhZUHML7zSDUI/UFTeZq08TD01ORcwFlJfoeX2
5jv1paygqyMOci4RAilbLHrmSaHJd11ZgKPdubrNW+jptyOJJazKmgr42I5j
vDuf7sXruuq+79p0bCCilgerw/F5l57JdKaoxmrT7CktuoQQdQA1jvOdNk1d
JJKC4+aWyfR2KQmlyQL++ZbcrddfrFwezt9yTe+Y75ApvbnrdvXS7+EQXahR
bweML1pwg1q0PBEiRa+Q0GcZOUzChyj9f/CnkI14Um+j+puj4Lb0q/P0k8zX
/IlFFThbqnSXlOiiwfWF/CIeAoce9uM9Yl5aC5B2RHAUP/L7OMW9LgRWsoT6
IN4Zb83qMm3bln0WbtsIqOIkDtBWqUtx9/7qUy3MjR7WOtJdhEQ/Gift2Npb
4KUy7gG1GkSy/MU7Rg4mWEkjx9QtqwkdphiI2h4pKb2eC4Pr7Ng8e4kAVi52
Oz4WCA/dgZLjsMvKMXKN8ZKnSDlcVnbvje/bXyzFr8eIiWpFqPByt/NbfYTI
sYBDCiTbumCCcgOVewiVAABRJ5nnxdHGlBriGdbAbmYjRo5KFUBZbEXkqh84
aIJ1DO4jeY6f69vMFZ6cJnnNhBqT6tX7cezIuexk64PxOLA/eYZaXmTLbepi
KAOmXZdy3xpJJgwCrIyqcS1pvWpcChkmYDeMy/00m+45LjV0h5KwMYKNOv4i
OMSRDg7w5riYMf7OoKp6aOjWlok4txoTVVLHoJ0MNdGxcDqCIdf7VYOcQN2r
B5KKgTbM89Z7YgnR6Ei9fodpM5SRhn9D2djkJSU1fDB2TCWu4c55R9RlVslE
ckW+Qd9ckWRYGeu/XcCfTeHGOXbrEZHQppuk1DUtRroatMjD/8/EQRQUKMzY
+fczktNUPvN678j66w4NrYxZEKC7Yzlmd7aBPumHlI3yyb/J+LSxT5jaEvoT
xKmSSjx/ky0KzNupKGiJKlGAWZid2FQAI92Oos1UpZM4p9xGyABreFBqo6rr
czjxcG6PSLCge9SzdNfpHFh0HnQR/mMCmY0JCEBtVikTt7BqBxgxQdDo5ZP4
8oQMQ9vZJZPSgx1JIiRj/soJ5Ahq7anN25zBTB+NGW6QHpWmPI6N/Fk4bFkh
7oU/0S2ha6mV8S1NSgHD8E595EG0hjO/0r4VJaAAHZ5s7qyEmXaM6iEPHM2+
iGlssd/m+VSp7R2GFSSrbBLLHs4qznSgivPF9Vb331sDo0kZfPzTUwJsiS5Q
QKPdIdnmKfvuQUCobrHxvNA/hK0GImgn6P9IvgyyvYiSWNmUxhqS50llriW8
KMSH7S+9dxeubazT2tqFfmmhpZ7fjQtcDQJTvYjGMifED3FKf74xSDJ0zNQi
amJqHtmUG0zy1x7Ei0FWUcsaN34ZHmI+khdLjGuv0vuQlduF4b99MS154Dd+
vPmPyfVgKIcgTkwCE/hE6WcniL1HaYrck/gLK1BtzNovGibIlWew4GwtzjmE
s60G7SzcrshpegqqpHJnXIP1CRFXNyMyghZBLBWNWBnrr6tDT/Tvr7IwHZza
zfTXqJzGtst9q6xve6XuSFQ/m2uDUqo8o6+wKpzZz4RXZgIKn1WPQLyaf9kO
FFtZ0iEqpA0mLts1ELGnRNtL0UTQ1YLZXk4PPUWOQvi82PxLDCcwu0A5wq2Y
dfJC1v0AQlZ+eGmcQke41mbuILap8rMYIPxINIJwWeP5t2Xydhc1Ct1BcYOK
Nk1qz9Vdp/4JJw+51TfjPcEPyCliDc1V5GipT7T99i657DcT3U2wetMNf5LJ
Nla1zJ/I1n15z2p1q8HJQIU5hf8/oxcOarxwdi8M1EsX7DwoWrw3TWYJleXN
rvh2DQ6imTH+GYZypuaHh1lFQuQRbj/u9H5V8IdT/3HHAFNBjsiKoIuWNBwW
BWuBFdYjpk9V51dY73myA/oa9UoahzgZ32yJSBuc5QfwtGAdw983hifC9Dz2
413IUEMNDwdSF8OWsKao2SgV3eOdc27HcugZW7ITwPYSgtFqL+ayJy6Q1gCH
CVmaWZoHH/xKAvaSE8RiWNFAkfOnJCI5t9KNFYjy+MzeOP011gq/5j9WuiBf
dU8m6+WWqJeh3NqavmckhUfyNpKitNhmLg2S00WZ16+584odDbyeo+iXzKNt
K2TVeE3rqPmNtCjAMU4wB8cf+GZL1N9XwJnIMErZU/N6WhvBOu6hG0yoVWZJ
J177lg4cZdUINh5LCH6pfA5Q4Q824yhvG1ix3PH8OeKYjyEwDhnZhkEVq7Qk
yz+jYWiAI93TEQvIE9TCSkzsPJQIfP67hrGu5WlE+ZTB+bpFRwUTjQMpLLGK
SeCUxMVZfCfpVXfX6pKP0Zl1moPBOhXgFkyaAVb3RylzURne7hmRjIArK8h9
wc7cGfKzoDWqcoZ4X1lO8Fj0EoDjcnTGPmGd1YJuekPk3DkAWSe8kUTvKZhG
6Snb/DsD6zTkK1ZUysy14rOXJz7gawZPN9vVvma9ixRnlIB7gEwAAqxKMZYa
jfT3QYPSVmUaIs8dv2lgaIc78B5w2Owg9dCYCjIJhZazxFRbQdaEmh1CTUFf
ZO9SycL0BbMgshlQNOxKgFoqM2/YG6DMwGH9LxdSXoSI6Ha3uok69N+p/PSk
qkkWU1uGXhCT9ERotjIUr71Tsz5mPhcC+KQLUFa1KjLJ6J9KdNmXf3Bk542L
9oont/KO3jMsWDiT6HjbsOOTA54nlylZCJ82THATxnv6QL138O09fr0JatEn
p6hNGOR5TRTV8l/ubMUuvjIQtrThcqOsH1YywVpoMr98s4bWzpzDVBlEpwRk
TW8bAsLp0odGgzhF61/nfxWrv8LJk4dtvWf4m+hYPnngAYJAOk7Rxlz+gO44
bPklJ8239uEZ+4iFG4IR9PY8hPt9OG78A9EMMpXbXlTwRiN6SMmeO9bd1dCP
iEawufRwJamDT6/eW8/Ocsn5Ce5UO1aaeZODSy5jMIYFkNuZ5gJwKkX2vLZ/
pWTEDniNnY0I8ncZWk+x1UWPZiDrACTdCGVl4ue+IH2ulIViQfZS3yCCwsU3
PPEbEjPczTF9IX2lb8loIzme041Lus/IMh8VgDCURvzwe+9WT/5l5WKIsYoO
J/VUveJPyS4+RS7/P1fuxkJFXMsnYwqUTfVLqxSz408cExG/DV9gU7JKKA8N
PqMcMbRdkaSgO87RLlV65aS/JZCJnRfEF4fb0swMuR6VfiDtIpybJ0i1wiUj
gTmq5eJWpQYrVPCjHQhAgNw61UfpB+iGOwcqfnWhlTRe/pTJ8alt5HYOfR2o
/bX7Uf3U/6fsWJ2nq+7olWEHl7vRmsSdu+yZsEuVGfigF1HZYQtJq9nD0ne1
+GPIweqr8YDpD3qrO4kZMnjO+9pg9/LrYxklzpvy6A3WDYKMvuYnVJhFvtqD
YbYWJWGkn61dN+RQFlkr6llEJumxcMDNG2AOpXwrxuxHm9ZZNAbWQg+IKa3S
NP3dUN9hC51YXdn8Ted537nS52PRKsAkzhZgvKA/lPRs0jolINEAaZ4RFu+m
DQQqefj1Evv4qiKfFY841m40J+DX/uT8igSLEdGjhqOuucnnVn9KJiPIUaDZ
h0n7RMfoN3MlULKhBSrLKu5b18VvthewKD7Z6p+t/ybS8gf5vgH8tEZjPEec
zt9tYnP8p1nVlqR0eLWz3pWTffZaAaW6xePyuXw4vIFIb7KFkN5/ILdfCmYG
6FulCYqmea7pzSfK8HSd3BSwdolz8AnnzoZE5EsjYQOrCJiZkCOBnkCNi2Wx
X3iYTbow3ERXuzqUYU7OaGP/oUh8lGS8i1nAhyaIG9buMmiI1bm+Mv+TpH01
Pd3e4RgJsDLNbVioeqUCXjS+sd9ptw95cmhli8sDAIMfnDT87RQfBK1Iw/Mh
dBp8HGzGMWW3tHDZPgGuM812PXTHZwgf6r07rDAnI1SGkauCRDtVV2LpHor8
aqxEpBaFZIfKac/FctdMXgaxeF3/4TFypNC2W82fkpgDa11AcZ7oo20+rJpr
sC7l41JHvdco84AcyO6ceKOqs996eebMRq90hO+noSLk5y6PM62gdV0HXLPp
gRX3sGOGrY3SMILvBkNiPrvaH7LnuNqzl9dowId/W7bozmHn3P3/WpPsfN6v
bAxlhBlRH/OzElVKNleRn7eU6jqJSs7iz6Cxscz97FMmZohnCPMUv7+Cvgxw
ioNmiq65skJwLBLp1TSOHZ3DCeFwUei+HmtWztkGd9ruZXUaDgvcGK6YueZ7
iEvlx/7WbtLfQHTrC10J+AGQLojlkEP/JJlnJbbQZ6WoxfYsU9d28c6UfLti
pZ/RIpS2NIC21KrlBB9TmVL6OFawDT9qrq7XIE37TQxtVgVJYEMFNyIISEhV
oeRvbfzJexNSpWwHbOxLK2LHrbwRqPDPxqasnIXSAj9eaTC4/r4V2NOSQSvk
cq1g4VMszHP5bjOJ/gFvMecoL6ZAqaWShi2uRkqeQI8q+oUf+NSzZy0l1bAn
8CZ5o4Oe0EgGHnhoRf++ofDLViqqAX6VSiBRf7x1x5DVA2VLDo3EqQOtBBOS
j1nv5HXT1hxiPCq1ixVQyR0UwquQjNR8h5vXGkrfvt0PeA5TczCzi+FFusgT
Nz5lsVW3ACzB+fqQR3SU4dDyhg6N9N4W7EXM3k0xu9lCnB2NDSekqv/nkMVK
wMQ7obGs2HE+B1HY7EQ8HDVNi7VFIp2G//wN2OGaiCKEu5Cz1AfEYwXgrT+z
JCorumilGES3DDlvXn/TFsn52wUrjsMs0etENw16NeDUIIPcaR7lxIaH7ycY
zLnjKoDfLnq0/pfpJ5pu8f9+1IbeBFRf21xSas+eh3YzzvPLB2ybpHf61WQg
5b1AnEZ90I62T8Y+cUsyGkGsBLisRBnoLX+SwwcCoEeJL5xA/FdlQ111W64U
suiNvjvQV3C28kO8hbSjYkYJLkMHZvRikxLe7IZST4/c+ma2WoPsVVcmHF7b
AwnoTBGf0YrZLaFwR7XOiGMdIs13ngX8phElCGs/jqj/4yveLCE1a6D3kqei
hANPea0rRYQWPUoXTKv0PKyKP14hjZ33s6IajbN84XWeWApyQPT4Ylo2I2g4
Q0NjIM/ZPsXyiYCsD8duhqXmeofpgX6pw3A3pJJ+lNGq86j5qC4B2MsA4Nbw
peM9FfvlU00a2gBHE1CmTN5oCe9cdFruAwt8t8W1XETj9y0OoGYpsAbWWQnz
VSxmaWmjki29PghyXYihMSfEEGEDIoRjWt0hUKox/qpzTGgDCmtN6pBaWL4v
7XvSLZhr4UtVFD7it7t8khyfdpNwaajBjVpFzmiIzuksFv17jxLa9AIfF45v
r07Zuz5jQ09ZJlThxZ4pPqwFsiudzTZedg24iLbH0Dz+h1T+eli9rzTN9TUH
BOgQA2VKTLST+pZKUfzfP7ptDejiWid48y2iweeHmiA/j46+THSBNzFjinwJ
F5EJw5uj6G4ycwD8QfpJVlOwiOTlId7iOccnEKJ8mtACOtGWqc0BexUYvaxB
DckQK5T7sUx6B5FlJ4UMlk6GVG72/9J3Qf4ljeTu+oHs/jtH0N37StXDfxBM
1dAUA7gdkNZlzUMS3LtLLbNVkj0Kv0+yKbAhbKNWWc9GMxRGWxP91hOEBBD4
qczi+JZVSIgzH5HuxeIKQxRlrqep3KbZMuM1WyzK7TkAbMYQMFQebIswZxwP
BF+Yinlx9FF1KiUQVf6qV0k59oUsxkDJyhEKfcj1sZQMVFwZpk7pt1aaz4o8
1hklSSShgsosrfPANilyfPBtEKPlRkj7sJHmggCMOmuEEankwlIzJXntO4vR
9IbY+EwY+NOo4srzBeMxUttRAkFtE7LkB/Fg6NvnUnZLypQCAqUGRJW5oi6R
s812a3Hqoi5vDQaWMbjjSMmq202QV233MzerNuHdHCnC7+zmvhwu+smKSLT+
evIJznzZRcJqJvZByi3ym3RoRv7nvaDAP6cit2BZOxkwfjpMLlg9zjv6UYxy
g6jNTAQpznATTO6rK1nyM20R1u0v/FQTnOsfH10cu/c9nMfDo199E46dQBYf
ASspckQRR0ngNsLxCI+Iiv3regVnB8YYs1PxJvFfAzTlBkEHxx6YnYLm7CB7
VWk2dnBMEiRxPqYloRLgFtUKYivHWi72utwco5PhUa4MI8g22YzheuR8hfCo
aeDNfu9O+3nESx5UhJIeEClsuL2B3S0Wf7Yf2EA3QjEp+0MkugVatwFD4wjH
tFgjHJ4lW4OiHiS3mq4wEB1QE3DQByoWbd3TmIUYyDGJfTAJIqmOQqkOsuCc
v0mdT6rtr+GGY6yBgYuVtoLCXG7izkfK7V3pj/RUQRc5ojEqqcqjNiMkstob
xXgf0YF8v43AAhsahqAriL2thd2t9nn8bZHYRYuEz3OzvP0L5BTbLtKWnX8W
gsy4CRp8WLeLuQsqLv+zaLZX4HeH8NDU+6B9fX0xa+IEerXiVBsVdB2ZxawJ
r5MsDSFjAG3chFYMtWUNd7SXZ1+UU3wezpOSIzQMdWPzZJWJU2Nl0dV+xp2m
VRS+cZBJjnBY905oNbBOD1uJAFs6HDQEdhhMqVBOruoqxo1VM2vfyO0OE5tC
Poyf/m91XKHqIoW/WMlgVssROLjLfYg6SkO1kBdQbNADfLzYceKW63NpjrMz
zY5QMzsShLek/imArrCbb0f8hpohZpSCSBX5idww7F+sIbFg8PIAnmv7eKNg
e57rKZ/4N2NzBYd0GOprfIeLL7E6nLMZR7wLz8gbxiBDJjSxc5Dk6/Ef/0tb
9gw7w1VlYfw0bv+3gJSs5nI/YZa0WiiTu2hCwz6fXUNJ58Eox5+PzpOrfzH5
+al4d0g2zmQtTr5zWZ5mg5cihMFX31PlFzuWFAnPxxKSKsdOIhtN0h3eSfGv
qm1nDGfa78bUbsD6fkVhqqxlp1JWsXb3ZDkAqW4dST+P371snLT07eoWFgsI
EIkgs3+YUjAxhKZzoUceADHUQIIAhnKOJ0RnS31VzCx0tZx10wjogBV6vFxK
NiEQxBZJxoZTfuTGyZVCx2odAsxbGBCJ9tDongGdi0RjaFaVsdInNBWGpndF
+lUKn4BA0tajL/k8Hb1R1yZsTKOO1J6uGIVC7qlh6CvGdGaVIW+lJdqzMW10
fjlDZg3mkvn/xVoWFx+0V0F1hdt7VOeDnHQ7mK50wymlXN9jZ1+fSlT+IC1V
Z9wXeD5bl/cK2FnIHhUWktMIDgtZc5NFXTumcXmmaLw0i56nAeXkZQvk9GLe
7SVf6zJQA8oPs7uE26CBjPzSTIKog/O5UdspLPwJviENO9tzRTYNr0mr1hRH
BqYhzMihac4Vrs3f+oCJC9/6YR7zDRhQ/8S130J2igiHcG0e4PHvQxAumJtp
r9CnldWhG0x30qcrMs7anpUiUJUaJVtxG/+gEeJZVdlRpVamU8kNJRtTvrMP
S/E2YOMouFUyzY/NK84IWXnQCT29AxHhIbeq2GSA5fplgUJxdd3MhJUXSsyk
JGzfVEEJGAPNQdRQgWtMywPbkAgJqwu/iY9JCo7jifSl7Knf3QJdhuqpKGf0
NLalo06nX4oHK7ehWWreyFHGhCHov9Z11SVDLRjpsl++s3TJ/tdTtax+ZWUj
/6QEgi/eXyM6cdc7VXrMHelbJMu6zlNv8+JprGMpD5p2IjCCZJY8WDLud66C
zD7iLz0UxJtF3Sqq8GdwLBgnvy3jUt9Gvu/S1a/5MMKUP3+4QShA6NdTx7ew
KYFBbY4YbVpzP8xStCdHxcXKsMZI26z2J52XKkUL9Ef0158tu1r8+X8qDxrJ
pXGElSU0E0nvrvLwxhpXnUEXudviKh81v84BfLoCy4OSADylWMxdHEyfiV+7
on//sjkNLXXyz6YNHWYsHbWti2r2xZeTZzwI8l4pAl1KPI7QhoQZnKm8WRMw
+Ik/TBqp7AX3x1GGt2qc02xWP/lrrefewHBNBT7F9ieh0HFk5PhcfCdm1fOl
xi1SXDTR0wGvLUCCIMktjrSU+7DdXtEwBMmVflg1f0eW3Lbq02nR6Qk8MGDC
XE9Z2DuY/lAKQfZzQoIUowEujGEqpWlznujBEu2U88OKSz940uyF/7tNolC1
KlFAM3l6PLWXwVd2EuRXyxMSvHrOBeLm+0YruQzQtFE1yZuyWyaInfE7DQ5F
GPZxKnTYtlwpsuAM0mJn1AtgP5O5ugtJ6hxtcnTuo8+c3Kcni1yqljvBEqFm
i24Bev8hpIRH04vJaj787PZvohomLjuvlkYO2cn8SHw6JsEn8YJCk4j4oKuu
NRvdE/zrA6B9Z/Vwt7DfdMfNXCorVy9xLnTciTGqBNnPxOVyR+uIeiuwuEwN
zkAOMUrwTuXrqAHVrXD2PLRuQ5WfokgBuliC0SjDjpfwBjcAaxLSkYI8ykd2
VQgh2gqdT3ruhh1PpyigrFUhcbnuSac+4/dAIu14SYQjMSqi0xX/PZWSpCMr
2uwwH4pr0VbXKsBjK8cTcTuoo2EVDrirAkzQPlNB/1yUAboHEHFcy76++UcY
HRLi15Pnmn0KS++395ukXmWgTr9/zi2q4u0f4g5RlhEPEekKcUDDpg3SwZ6F
m1o13F5OCzUFND5v6cGAJ0iGev87vfAWnPs/IuXPWfzjiF5u3707yameJp3i
IXPBBT8Xiev8MhaEnJ5W71/405XESsT5XdP4kJKX68T6wW2c1wsOqduam11n
VYjGZf3RLuCo/QyqeC/SoYr4ZjDFmC+5lYbaVj4TZrB62qTT5YvP/yYGIVLu
Yd/MiJ4dzs1yIJQQrex2cLwMZyJJwv4teDornLb+AqHYyr2VZvvj/rMXwu9f
642r1tNaHtqFnuRxsJBPtpBag7QYV3FDqzuz84xg1b672LrRKp2uVGv64rAU
nMuAPi6xKFN6qyF3jzInhM3zX8yVDEwnkuuvJGWlJccUFYl1myTllXtIBWPo
ijqO4DSyldUebFvlcxGzMSSifp/5CXOti1liNOtHd1slad6eElARsjPCrPPh
Dim7Xo98qWi/W4bfV22yfKBWRZO/jrd2/F2WiQsr8cEmxzx5ezgWkAOgiT32
KcogNTijMERdVD2dpbY5C1cyeVk0FzuVKT8qVeSPQAB7bOPAlZzC741ZJb/V
y1RFWiCYLMXmvC3ORZv3sfQD5i4IN+rgc7/7WUmfRTVWWfbg6mLGGpbh5aaI
KinfwKiaQcojCUW3bk34/x+nhHjlSF153Ik8Vkvwvp+bxV+W6iNlbXjXUGYu
ux/cePR/ZDVghUIfO3+20QwcDi0SZ2uBnOeJJR2zsf2x+Xmrd4gGfF9IjZFd
5KE68gmg7LGM/J+1FVUfMgV2eWJOlRXdZQ+2Yi6aejL9SxdmKym9bNnWxCa/
RdTqLweqRYobFQ+4SKDYXBTjGXzOcxh5c7yYOvDxPNA9YXZ3k1T6swZDlV4n
f5IrHdz0pR5G7tqgaihHgFERhoKx2caacy1XRe4IAG8y5VWnW3Sc2KSAe+99
ZREMXE3mOk3sxjH4EeH+sgpt4NZ+bjDDwsWyy5bNW6o+Tg9mEiMMNa3s4qIh
klc3BOD1E81jmb4Rx/jKklv8j34ncI0U8UL8/qixJe6NCNrA4LDB1WcrOWem
GCFJUZU9X4c+s6Oy/VU98mkLHTzhD9bbgp5EmPSig4h8fSsSngE3+dXOT0B6
s6iE2zw1YYTZJVQ6j5DEEXY6AFmZEUzgO4a2hQ8Wcwo5bDIara2vu+E98cBc
UsiDRU5Wj6TJPzFvUlQnBUJvG4hAaFUU1Ub3vLAU2yMEgATF59kCYfn40+Gt
WaNwg0wQOMI5QTyhjCuqcy1jpY326ydfdudnw7BdeNEwL2VtaPdkIzlhRuKd
Ot5VKiqa/SiD3Zr8KHZy1VMDgh7bOKi7xJWAaL6tR4V6VLgEo35BKyGVxR0r
hXLPleZNX2HgTRcBCQJClrrSCXHiqNKHq1KPRF9PdcyqaX5WppxT/fZ30R3J
DlofCT+NHeYyhxOM3eBZvgPKvaWtTsR5QFDJ5nvDJFOjn8yLrpQVQiCjeXib
Z4FyIDEx7BRoOFA1JTah88VCOLRtw2GIjlqHMfXSDNMgVfmdVZ6UqTBzJm9h
w6DAFsfpUEFUMEWDQJoPANLDWIYOeMnDwkJpYiEdoeLC5Y4kq5DL6tG0Q4bn
DtTXEU0JRHMkwTbteIB3KxWsSc+eGpYHTtIm7dcjiy/4LOQzH/rEmsyl984m
kw9F3itsIpnCqnHfI3EE6T3L8hOoWnEHNIe+6oCtuv4CjuBuxkQwFQhgOomc
4wVcO31nMQE5WemQwPCSCxYCamck9XVUkZS256SrTMDO4dhaMe26+W6OpOtf
r2I+aGhkFzqKSKQCCK0PveFrzqP4Iet5/MybpNf5IdzJBJUy/t3PGNqMGylk
hXWvenx5gGL2rN4/sGyDqVfoILxonsPG6jF+/9lzUHIrEdZJVgZt3okj7LbY
YGkhHQnrUMVeEnJyW73Hpv454ci7X5dliq9YaYz8ROv4PBH/FmtjijjAdGPu
/B9mmC1cAzk/R+RtAxftakblFKYfyb7Q9d1OvzrSl6EZkmh4cx04Ae5EFBnA
ZzN3rzns1APR04F4C/2yhcuY7trMK/DInmCJECeeI657DCVzhobFVnkaTRKV
mdSFCZLv9qu1JqZv7WUIU6eEgiCsE12oMF2ucDoDF4j1Lvc68G6rgamTF2J4
2KpltJL/ot5AU7+jCA9CyErxfMXA+5217z/t/+IZV3MSyIfMPZNE4QizsLQG
zrlNhSKcoEstGo7yCy2iIKOL8hMCBnN5pOumRSNJSl+2jY1iQ0UugHpnzA6V
NayuMiUizA5ZFuJVyxAz7oQ3o+GVb/FMMEkH8b7mbBco4AC2+Zj32x6FNRdT
VvLWhUOZxjnyBJ38vo8VEJiEp+3deP04SKeeNSa5BuD2yyxieLOembYSPgrK
qtL994KoAMD30M5rPMEfRnn4s8R2iGoxw2hV2mDbbuzgxZPBgEONA0DyAsyb
6asM8uoaPar2oaUuhLpM+OGADTkQX22VRTz+qEr/amvfpPlsBglPpmLlDcHr
jktQIMiQ9n0WOfXdp+6IoHfyi8pU8+4dzoDNG3O2Ca7/I4hakwBUft8T9wei
7ma2kpqTIwy3RnSaVjOgZWd7O89eIRz2/z7deyL3UfkDY2znxQmkXM7Lj446
IVqL4+UvufA+R4cZPwoNAn42Pn93KIOR7yTSFa4xBGC0FRQvwIfnYMGYm69l
Iak7tT4I7APt9FtTQ58AT6TlzkWCvloPPUDVd0lFnDjQkAlEXGYlh5Jm9Flg
ARqMLwsD0uOoMSBlv8dsu6kpj8RdYg4WJUuwEoUbDuHd9g9LFpYC6zpSqfxi
mSChDaQH5gkRZPYXdn0Ndp4ZvaTx+iHluSJ42qv/eocMuAyOWaUyEefp2ZD8
LYPmPwLMe2Ox+gsQ+p8XONqPP5kaHrbzDg7eQn5ekIjOY4G4ShRLNFFqiKYF
pH/DmjS6WBAZfS0AElBV5MuBJV41725960K9DWsEc5MQK0ysIF+ebJSKOr+u
VXuHhP6MUwrgnKHcMItVGVlYeV/CzR9Zti5TWxUzjAL0473e5cL2dr6d0d2P
NXcVg6/ECtPFWeVFyGx/Bx5bcJJMbAX3sCLyuW2WGbvVSbxzwhNvQh8VsEaC
1tjpTtuOtHAbA3qJ2J/0MaCtrIIc/Jm1+s9xsQxOLPvtBklfI+w5BNXZonXD
orzMWKS5zcBGA+dYFqlUtf4LbZlMWg636O242bjTrjJ7YiQrLpAFmTvStObw
Iu1JnnWC6Uo0muJmuOTh9LMyTq0WhdFu1neJKTmystdrM18Gvif0o4Jut61v
/cfx8vHyYcODg97Ogr6IiJd7BfrwTdBA0HIqzjoUBjTeqJJP7+v5YfrxtmoC
WjcEZ7d4wwS6XFGQ5pKcLsVUjuYBwRD8Ns0AApgwmXCrVudSN0fg3ufUzQz/
X24DSxHIFLMrc1mNv12FOuoqXSwPdFiaCQ3hrOxpyTpGazDqcpi93V9uubJ1
UwfzcdlQbrtoRjmVUrAlIq2qhKEzSrWVOtSmaP2cQmAZJeEbaNW/73xNHeP/
A4qCQhTu9Zxp6zVKhJBS8wTelOyZuDBotCUsdzDltvR2VUPYuW/UJhrQvm77
00F6QmEjqO6ChuD3Yru4asUuYM8pAvF1SQtFbWOYPyeY/lEayodceQE0gjM+
fQ64F3Of0vIl29tGtgcoUzhuA+soNmMOZeY8erflrsnA8ENssop6tJBHNomt
00sTq420sMuSoBRleeYFRgaaKT+aHIxNjzZpyN6/joNB/JWFQaouQSSF99Yl
J3EmPIkc5Gb3tvz+7OVwctCG4sxFxNbfJE/IBGI80kJQ0ErvkzRwnuTgvj/Y
GblSwFCGd+PD5ISnbEfSGUoDh12xapSoOMfTfbdUrKDkuYkCGQv+ZdZdATwz
LdD9VdMN0lEq65htVOrP0tUg/V7uGqv6vVqGTcb2JdrTGcUfyKXSv63C0TBL
TBJzftxOAdJpx9lQfyH5GBxMwY3hNASTB7E366y1FXeecUZF1G0nSUsbhsEg
c4P8j33eDtVzrPqhXy5QadcXzkXBIc2lG1bTVnyXxdG8kS2oB07dCl7M0FZf
Glb4oCfOpnlqQgwNJ3hukEER8X1BBoy+PIvRADO3yCI8/KbkZchsKZBns2JW
cNZ1x3S02Hs7/ZWZfCY032lvZCGjgfxrvMf1ne+7iy5FweKgDHuIRd+gLX5h
5w+nzFd0hj21Tb+oPTsxwlkzZArT6R18xkQGYRDHPILDcaIza1xtdWOfSGI6
aKwJKWk/04ewMgK3KOHYOGzm9YZmlP9/T/e8xXnFzWWmNN2LmfacEWdTyt/s
fPpxmzCqGiL3x177a2pHAzzvdGFwOSNPu+XrrkC7U8aoHs4OyvhtWhUxNyMP
rlGSMMfz53Im91W/kCCVg1T6LR6zW714iNtiwHzmyhLRIFWpMSADwlXLS/JF
zJ/ZCM9snFGLbuqv2FLCXqSGBLjCmxieNYxDQALMY6zyIeXMMb1ZBo0bKAHE
gDwessDo8Gil3KojJB03m+vncS1rIgbZ1yJOj5TfHQRpqQMjBX1gWRMNEL6+
IHCk7a32Y3cCXaXUdUyfyfqPkEKDJP9xZr2CkkILJfJV1ZKrFgP9WeawPBot
LKWdlQLusnsbnsZTRLjynA2H0xTelTo/OLKdmChXOCbPIe0VIFZRYbssC6vY
VZPyu46ETBK5MqCikFN9r056Ys81yDqCuw9Zg2zr2Ny2aXwrgQzRPbnwbW2z
74NHEqXt3o0vV0IjGJ/s+CNjZ8ZRVC6WgDJvJqwYdfbw8WGN8BxA6WQB7F5b
FSprcl9SMABvnyk9NLLZWtfu1kdA0HVeH8/tOQD9xGs03wLD77Xc+YzETHIW
V+0vm3toZjY551C5FCLWLdhWIP6D+NWZLWjDeco4uM1fZOzYIDmmVfXFQOSm
OosslIp99/sDd3keyBaZzVfXDB1i+CyTyX6OOZkyMBaiT9UCEAMsVJ0eRqTk
J5Rt/8buKjLkHIctrsrgoKnCHTEgVykd5gmNfforha/Sla4NldPDmos2wEHa
r7k9RyWGiCwLYfY1K2P5LK/WbtB349fJgayLFGGavyzJlymMqP1TdT+Wlyyf
nSoLuFRAiTe5xC7AFcrW2BwL9DyhB8Mc1wR+N2qXDV+5BMZYCtJ/m8ap/BJn
GGRcpLZ3O2w8xvSizFiGxAQM1MD8XGZ8yRX4l7DD30GeRtP6rUrnrA0AuTM3
SCNWrICD5C6kk9lpB+ALV3CcLWeVPZlk/YqQKB1ciGLJkNiIlSlhQoQk6IBA
UV/bXsbuvWF6UwzTV4PH/5MlyBAwH6CUio9GQeFdMD1lpzEDxxXuTp//DYbg
n8AivDYkVvg1iAFnoRfTAbL69H5GiBYYoAJGRLdju7hQeei9h+30Q3ln9DNL
nodXUWr08vSoVO1IdS+Ji1NoMW55hcnzpZSHTVzY1EAkUMLI/yxbgAY8pxui
RjF8Ukj7qdA3mH7GVRPW6Wssv7p4VjqBSltRqDgWvc9L2AbP7McPJnmxq921
btkF7iNCaGkbpWUuqkcPqqW7tiFMs5iqmrqTKJRVfDtHnMIH2Z0JBDvmskSh
39Gfz4MaVjyd4sS3P8/A8sDUvUfPqUzIqF9YxdlxP04bU4VMZO9oyiCI2RsL
dIp9ypgvlMQk86x9lsyqdwL8/OCYorh/M0VvMuf+UF6YVpscCLVjMqBbphwM
uOWkxa6lQIVdI0k8yxiZxSeEc7O77FiNkOHDQrn+TmANdN1d1unFssV+2cim
SdMp7rEo/iqjac/eN+yNZ1Tdfc2VUvD3Uw6XL/0C/J8AX1vfMtTJS/a2NzH4
Ke76cm4PoVzmxoDyH9SYqys7Axj4cXUgqFe9y48MoNr1gPM4+TOcLMI/G6B3
5uCaQbuT7VXa2KQlTbFIIItJRC76mHJJlFvTgGHTDNvC5c1lWcspZe6DoR7G
fCMd9e4jWMlp+nTac+EKL6LJ8hdtKJftTYnDRE3mkoTgaKQxirjxllLD2k54
NJJbCdACqoGqxIlcGYxzUGB9Hd2+JsuCi1daQRwPVZMa2q9OnZTS+PN2qNRE
Mm0VKQxnDznmDrnhY9caQDyq6K+zHMhFhYbap4Lv+nY610HyE7OUvoISIGrp
HdcmEIEBTi+ZkJ4USCC+d5ZNT4x5rF9S/wo64mtDGAMm9+02NupQ4+GrelWR
7nVlnNrvsjMUO+i/YvDQVBUbLGDTY/4yvFDIoZBjrwP/sYD9cyv3b2ZzC9Zv
SKBcokQM3oDI2xbCywAREgVDpqmLXJMiMk/1XC7fcVDlLGmXLpneTkAT89Ez
h+QOgqifi0KJkrwDJkTLFoMYw3QnqpiMSfzD26OQG6DGT/89pvwfhEbcEu7R
7unN+XEX07CkKcCtEF01EOt00Rdl70rLxLJoU6Q2X9FN9Og6VjhiCaL5DoAH
4fQWZBhHVw/7pLGBoLiq3OlHwKbLz0VDze2hvcrHJqAjOEtmsr0sQlW5dJYa
mc7B8mPmbMpybLdtHZY40I7RK0vfxpTNXla6A5YJjIj95Am6xRzhIou4dQvu
+9YhTDA3ZPeAxrarZet3dpVYdNVi9EEcM/dguoq/x5wjocSeUrTBVUC74g6d
skzPyQKDJacOi7pthWFM5H71MhRVVKsuuypUTTFST0TAUCt2RA7ZonDVB4Eo
r34ZP1MrVz93sYWWHS8CGq6DHeonxqs0Sx/nyhHugXhaRxXA8ZcK4KSqtNIH
WJ/0pY6/vlS4awdlt/Fda5ZHlThgjPxqkRVUFw7UhKbkyyO6UXMqgKn6TPyR
vOrVHdiM8s+KewWclYI5YVv/PXiz721xTdVEDASS5i7lmBVbSt+d4WIu2L/N
P5B8U/vxHamG0vTKGboO0gvEddQ33SKdRz60gr+GOxqBFAh3tjv5sW62kQed
OBCOyYK5Jh/zUA75KVVAflCCY0kEILdb1CM8aoy51FtRFL0FuQ3F4OO9mnyc
4LirIxQzi9fqq0RQOyrOh6z4+y3fJaSwr+AOy53JJ+vvTFcZPZt6YXUAbNT6
v0QtvAIsWJO01Iy/aWnwEzc9Q0xSgwvK7PPNC/znkqagpngxlt434q8W71G0
y2PEXFrmKUsjCWhMVvoaWTnYaFlsi7YPGAO3TflnMGcZgiwq2AkjeBEGJNvr
IWyRStV4pSllotD+mSD0ui085NbZ+DUmpXaBE5eXpmTGCvbCD5pvD0dn18Uu
RNCC9Lkc+PCoVc78o36CSrzXG4JDAVWy5kpUQleLmJMbac8mRbENJBllD3pK
C/4IaAgEpG/xypkkeg9f30GLHktjQxfxANt168nfalPmyhrq0ZIR4UHvEBOM
6LGYJyypr6ic54cl8m3U1MlcY3/xW8weLS4F6MXRnwYzF1ABqyki6OEtHtFt
Dl/FVlRWCZA4ncG2oh58oOfxlN1ss+Bgn5vqwfkFUWxdwUqeK/lFyeYqEPoV
yBeGA+8jIGqglMV9WXJ+IpaLfo/QdKdE3ATcsCX4IsI0Oq/bChCRSQzhOSXa
ozSHH8+udE5YlkqOJcFB2GIG+knCkMcuMntYUknfF3VUsjoQYoehCMCWrNl9
/42xuDljal28Baeb0O9K0D3I1aRHYOCkOcxUyoDAQET+iyVD8l3XyI/0pbTW
c/Z5hzQ2viubHLZj7+j8CwrZyGT2sTi7WEv0B31J1b7cN6z6MuXdkmstr+ZC
BvN78nQ8I8LVrZXG3PzCMcKxnEM3xr/F0YMowW2wC+D0hKluV7u9P712HLpR
aMUMsNKlvFe3/jE3OC71MWAsyYRKCF8yvIMqxzo64z0BvufojRpbWdbUn6IB
nzV1Ihi0kzjHOWlULoeXgO8SCKzLIxOjZQRiQj4nTj6fjZeFNB507p0wivtJ
N7wYfNhPfegKe5XVX0yq9n7NY8eI88IUU/BRBv3pEhBuCct221a/Scy+6sxq
jgk5lvDj5vAkEEW5pSCDiLr1w0TQKa7jQH9ldo5usyXgMEPQR6Q6WjwP8REC
dlKVJ89muQ6ItWZ6oO5eIXOaOcoC/gmlZa4dpi6FlKMrpwob2ZWbMUufAhCB
mSK2QvwkqO+k8Ut3LSv87qjpqGmftk/iO12pmiqDdCIop9Wbj9c9SsnRluXk
3x+cq8ZH+FxpQpfV3UM02tlJEwdp3ivOwUikY7aqGL4jGEb2ov41hWFQ7D07
UVNcgjJXhWZMsLqfhpn8ESOc1VL2Ns4BZBTo+LjLh6Fq0ekBFJOaXnwFqPwg
DfgQcdoF3pbx3wLh2AYo9K5yZKl54mve+9GeodXjTExYH6FDXh4/5NELVDDw
jVHcQVYeLY4EkVG4XqDJfCcYKvbDjmiXbZ5FRZrSmTOa4ttuv9CGL/oPVRkV
8IdYGz3HVBEgaKNqg9OZFaY6g/cKa0KMmmMJYuxTFsEgbp41L6P7v51NLO7E
FRa/vozcY6EEwvbydM4H4LfMzK1UVltXeVFEP1zRRXPjQykU4BB/FoPORmJz
2+ios4cypOrnncI6u+OJXtjqR01eRZ60XQJbTy7dZOdaz1J1jsT1FcmFVPYA
II2vZurPad4c0sfdbLaUpAOlVP0b1evCj8IQYSPa3RrkfCg9Aj4PUtzQ1H07
rpyW4G1tbLoH9HGzr6JQZhUTnsoFH+6amp5SHuxen4MuCnUxU9jCXbhepgr/
Qg/9UKRhRBfk8xiip5CmmKIAUQ29vmsDMGk6bUoUnJe/1WfG/2yOSKF8ZwEJ
UDb1gjwZafZnmYM1dwLWsfsMoUK5CPoDQFi/yPh2nqGFAS/dS3vmLc+IOvUQ
RRV8Vpkez/+iwFc4nmFKc7DGVOXdnU8XL+PttrhQWyCaegu53PbdOZ3X5N3e
2/vG+JKXSV1sqo4vNwd8hVtduZNmHlv6Q+xWrJigneBp7P313ycE3f6S01/S
4UoIkJw6US6FL7aLPbB6mhjRuPBFGTPRB2R3yoejEd0oR7oQxeUQ0FxCttdG
nc/nR0aDZUdNin5nrVx/v/fCsxDcjY6Hq/WEQbPJx8W3ZIuCxUUUwgzxHzLh
XoASxkfXw+4vZZQF4LuZ96cR2sM4PH4zN5WP9afWKodEtlMS6BtV8IBCRgQK
G0KqbmLYqz+pZSNvuPNzquHRwNZ+cMFSR/DCSAqFus5AjrJYpRmLDEtLrexZ
0Gs0tB6dK6SyWBQnafdok2eo5JOrJnyq2res3BYShY9PhQk3xOw78q68ylpM
3eReFWME/oscJUyg93mpSSIII+jke0PuzVssc+YedkYQrcgt0WA+I31BIZXZ
OWNjm6tnPH41i63h+NFjGHGYjx9P8MjqmS5VzkN4W4t6ezQ8YytLWvWbgFbo
5AVd9DMAsLQNfZPHYp8p2054J2f9VV7d2UvWU173kzJyXoygvl1BH+U4jaH7
t82ZK1nk0PIlJbyE9JGA7yJkedlsC4s/cDhnMYNpDZPHLoTJYM4t+1rO0WWI
9EgGKkY+5g5s9znnV8r+M6CfnE6/aUn5xeu4Kf/TU+p3z2W5JqbOTohmavLb
5gSWz3saNtp0tnWwAaYELBDx1syach2+CvySpQF9wkjjWEvNVwn0HpKI9u+l
BKYiRfRvEovW3ZZjGt7atOyAGTQ5IshaI8CpAzNsM+fXRUgMWFdmkI3Vabrc
cLt5FSbtll4KKa2UX5i0Ji+TKn/kzRf7M4oqU8MKvlcey+uHy2n3AD0FK9u8
s56Y1DT/T2gclOIRh5kaE1Dh/3OxrnX5xmKCXSQM1H3Y8U7i0hkalzjJk4sw
T7ZbtAj4DybZ/F+v37OJRTw+sRtpaoiCG10dXFrvgLkFUre0hLWSyjFrpJQb
/xlN3JhvPOxrD8gjduziRPJOaVTW6Htxeu5SsDkVcPM4WNOTq1w/pFLl6XhK
HjZxK6OHZ74WITZEK5q+nXTc2W6npvkMTWIEMSyd5inOnhRfU9vV0nSRlO5V
y0J91C9qk2/G4GIUrbIyNiDxnh1IMK/4l+q07ldAUFZBSnUwtPcIE/8/EJLs
CQ8rqauQFioA8XcJrLPl8JY7gPqOTYeAenjs/PFog6WBy1eaaHqqX0V0bkZJ
8TLD67zyQ5HTS6JIQTiTQBE1i93Hns53RB4j+BZA28tYhluQ9VWqC+VDWZTO
7Rbtrldi8UltFUgUBXKa+o0+efvv25aL89C7TyNogB6f8um/nrTSZ5PotGn5
CNPLNMc9CcD4OJLwT9YkSQSGFvXfYLU217Xjz4o7CSStJ4173Ki35wPWADDg
gwuXK5IOQRqWU9qSf1PVLY61g+EV5R1g+9KLhwNv3HYuuMhEqOOpwFcxZ2p7
VQ26VfZoYJd/W2IS8blWMsLesDqNjq1suFfwigMsV+Y5lzFeZvKOOo0Usyn/
Xaw95JPzSBGV8kRGgr9nDFfNle9y2ssBYDtjzLubdiJOq45alOEZW4vpJx+U
3M7H5JSINpP1Egbe27evo5Tqh0n9mQDOzHHsmBYJyYT4C+eT7kkQ0laQHvKz
6bI5fXClP/uTDbTwC2xmM7zYmrR7Ik4imOV8GpqYUkOYhr6LYDvu+083go2a
HIMTUGw7Iw07glJEjYJZBrjDalnB40ou2ja7/+TkUfhiYXnLuvi2Jbap/a48
MbZy5YUd8xwkt1WqJXqbKfKMOJPdvi7cdieTFJEDRN1Lk4D0QA0BpfJac22f
fxQMH/4U79J1Jm3fIB51VzGXKpu3ioBp3GwAc0a4VQL2bIOhEqNE8CWD+KWN
Kcfj0/PQS1ME+Zg4KcdycrL9kI/0AvFAx1UtzWBAZFUolchZVrb74wqA5TK1
L1Aq5Rw7Mezj2c77oFG2mQBRgzK217pyqSB8Mn5ik/Snl4rn+da9XUJTY9ta
lEZ+Jg+UiLK7Oj0keFdllI8o78hGNZSRciAGIq8BSP1mS4rD75FUCIsugTu7
Nnky/e3eJBunhvl8Gk/OAzJRiAuxdypkHYeic4leW0taxPocH4LSMyIwQGZ8
m3soZuDeU88J8DqESmCWezjqWBJYDQ51t4TFvk4Ls6ulqLbAHuZp1dCpdIkq
9z16GmWf9h3+qrWd/Q862SNKwvS/Q6gsoi4rBi+hEJNrFACzuaeSBVJJ0i7L
0yLpbrYdS2+cOk/C9kdXRyAkPclMUoYauWgezX9eC/uDVYg3PlFeULIifYDL
bNa3fElrPHfvWtJj5+sPqLT2sV4ahKEzo0zj81HmlRsAQHN6AcbKKAzMBZkZ
vq1TGMo4tnI/YR8Qxrek7l2UYTzmPhsQ/GU1ltCjsZUafV1ufrWmHBUsGox2
2jplzox3TWBK3N4A9jDCcKZSslGORmb4Hn4n7rOhEthCJC9kfaAvg8fw4PbO
Sxu6+/YkngYJPTNDmsf0iuX8Yg8ffdd32lgfaw3lZG+iwYPvEftnK1VcWq5w
+DuuRIGnnKcRA9ixuwZ6Nmq6COq5xzcrF3UsKI/02050YnZMD9HWkt+FUxev
ThgjkAPBnzmqKnQehMvNnITDDqPWkkpSCdAWjQylK7Dh7Jt34cpnlfDNKxYa
TLadqkyvXxFzBtF+PFqVMsSsVOqVFBCgCr0bZNTcNxBgGoZccL5YYzy7f/c3
DScBUgzICTlAQcbsCvDSSz83RhsOoySqb57XO4Uz4rs6Gu0yCFaYLLfDGfLv
udWKl2zG/EqNLmVQCIMzvSAQyNm7K4vVagtk2Wk6aovihzd1z6GcOYV0aQs+
rG2lpTTY8n/9m8HlPbFqJRHHNmWojxJbuOxfHG0ibkgwC0bM+N9IO0wyQrlJ
kSN5r7KnE+pICRcgahn20+r6aGBtzXkD9kP4xISyYbANl+tu5jCcAwGTasI2
P2jhMBi5fNVvlvbiM86uy+vJcOBRTbl3WLQwugdsG+TKJQd9Qf+k8HQbBf1F
agumGHYEZz4fRxv/4QyaDghnqXF4fD8kZsjxn1MBQiHqmP8sjNZOD7NA4dWE
mJsk+yt/fj48UQVKUnvzcLETnFvjpUWgp1KaXQw6aSK1r+tpD6mBPGBhNped
rLyyCNv7KcxaS4mVD1VsyxXSXcfoKUxrF0/4ilxNxwuox0mIMCuyY/3AgqQ5
uDKpegGUoVtdTk5wTQq9XMoYBcOgPDI77SVg2seBgPZ2wZ6jTIZHJNN9k3B3
GSjHF85oE/MCv81/4eXLVOqywFWfFifm1bSOOtgqD1irqT3KuCXfyZU00/e/
qE1noL1UCobA4LeA0Bn3IA+fMJFTVIVYT3v8/Q55WYVuDMgp+Q4/VXkc5IU4
JNRPHN59MwOqOYlDCV6kd8hqDLYFkvsO7TZzzynMbSaJMUCQI7ju/xIH7vQT
eLR7YVa8qqnBrA30NaCSFhlGZ4YlwCHr3ovL3hpYLvixx2Iu6FmI67plz/11
w4b+kbkeQPMs4hCdTzpDWA0LiyWLjMc6AVTJQA/UWRJttv3VDZ2JQAfaMOuF
Q+zLcs7NvXb07kjYUj/Ir/983WSKe9uxTArBLS2zcSUXIemuSCdovG64YIyo
jKPJX7hfQ3LnjedESlen3h+vKoJr3TOJYhkyACYOO8/t8sBrm7ewNPjxr1L3
XF4Hi0dz6X2nYYXT1L2TUNZC60kCUgcEC0bFY7pK2bD/wXnIvrwQx4OtyPbm
FFH1tD0AHpylzoKWJDhjnI174OPWh0YVCZXZfIvUZ4At7IuC35RTKXmWuUZK
iTwHAK4U49bAjdw3AiXSofkDzrBq6Gb8zK7sRtfSxymIilNyWq+5cYvH4oOc
qqnYADYbxW82IhJFKUy5GticMYHbw1O1eyfiFjw0sXbQEh7M50zON9rFtVDL
PAaDlEvRFbWBOB8XzBLhJaPzdAnKiUk20A04Tav7ZeAZnvcJWy7KEJTmd6KJ
06RVP9aLKDnoIXkcFaJat3mqONbutvg/iIJQtklwmN8LlcA8jhehxbNi7NiM
YJhC5P2HdVqAncclyfzLLexC37ByMIEj+WXb6qvthbNUZkSEjuc6avkW8V9r
SVQVrvvqntu6UUHHFmLE/BCr7UG7paC3BxHacGTGpGziTDrMWWdmimcCQfO3
zKk2TMyYFC8UM+UJIQO2HKRcA2q7P9Md1ZymnHge4h/74/FlHmt/eu8Q/Tq6
m4JV1GEdBD3lizhhRqFvTf60PKhwIrnsFHjs4mG5O8WLReDX1JLK59MriED9
k6vUOo5djaKsuRyQyIwmVDo5Q2M4t8gVGGDoe4/BGlmh9wvGne20wBu4YuH+
OO+RD3SSaKTv5JbAAFHjB2E+E+hfhniuaA7Vpsls6jcpc9YHeKfG8nP18NqZ
zz30/cZukwV+Z6g4ZoxDUC72fIPbnUWSj/srVti9/VAolq9sIxuQvgWqYVbb
hAOjU14WK8jNziJrauAAd+1rEPKnZ6j5LY/lnieAC4IF9UqZgbjQ4nQfEdyQ
Mqx1inEW5sq7+mradhbEqE2CljTOTcFFoLWwirSZR+qxEiOYn5aJrWtEXOV0
lAKWtBvz0dXUfdlHZeFfpd4NvfqnViJuDE3CMqmP22KA5ZR6GMrtepZa4du9
a9/a7po9b8eO7cLaIrBpz8+ccfuFC9P09P1Fb8rSelLbkWzoL7AGF/twe8Nh
1O0tX5bOF+6LGDLBW9Tujuj7BjU+eCRvaqj04cJ7VBLkRjvAETd6feQYPtkP
X5h9Sx3Z2GM17QxMjevUWrlT4UwlgnG9VNN/pL9CvnFv227TBD8WwqA57aPQ
lTscxNWDziTinfOZyu2kA7J4fDjmHruGiz4S0fUzGi+Qcrtag1VSSYihgUo0
Hxk7+N3MNXxggBh+Old2yhBcl3iXiHJhjbhOG4YkB9SLofuNtpl6lCaoJyfw
7wZRxjj30KeJGdDxBrYMI7DRfEI/ZcTFBDeeK+INfAJWzZHnKRM9eqa5XnkZ
TiqcJ7V7TpEdSxfn0rFZAZDlorTrYr6KEw6qbkS6dEmM00I3mx5QK81McnsK
oMvjm6bS+PuM61Tu8sFGY9AFZ/iJWZsqFxaYTXBeR5Rn77lXCQmhrqMVgNa3
i1j0Sw/tDDj5bA8kjSh3m7/vlpfQo8SIHIkjMeCJUzvAvf4drPZfo+LOLpWC
+TRphv2TB2uZy6/gW2L1cL2WLfAY7uIk8rlysb5HnBbwJj/y6iyif3JivofW
VmdyreFF3HeAPgL2OT9cjpHYmivNELC2J6Clb9ZbO3K/cnFR2+qUq5Y3bwD1
hKudpdyfCeG1YAkjRYttgO667wr9iii9K2OmrRglq3VmeMvFIT6sVzolCjN1
PI/xWqw+Ux+GojlbQusVFBe3kt7e152vaCkPCmhRmHFwfiiOvEbTrXKG5OJ+
iLZ0B3YssOeUFFBJVZRiKX4Y3SawDDWeolEAV60A+LKzdAz7vhpWOeXVfOpc
+72Btv+IwDHV3oRh7T85hJ3Ngayirx/nOp78hlGJE9P7cGuD8AVS2SxqTZ8s
40jdXF0JyH03Jh7kAM+9cO3ljKy0xY5QrtUY78yQc2c44ZmxOLmYJxs/qVot
L+CYi7N8PaebJAWD08HnlQHNw8WOIK3iOtREbBbXXmgGh+RhmGvTwZUSVjFo
D9a+aUF0zu6emoYjRCdaqDy50MgvGrRjNmCUKWVMEsaYnghQ4aMFMceTXqVH
eJfMOYwQ6E9wq4VCXzEDMHVPJ91jufpni9Y5WYwLO6ZtOy75xEfAiH5zex0I
Vsgz2L+gM26WICVQ/vzsO76euS5X+LyR4060/W9/3j9Um2N9gXQy7afTnT4/
dUiMfLblUzt2Ow4PsTM93vx6TkuEDeU5aX6L/KVmcB/qmpbsZ6BdTDw3Evu/
A2j9bzSFcULPhMP+RotCUuNi7VineLecLcwK5ipmAkxuQ3K+3ORKH+yw2TBe
RkQrIG2iM6IxD24Ko6kDWUZP7K7QxP6Fb+omw886y7llvUraDf8dycNbPJrW
ZW9HKsc5GzI0h99fbtE1vE7BbO4jqNHRsneAUG7a0WReg2SHpC/FGsRge8vE
ybz9U0lxTxPpWrjCfrhzVGq+fe1WHyFEybikm448FXzFJD0te36IhadRzTjK
k8RpeGASw15Xyrk91NqgSxvIjMgI6BJBNQ5i08vGA+Ie8qQHCja1bUkDYKVh
aBDv3ovyrfPjkE5fUaHpv7Bn2it7wBbYJdKjpzgcr7KwtV98SiYPfHMaYlJU
IzZPMIbROcdKDAVQ0OMdG9PTta4v4ki90Yy5X3fNir4PKNF7U+0UOL6/wjrA
9A6CdfnsXYzIS/X8aOgBqJGWtjlcCiFNloHKKed61aWfaZOnvOAOUaLwmzg7
4lgomp6vQPTjtjUb76Y40MdRbA==

`pragma protect end_protected
