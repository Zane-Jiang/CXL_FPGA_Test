// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
cXhmmNLdhItLUIIaXB4zY/PNgQc6CiZAt7fNJkPAv254oaPyJidRl+D6jCTrTOH3OzlyXl+pBelo
maMy4r1s9hE0+AtT6nr82lq+MN6Ak9eaLOj2tlW6v80F/vj4KJxjMBLZakECMTVVNQ595B6Oegt/
sDc5Z1yfa1N+DwLTMQ3k+HHp13gfw8c1Ckk+zW2Gt6x2d5vPRydKrxSiAq6owozEjfgkBqvT6+6v
WY/VqAWEbgXgr0h82c5wwUjewf/jGBcPAlkO/9k09nfiKvHYSyznrh+dsqtPcE8lk5rvkFPa3K0E
3Dj/Cmpg8G/wR3HBXZrkCvX4rngzLN8OR08IFA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 28640)
98O8l3MB0niUmp5tgzdTHw+HDohb0vtC3fyWfsR17AjA6xjzEJgr5kz+vWYjDP537IM7t9WkjpDF
KPdBQPxxdnUN7TEkwp0ReQXI319jAFeQMmZAWb2p+DNaH3ANQVt/U9NxmDDz7issTtcvk43dZcrg
LnA983+Wns3xddobqaS9YcCQhR1JDVIN+Mys8hURuO4yOaUM0FPN0UUcFfppe07eOsJH8kD4Ky3l
fJXR40ZXePQbCw1rLBrExGW1eg2PZddQ5oGWLhs8V0SYeFieSK/K+kqzPkzWHu9MTbKWsPYs4cjg
Neem8OC8Ve1L7w1YnXI4bHLbkMHk6QcHLvYbEv3mCNUEVpf1FpxSt80P80nm1d0Qfg4In43t1I+n
gUMjfWCC9ioxnNJH/a7Gu14Pxqwc2PYLmVduNvWCTU/OkrNadozk9H0zXpu37nYYHcg0Zk6gg46f
GIc1DQHfoo0CCuXAdFPC3mWrEIMPEmdIR1QM3W4emOJIEFCTBWgt2r+0ss51w3rFHpamfeP5o3NB
fPeBdd+yCdcQ9aZ+CUNXXsGoYDaXrtuQycMVlabg6khsiZfiOJS3tgORxkcxZLAKjgqigX+JuoFB
VKertOtaELYDKugWpXQm+97BkpKbcOvkvGMle+XnVN62mqqNT0QJx6WxgBaZ3V6PmHcXuyGhD+EK
qVvOb5PfCKMiw9OZQJRba60o469uKAE5spO7Wf1ekImHEk2JDMvAOT4FXLw9gFf3/mlIeOJoJ1FG
wu81cx5Gug7R+roGDYJjbFaB16CJprwaijDe02BaKRopqAbVvCSI6OhivpzBntfsNJtAVRhCkbzg
OYliHWGe7NSRPEJ/HWsvEWibJnI1owzbVDqnlZVchocePWGxM5yyYhAOXz/n+hP3wiWgXep4BJKK
bG1R5IAvPvvhxQXMv76M9ZiuEFabgMdHbkJyaiNRKpQLZ7x+xt45AfNWMluKrPJ53lFIkPsZY+mt
5jDFKJRCzZqkez5QHLlLYkboZp5fGRqbWmiDGSj3EQzNBNkwS0G8aX4UzhceVofElkW6YS1l/1CX
CiMQomFASAEscBI6emUpApTlUy9zWfxupMbtZNB8HbKQDXypWUSJORVopnF//nRrE1piUEoIABNM
siLz7StJA8dS9EtWRaXzNrQEMB9Wk0LZYK4NL/mkQ29t6Vf+iTMWvG4aYafDItoDL7oWRfcK0VKs
mMnU9Qr/HUif/Ybdl3NCgcS9oMe2vC5e2KYTXpaAFZPB//jwnVahBZeN+kf/WZL280oWzHaELnva
rlqP0aLchod6Pb1FFz80ZLDbI3ic7ozr1nirOuBlWTKJp+SiuSKfyEmt2Pnhe61k3j9KudLjgTd2
ArjFiAdg3dePaiOHn+9aDt7fTOtBOuvyC6eiUJilg8LuoEgkq4WYNcsRX1YW028zGF0+61DrnnJw
WK3YewIZsj1mvMyyGU1sr4kxpRS8KM4KncZopjBRhx5rIPESkvR0Z/r49+pS6DPOMzESjl0tw9SA
KHypnTsPHOrBgFX0s79Wfo56AVQzgcN65QQi5hs6QIzbkFZ/IRUDnavaMhAvajFNOgJ+XjEOSu+Q
GowGiB7GCIMZmUuIhybN0cPoTJz7zhX6gDPqOkJY/IMun+syBB6EUOndlIxvdOkitEuAVRvnQ4Rh
2o6UGwOp/q0lxSfqQcGGJy/AYPSltI4QIqreCxGD0wM1eG/zBrgLd/6qXNAYT4M7W8nExb5LG+GZ
g3rnyzeFphpoqjltdd3+WZ4QVXx8ASbsO8yo0nuOEbj3vcsole5jQnI+r+NzdocnBwADa3nKxSfp
06xmsdJ14QwTTcD39Yc1g+H1E5+Rix0gbvrgoyC1zA3/Nw6FdrX2xiCixhjWDE5oNXSCS5dkPc6w
QQM33JEyygt/1wLGyBkS+4+JGvKBp8wWaE1MR9kHJQZMDoHM6yBbIRpLGPCRv3ZzKT32CSP5NDOD
BwvwU8etquL/nt0yL6BDItPeDwqZgVK4J1RgKiENDyFGT3bOoGPpDnsllPZi2IRU5tamO4AjC0yu
F//ES4VfeQHyl2kSbxzeFkNVuf5ModuurIVNyhLdnvoOtYtlFORtb+HJ1XRuZjNbxP2VmZlahGXL
z0L2+MChmU0nRAFtjf6hGL1YUt9yE7iAhD4xJafd93cwdd98NuAtkXjUXG1zeJGRYm+3+fr4Laul
eELhCNYO9wrvhhMtJeVoBhoQpUzanOLRbVV3LyryQtKfxzHn5xrkXyXA20O3mXnZWH22ZTqbLtwX
a/uJDukvNDbRYFtUZQPUs1mwroMWeOHW3m9H4vpEnYuw3e8Udc7/7QNGn9GamdGPlJUqNe9HQOnU
P1Ur35vCiV5KoysnFGaHoIDjE8frQGSqzVNj3WTRFHu8rPG8N39ooz1TNO5DJXNPfBEk6i20p2k4
i43HS6OglU5D7S8mvVm1afHmKUFe1kSSdnjl9RN7Oqizp0w844/4SYTuxOR+Nk9fPpsZE3y7ds1t
5HShve03T72Pq8hS30n4JClNSrKLfkG6Xg+9gWQz247JTaGp44O0YxpJOeSEBz1BuqgHNNWyhZ5/
ir4zWYnzqzoHrYgIP8iW29y+kAtPnvlKBUwDUdFhcS9YU2PgvDKPibsZcCo1uCSRaVEM0BnBHhir
fGtD1Yq17KGAfI8SK7eJGsghmr5xaLmyymB/L8X7Tk+sIBbGPaAwBGG9q1dOKGxu3ZVl9sGW6jvJ
a6YnbrIcJKSSVBubDn7SIhlRIiPIJuyxHrIYI9Fs6DhI17IDVvdQYxMy0jCMx9kbN/5KUDbS59M4
ZQ1LQcQlAWYPKUKFvsBnEfDFqTlQzdnogZ3pLEJeuvQnV9eBWslZkpC8R4O2kteBWYwrMokuDmE/
zyT6yD/sAK+n6/YIe+H9cQcX63UGSOeB6A72IFsD5cbd8AlRt/klS0zIT9dhcNSdPz5+p1TcIxzt
ANTCBSPPNuHs2wNFN+tnExWrt8/p1rxyAh26Ha65LgwlESkm0qyPHUaDVdu5t9sj7HOFu/TdrYuB
Wpc51ZC2XVhEVdRzW75ISKUU83ERwenE3z5uFXao8ZIzDI+iwmIQu9nw9Nz1X0urTdZLREk6R/Z2
i8KmgaS6u5wjQL6BO2DH+ipE7UHAdp2W4Bq4tIeThzAqTsasZS16DkWzb5tXv1io4DYoXSKDdiR0
mTwSFPEMkZGWQPQ/7jurl5iENOdMY1xgDWdu3CCfXdXKtv3tJRpYR/gTQEd083BX6uHrxCNb46av
4RW7oNjo9ap+Yrmsu6L6VejG/3zZrOOCDUZHbIJhhxwi25++aNF2V29ljuyC1pQZ8PS5DDibxKGc
mBceCVbmyT3eGkr+IC4ga/WIKtKkAGSTGBfryneh/2OQ/L3MZ+CsQS53Z8Kr+VdvKVBE+2mZoobB
Wsp9IR46ll6NpqnajXbWQDbeBnBM4cOwYyXt667X6MsqKa+d3ZqskjxgCRL9uoz+vzKIjsdL0+R8
3dgLZznYCb9Fq2nbNsiZVfBnsziJ9qQ93XYQncW3ViJXsRMXKMX/NUyLtWa0Uu63WTnO4Nu7lxW9
BE37jBw2/nB7Z0SETpgcso4zz6ltMCS1a8r5dXmmouSDDovJEVpDg0+PTFSkKMorxAJzFttrNfUW
Gm7S9/Y49s+S3hjKzeT/m3lEM8l/DYPfo3RY/8bi3RYWAI1OyfHiBS3NhrxiRd/JkKFoO0YBNCZn
brY0PXO9hC8qOiH7IJ/fMpRVEJ6vK8bp+sDA6/Rfp5swZF58PY1MVVDBhFajmKUaaJbEdkUkUJ3P
w4fovTj07CX+gf5r3EKjp69f+FFyy7acoJxd9ZoHfDcWYn3RNU70l2xq54oONSclNsP8Kci2KxAB
7wgRYudluBC1rS0TPctHt51OcryvE3PlI921gDU1RAa2XPw4mHdT+C7D3P2vt7dpKZ4VS65n7NLE
H64kiru0TQTIO6goO7RYWRBGmw7S7hhabom33+GADt523EOk7IHCFmFCoNK9lzFH515XRYJw6rpO
p2DyaDYnySk3BSPLAFomURbqoX9yG90LQyZx42mA/kF3DKW+umsioguIgy0xuc1AbzN2jOxmi6bN
1OgQ8G4fiUT8LPpWjB8lO/7vd4us56hKvo8Wl6z1MY22VLV1kKfJqz8KZr2B94gL5lhkP8CHwcuN
IAJAAmRi8A+/rXCtDSQbVydUAdNqXVvbv9bBNq5hqlvHf4LmBKpViLPSqXncgOYyypsCghJx1Cnw
fGBJxR+sbKTtgPT8Uua3kuvB5vcQ4K14RNYDGhQ1hOiCQ3GdIATiSMDipZi0EYd/lKHVIEuuWyCm
ud3QIrVtgUvjvukzA9M74w77f31GHYx44bvQnXdp879INMLEar+wHyPyMnwv5CUopnhjyyTk//rf
Jml921a/3Z4gucn86sP5eYbnUsn2eRce07o6GAvjY0fo5dGO19Nd/L33gztyGCkyjvHXbK9HkGA4
lqvqtHSqXFhPebPTYl75iU4btyuf9/tg0BPBaN4/v4gkAjciCERuyo+G7oPcToL6clvyJM7zrGUY
185mUaU9bZmSOjE97FXYESBAW5TpHXsnRt3ytmuFKx98zQMl2FNM6QPonvWZ0Vnj69Ks8hZBGl8Y
h9gee4Qeqq8tWD4CwqkuARPdtrNXVTX4GX+Xf69EBk6jaT/X2KyzjnG94jUujWBlslkR8UHeXhje
kLcpDtQrsmuDwFzFpBYYAlwc31J6ksWiWgtgZ+RjQJWRYvAfpAnmqBY63I5+UlYVwbjZd66/XfCi
DFszYYq+ds3b1BC8Uj31NzWmXGIQMQphrFy5KUZnA4brdXt3rGFtFIWIg1nbvlr0ENqRK6rBqc9W
zGF/4oiPImdswhnxpPHy7vx9PfvR3PefX2VcThD7H233niRKMzLj4qgVBl8QROGDQUiORxmnl75h
cZm1PUnEfPdswAQnwcr4XCBQM7BlpSpClgRtOPPMQ4z+4I//Yvo7Xw15YQTF4YOCPAeWurXWlyv6
D+7CAMGqzl5A/7Poyktp8GILcLlzt5KuezNh361u3HQXBqBiw7moMHdOw6OQxAkY2Ycvu+DmyduJ
CQrOINy2WlrLaJEJ2IyRQfDA5ws1Mq02TPkyXlBEJjMpZuZt2xi5IjCqNk1ObXmCBT2wb8MQ+gtP
lsZbb8LPKfdD+CUyB4XlfYlcDl516ofjqebBaC30b8uGE/sdUhcNEq8MkMYfEArCs/YKWpYquK/0
c3v0Savrl87Kbp3HXsfdUbs6eKHeoC1CSuaG1aPvbrONy82JR8mD0706MckEOnzTBD7wsyfZPC+n
ZM5ESUEdKXmQPslCwQek1s5l/ol9Az54/nB02EihmxLjeYwpgQJLgDU4V86rTns1dz8+HAv6uT/2
VCQvkeX14blo5HPX6RqBJq7JEYBKPJKrD0Tuq2rvQPWVTp2uqa5wJEKUc/bRlwSLtMmW9L9ask2i
XBjbbQi4Fn3vptbV32/ROI+LDZ+oDepfVP1HrS1bXBF4QaB6z7iwgLx2Borh2i25UyWVtzTmMbfz
Ufa62QimeoqTi1HvtLV+Mle69FZJMEskQ92o/BiO8/WJBkg9CUqN2UbyBdcaim0uHOxrDnPtaUre
owNCGk3NJX8X+x+bJ+zdN0s0QKXxxuT8IF7xUPlTLKq1h7/8B3Ob2FgCb7VQeEsr/gtlL2yCDki5
0S726Cudlyo6uWln4g1O1gL/5myXcp4yjj5q9sn+tXAtkROAfnI6luQ3WbV0iAHklDHVi74vP3fN
3+x0wHNlc0AcRqC01gB91wcOIqK1Z3GO2oJW0P/WpKrcLqMJgCkHSZOuwsk3o7v6VniUg492WLcB
nmewTYfUcTu3Gf+7q6o5gAvuBuitYjCnOPdHCGrm2YSdrgoIedgJSPvx3Jpcs9g1kFdJ1UpejHTM
vyyTaN7FKlA7fK7ZhqFS1VAivpbnC0O47LtODmoVKF6jsv0sHyFrnIYS6bmtX/C+Oiiukih7EjIP
gAe1jSl6orcY0ZVj0q8MFmu2kTfi2dGAX7aofK+2aYmzu8uqxZyVntqJRHBSi6fLEk/jEtLjFJdb
ZAMssQYUB+106Vvlc1ftQJ19N5foFW7//kFR3kQ4J0osUorL2JEKUXDZ+Qx3JbscjMU/QOn76TJb
GSwtxwuBOvU/8Knr3gDY8IlGnPsqEKWFcrI3hVf7aK1J/WI6FaBRiRgl5mpoeARtne4TULfcx1wj
m53FIKirNDX0KPNr2bmVICntMzyJF6sZABaGorZB7jRP0QPe54vVpPI9TQ29C+CDP4qOVXYgpKRJ
F5Idnod0PyBHKbJKglsJZ6ZKvhvGL9KyWHbxqQaAv3cGync04fxenTXGvCUJllAg5AvTxyPLNTZF
fmLrBFcroG5K5CuB++5QqQqTWUjKjZwI6zzZ2QH4Uog7qRzg/65TvuuJHVKNzIJMoIGhgBYndM/z
G9w9PPnaV7enM8z4KBuj6aENNY1FfIjF4OSMc7jOO35MNfc2+5Mzj/P6ARlFN6Bu7xFPa3tQ+30b
WuzBGLIJX7uPR19qn69EuDeAIGc0mde3dNJ+CU3QF3pnDq9MVgvf7V1GbwCD+bz85Y29Uz9XxZmA
NeNKy6KyO5vgYCnm6vJEuX+FCvBvbA2whR0FagmRw6fh3If0bF+99Dij6j5tMBrYNxXeI7dlVYqO
owLFbWyJNkfw9aIdURj8a04brTRe4IThoBTp9DgZXmFvrM9vCE4hK4pthrDcaB7sUiCNEyxcnN2p
IbatKPh1ZX3lXazPnDFGi5jtD3xg8kNXCVUDWYm4/+3w1i7o4UBeyOLeo32Vfle1ceG6KuTHKnKn
Ry1/CfijWwcgD8Xu4INb8C6/duRDH+gNGXo08eGIt64BP5u6gECoAMIOmCiG7Rg/q/L5q24HfcGb
3qa3bmzIeRgmX267VWUIKqYKVmOGhoC75xizxe3rHo/Siq+RV9AM6B/ot96/1Gp4tQj3OkO2myDM
e00HYuO0eSxtGyHGybZfquFjtJ9g1Uf656qRmEaSr5raBgCENixxD98EVxQyBpkrlRju0YIGlfid
7VMwHbxxhy+mA9UETamFLbFX8yqp86y9SKUd/P/lAIWbGLS0mJFbNmABu5hxR+nrnxzr+6qWm3ZW
S1yuEC80NySz989Meqij26U7uRniJs6yNQRZGUe7ye1WKs+AKIUKUDJPBXCu9vI+/zzZQsXAY+T+
ShSF2dMaB4biy44d5rMI4sTxePDsdrLF13zwGzvfM9O5CNlxL31n/RRMmMR05USWQRsVgF7OCsEG
Ke714rE0+KNaiLwOpKKg80QieOjTYU5UNksg8Fil0d2ufa+o8Vp/fp2PnNEzMgz2Cb9s1DNWcxFw
JxwABoEJm4T2TraRvAO4rMbw5RYfXjC4reS2H8gFbM4qnFPM2t1FRz7ZHYYRWv68rr/g+4u7didx
1f06th8L8E7AHRIvuByqUIcHJfVlb2i2/WpQqV/L6E+afIbUd4HI9U3asMepQvPoOOmi0haDalRy
fL9TN0EyAk5PtY+RI8EVRcg58Bdb/AX1qHAm82LPfzI+QGmkgjSf3a3no9tQ65YRYkSVkJ4h495r
bzBXzL8Ww4b5vkIsZrrIYiTHqlOzVmXTHoSjHFgTLVuwlsoOQj9MOZeB1hyqeBuNtW4EwoFQB/QX
ZMDmEyO5xMDG0TLVkOv2rc9UxPPTfkHbQ4Nomv1WuBmCUjzkQ3QYCjySuLOvMif5RkRBy2bUEN0Q
rUR+5Z5ycxCdDBVpeVKgFS0vZ01H6ltiSX90NmETGjbyd37cVh6Yl2YC/9eVswXmdy4sbz5rsXze
6Re4db373Hlm59d2WxBX2gUXkTqdT0I/YphgogRXaCKRla7Jh46WQ0SIkk/bEjgPbIw6fDfjSulc
mNZNotDEBUDcz1iHlTPi8kcmsViKofWs+ED5y+oUlDo7PWNZFBBkLHEAWkrXspygkSuwAWYKs69L
V0yxd1fFoAFRehl6alv3cTod3taJRWvlL35JiE8ng0Lqa8+PvJ5w0+GcamZYlub56hPYCr+3Wdra
bDCjQS8ImNiLVMhaySVaPxYx1Vjygw4l0GUwQV5p1wkkCgbMXBjFx+l2U/TSesAn3dCjl7e5kQHg
tw5Mm2KYsmXZ/oV1rEciP9eEwn0JD9X1YOhijy6ZOrJrc93WnHe+fbrFr09PylQ+PHkcYyhVt6fO
LqjfQ16AHWEkboKAsuyxG8V177supVd9MHoKlUqWDRkbrLDuzb9QuS1ky5AqE6ocR81+NFYwL8J0
nTDKgph/VDF3d0BvCaUDRSw5UqVjUMU0LWAGc2kLhtByBht8xK2fozTqdGNXcy8qU31Tyn2enFJK
ZDTeunm8dm8oyRw5EDTp7Kb56eaeZHlU6T8E8N3ZXHtfGduFDv5Pmz1islXwceghDLFq+RCNvaAv
dicnSFQr3TPyL9cpCVtekoVE3oYaszMzZyz8jXyQCdx2KsSUbu40KPZFlbylpMp1uAfaAt8p+df5
FlhAct6SASC+6wwrdislhSgPaor/g9E1U8GUQBKwwI4OsoZmjE08HzspTqCsXPvPn/szJNDjs4nU
GPw0zuvwM7GvalbgvAvP4pUBCoQ8d8KXDzLLJsUDvCrqIAkMwvW3q340UCJ1tnsmrOQHK/LOHCg2
Tt9zruApijgxBQJIE/QR2lVz9gA52EvZiKylkchkXkhiW26PwVBRqB/HRoj8zg0IzchDZrj7Ab5L
iye/49tF/uOplsB7G8F6p8DJf9b99Ns84A4ff5UM9NZcKzQHPBDSSwGtC6GpGcxCykI20tanZrU6
zOaVzALhX82LvS6mVrt9GQHoR0pkRmSfHcPQmSoENGsvvPzUduaHDs9bib0YBCrla2In/dPfS/WO
8rg3M1WQpFPPsaS4j4+NCNwsFAWqi1/PZ0tPUGMcjrw95P0iVvD+zg0r13G4Az6ECuM087ytTAS+
ea1amKxXuBhSv+DHKfO5ecJaHKv6lomOO83ffXbk2NUtG5LxiYUrseSp/tCq7fDsAOAD53dMB3At
vM5vTC1TI7KVFQPqBeWFwFOB46S90aAWrxwRlC0mAWG6elE1InDInDtn0ygXvR0BUrGssd/o5Lyv
WQgkdiCyrTxWpsu0OQxHitM7XH9xnt/q97jLsEKQXYIWYux52AwlccSP5DMeoC2CB7/1O5yFX+Zj
w5WkDVUV68a8jGZH9r+7xjF9roiPp70tx8zh9n7tY8u7caQv30Q8aPiLg/BPYFCZHDrKAnvdhw31
WPlKxY6Re0MukrSz0fGMrveutRqKT0tUVwHFHLBKAaOX23wwLTFUJQlmu/ZlixzjGf+DOWi6B0sv
O9gUuXXcU2VVlb8cT66tHWtN4X7lMOVoRz8w5PRrC6ZL7cA8ni2HMs5dqepjs7WmgtFY6MiiSykB
w2pLhXzrw7m8aDyh1zVeOduCRcbGWMRni8wyGwmd/5snK+x4puqDEBE9AC1VNJjZbMjghF10wErw
40lRROK5Lk0gRtaQ1EDkKFAwOpYx62OM5mW3fAaLl9PQFg8GrJ/HTlr6Bw7V9ZqzgZWwItSbgvOM
RTUUngugd6UWBPLKDKE2XndhP/BfUlCdhzNrLTcCU1aI6JzRkF6+FhHWyAoQeNNDrRXbZMQKlbPP
N7m5BGI1GNh1NWEky6wer0vc5sgguJAEHKegGCkfz4FPgIZw/GpS74yhq13TRlL72Hk5mZprUIDG
Pmcfsv4bh0X3aHz79pAad8/2TpVmHKyh4qX0h8HUjpCogDkv6U9/YxBjSZhYuwdELFYUUJHJuX0u
JxgpegsaRWSzLiJp7Q/WeccDHZwsgxqbPNW6nLVJyiRuKISiEDkApvnrawVlG3P6RZVRZVw7ATk6
Q+fC1CWXLubd2u5HzCbnq8KsGknffzkgwmJx9wt7j7FpWEdG2gvrgs1EQmRuzIv1aYxtbRaknSXP
kWcaCj4njIJzkpXAnFESAORFFkFN7108jM6xya2MIbYLWnBy1vqVY8Z39IjSMF42XJSXfjLuissF
l50gWpT/uLXTzZ8BkoUxA41zNUynuXZfimnybCjLYIeFt0Jc2Hi1bkhNkaZqjTd9yCsM1ywb8DSO
D+c79wNK272lNGIVSOHwptxzIX9C8bfEGa2gBWpZuWoSS1LjbP5OlDBYe5TYSOcXt/UptYHGMl1/
P8WrqEeMFE9qyafvxgkBrY8IhD48G5ky/eXLNarEl0kYiEt8EjAlrfhC3T7H7iRwKtCy1ma64Vd1
sdmMSi4I5NY5XuwC2aq+xxRVLuv+My+fuPPJkCckEGpG+pK8HBZlBOFQqUWyUs5lioKXkZmpJ9LI
yIPe55/D7Mc2NeRa4JNE8TnPsaW0a0Xu3rv7dkXgWcLuy7kxs5XwvH+xLblEYjwALMRp+zpMrCTQ
+VMDpSFnxVpkSo0edH89rawsHvVOsUqgXbP7UwXNQaVzHyFr83cn2omJM8jHdAb6es24TGq/Krzp
svUS3I4VmOq8vwEOTNMNUirTOHqtM3aLiyh8L4I4E7HRS+hMuhd0XTZ2+WnYj+lDN4GBuuBRSrK3
sDPJy+m3Ejumbf1x9fAtyb9WH1PJ5WXjrpHwTdAQ+//lQiGDf+1W4AV87CkLI8lhoSTNAQqn2Ktn
dnvIZ1OiBJtLo/ojlJNxQFbS5d5M/g6NaD01sYUL59SuGbA5IEiLf033NltyvKf8V59vKOXF/qxh
/932bUEgtnYoTnlFwDbqCjam3lkrP022cANe8PaNc2hWRcjJbyn6H+qoCHaJqYPnE82GP0L9JhWN
yEu+or3NLTfysW20B6LdnU/aKxO5Vd1aeaq9lYVwGeRMjvN1pRonAb/fBJiuVhJEliNv7djEgLCh
u1d7wTVsO+/XMQlSgTwOoWXwc8aQedc83UAq3ZNoWzpe2SzGYofAwdquYD15/5K3BB4nhRXjPslR
uNtV3zLHFO1DFFUxS18se81ujO1Q5760zkhfQMmM6+LXoU06mLivmz9KYIipKV8vcOOdV1uSZJTM
yQD4J3eQSNt8W2MXLmk1gLgKgRcG3eFic9dk/G8Qf/BFMo7MPMZ8jypxX8AgS8nUy8vle3DPFUJw
AtROrIaeoW13gkSOWc56V8sJNFK2UqzVdPDYQpcHBEUg8zwicMGECU22xSbBSkdXcRlHQUfpU5r6
IGbTL5ataBYRdN3Hk657GhVdlWMKgFTpkhKdqsQ92xQwioEXCuN4+wLimP277UKLIKSpYhhMkMdL
qxoaSdaQ7VeFbac2SVrnktpgWTd91ZC8Bd8dpQ7e2jIYxpevjjIwbXYhAU62LVDGvji56+FBf0fZ
yoYhxP7EQt6MjnP1Xuc88tNioL0HJ59ek35xI/xMJy5cW/9N6361+vTBfuW4ho60IFLlqXOlYPa3
ZZGUqSPzH1BxFcwuIsMWLrtaUxBTjOoDg9a745tDDAw+vW50JghRr9zZSfpO+rfHF19/7tXDtti9
03VLI3O9x8nO6VC+MopGAkQxCPwTOUhn2HwMGcbot5RcmaUDfAr6LAiJ+Z6SoXn5eg4P8UROEYER
qGvb7KCqIgxg/Tm/FuEW8XsH9weelU4Wr1q67CPoVMjyQydqYxExalfXzJsU3IK6QVN/jjpP3ptI
vUu+URnl5qqJJUP3EoYorqqhZEnEyzj2m+o69c61ToOmxJ5cs3s2ffU3iVFfzNSw1w9bs7EazY6E
aC8tJCWnoTMf0bGp4Vb1/14aSbBgXNhaSJTS7epf9r1h6NY4Iwq6xYUmy/VpkqlK6SwDDWGsf68z
JBYAvcaOYSP143UKedFMYPeLXIcwdo8ezeu+hWS3ScKHnVSCbf1OXeGpIyi8ATlmRV5Y5ht1bnCK
A6QxOlEU4M1h8xI7hdXyluG9Eh2I26oNLprfJg6aBfbTsK/neNEL9eUBhTtw1sHAsKLEiZqP8f0y
Zmfmr+DPNi2O0d9Vw6IIpFLwOmD4YMDH1VU7fmRLEGUBREAhlNVyLP/r52WC3Zb1ZaqNTucbZbRK
hve4HNdFLTmnnYa3U0eGXhwgpwoFe55k7XrGSLxNV6Rt5a7zk4iNS5uDXQi4nM6b92t9QUPglzzp
OngCC22uTG8G5wooOsy3ZVELpNH/aUUTEk1yY/C9n2PuuP0DvKyEikCbuZOtp6+nVenIJrqChyhx
gbt0XH6BuiHWz0uBqsEcjusU1Pe83B0V31iRGLbvqesXVXfIRjNOO5ztE7lY5fQrCMM+KbS/bP99
1yOBkqYsoZBi7ei2ugqsU+odloKXSsyv8H1cE7UTOmEum86LY41X358avglNebATZ7anMwfdsKrP
SER9bu7ApmLS6++KX+YNBz4KuWulVQknIiL9JAU73MTrdxx+sZvm0f6qizpqphVF0SFPCLOhx52O
RnBoCnyX32qW1xfaCXo2P65mp2jgv1nm0bdT8Pze8OYumXPt/+HMJEdsXVRd7s6PBxW2S9alE0f0
Yzc/0dG0DplWYHUoMEDxJFwP6V23JWa3a6czJSQ54KAnM/0o6n9vS+bHxKB6TUrKm6BXmXkLmgVl
BrDq+wRAkSBEKGosW9AfZuO8w+TGb8fCqa8kx0J1NgeRRnUm7rVvLu4o5XFgjJZkrqwTtfu4XFem
eTRL1/YQCoBApeMFzY5kpjMgGeTK7SND+nlgGWmbtFfa4ZR2hB+cr1wzayPBeMZ8pN987UlVniv8
Ur4lyW1y9kFQEkvnU+/By0O7Yj0a7qi/EUyjqDW5Lgr/yfV6QhWx7n/4yfHBD2eBqVT7ZemLFHU/
bUZyRF2LYwxUPsIKXP9V+ZPQLEeI+qlEi0j/8Jt34RAJdCdDued/J8LPeSbiLT+UzTRzmkJA1SzS
nDmTp8gb3wdpxeXFw+tAk6sORhp+yobH3dBMEcRI5UPFV1guGOctvFdJW3J6GJXYt/qN+oS9VfEI
BO0Gu7R2WEOZU6HPkfPBCFYGaYx5mXlLB5Uw6wXLqzqOa/lLPqBgp22MIpMDwhp0W2CAfofoWsiC
MWpbalzyM15yyIDPh5ZN7vdqMVtXACAVBGLHIQVRzdiN9snvP0kCfpsBQfteRPwNvKkO0oM6P9Y2
bEoypCYfwT0/4zDdBU3kcZMEqmRelQZj+lU0Wj64bUF70PomWiRGdxomq39nZlaqvUMlRqb7onRY
DYN7ZuS7umWqhwsem5FU/ttH9181lS9sgZ22hLyPdnEPu7LvNxDNIT2OQOIyhq5iWd5FaqYwZycO
uQXNkjeL6HxdAJCiKUQLgiIZEa9EX2YU9+2g9DlSmKHTPp+kKpT/OGOUIbZ0NMORAXagQI8VbCUQ
5V0aZMWOeyvo9/FjLkfe77jxYUtZo62q9PI3z1IfzTsJFWKiVMvqpuo/bb7iWgYIN0sqpCqJzVJi
SNAkihL9okoIWWTdPuqw/Gf3nd7z14pqn8j/i20LxrLLb4eVO+mzGAsWD/ZOigaR7LX1zG9/H8WW
AChEOb+6zHRtc4gs44Ad96jwBh09k+4oRNO8nEzyTvLePaKOGAFkKdPIZbWGdXwYoOes3f7244zB
UCr3K0Iu8CEak+Lw6Kf+wHEetyrxoXKnTjHwVz9Nleax4Lpwh0eG7L76rXQnPT1Y22rmbsxeX9eu
35gldduOkX3K6DLCQV5AyCZ234SF0x+z+s37shQUNWPARPKVuGn2a9I7DtbyoK157YQv3wR6/dVg
tO1yuKqh8waLJpKbc7vKNEl9bOLhiU6tuMSMsmCUoT0Fx1fBw0ADwoqzlojSWx6WnT/DyA8P1Y4H
gD1qBD+riPm3AcSF8hEmfjvMvsD3Qgp+CkMkvN9PP4xPUIJYoBcJh23Hk0NxqZ95OI1lkrDvfAcg
xXMCHSdjrIdNr18Yxkh33lGzX8MYTA1fZJ4PxRXXnS7/qQub16Tfkx0eYL99fQ7bU7rgvGRZdHPY
DMzVJj7KRTdt8GdodFVpa6h4UNTJEaLGl08LvhhJXfXo1NgMn8cNin9vjy417dsX2ESsOMR6O9/W
2gSiDnU30fa89ymzqsyuBn1TIhtcVtWVy+CbsPwnd1XF8YRQdgBOoRPuezTbclIJdu4RbGBLyKoq
DyGk6VZOUVSNT03v3tGYAHThA9XpeFFkpad41qp4MK5Am+vmTalWA9ufW3bz2P9+rCx/aBzfl20r
0KO0oSFHekpMZ675Aq3Bz7GPyT0tk5H1s+YmxhvuN0ZdaH3dd8FTjlbVyg8JYhyLvoBvNG2E7JYM
RqfsTZRFQtZ2Z1vCzkIS2+6QQBj9sOuLi7etAf0mU7rrZUiXhOSz1APh2UWsT+olU3RYcgf3pwF4
yu/lA+GVlumNfuXBoGRkI1d62FXIFaxhpxrvojC0kA6frdukf35DnQExt9ED79HV6x0jSTUmqQRQ
PdjbadPbB5HAr7ZzBkaUHJbBSx8r4mrZiHbrpHggBpon8GALLf5pUGUfdAPfM/Xv3bNhdrVZOUjj
cRqXmHWRMkuY9PtTsaC3g0aajQ4u+LWYcA3Yg7K11anFsKXBQFEpR8JmdxrknO0FrFoZUMpA0LWX
XtiNiZSdFcVhN6ETwOARcE8WsmmQ9ffwNMkmvEXXRypCKhLi6Ig5hfpsL4SPne6d4TToQgxBwbcE
x1KtSRWHUbYer+IJMb9NIk3hOrSM0dQxOjBgKioZUcVJ001oyHupcliJWQihUZwt33QYP+Ym+2qq
LI9Gf1vhIrsTJS0Mx/ROyNFZiXtZlu4F3CCLqed+R8nvfDZy8Z15zKHJWvnBXZabT3VEs0M4PnMs
wKI2Pp252fcf5GFP1dgMdYDIymfSdwBK1127l0zVMTJONKvKxzcNDsSCqZUdex9xuc1A26h1ykIL
ZWcXZ3SY8+XbLc8DD2HGapPMmgHsO+jq33S356ZaoOoX/aALKio/KkOOvoDmoC6yx15sxtgZNSza
SL0qaE+VDK+atgDAMgLJKVt5uqOk2jZ+EFXSgZADwtTE8E99/0WRAsdArLFRQJGAyAO31ZuxQVyk
2PS94ah+fmgQSo4paA/G+iCa7EADE1GOZOV50b7HVLxSOtKc4TZbP18KdiKkB4z2KswzN2EdAa9P
5byK4Rc4X5jKonArM/Dgxft74oYf9+8Jl+06UjE3ChVHlQ6Ewu73BTMIZ6ZXNqmxz5/b5hgQ3BGl
9fOX+bOaU9XMxrW7n6WVQU55CpRzZgRFN0qSJPavef5jajZfFOEnIiJF95k7S5/J/bGNj6qTOc6f
bxUF4OLgeQ9B1jh9M1bEo6XRizXe7lIiUCnNpXUTgbGtc3SpmBz+8at6sPD0H9rR/bx+5dmaKBmh
Um3t15WwtsoEtxWnoJg6uBgFZeBhGpzzco7dIN0vWDBWOLO/u2LGH5n8qc8LLJ4mPjDqPTdvwUk3
C/TWn5E6g9tlQIy6m5ZJ9KXNc03Y/h5Z1+Kfe2Gr9LDnGD47sWKhuk3gJlcvje20izhNXUMt1dqq
quJWfAbVV1pplKbPCo4fClRryQ/plGs4JVFXjZtbrQP6bGvsg6jN22wX8kbd6A5uqj2l4rzxNWZ8
SkRR+NyhBwtZxpWow98UaVtaRDrVuaXWPoEr4764GRachiKxRQCp5IpVj/BRNZxJi0p9+Om6FEnl
rKThf9C38+NTrF7UR+DD/LBe3u+P7MyDJNdaznGuYcwhqh3UawEuX3rQPUiKO6ZIndkXSHg1Viva
PO9ZnkS2pDdyTUSDLuZHLrBk2LjNKUpxeclMzVsi+LFk+wocOOl2X4VReo3mfyz5DGXPg8+NL8tJ
SeVcSXv6NfTqGZSSJ1AHZfBW5E+WiZ5ifX+Qczr2nJlwGlKZ3nvCa9rg/U/2NDGMZgbVdFMw2yZj
mzy8joKloMcdrL2Wri6D3lW5Ip7qEPcHpWe7TBNizDBzPSmb8KCi8hFCGIbbBX/PXAKwJCZfFdi7
OQN084WshI63xWSPXO2ELWkf+1byfgXPjY3G5uiAssV+UBY4MVJJ+bDAN9sM1aEya7QqZXm3J8dO
VIOlRz67c8rNoEdgIpVelixPXRzpsQxDU0+14oMwlgc4bOgqP7Vty+vZL1KeyHmhLa3+No89cZ5/
+XGhz8zjWVQmE9W41JNRsgtGHonLboWruZc6l31XdEDZ3cbTf9Xr7FJrqAiM2rMiYSkrGoYSwxzi
Dn1qN+XbBwGB9SCozqFwQPaabT75JfI122CV/qJ37edzVUL7LlHq9fE1h6FyiY8mLWLY+xzkR/9M
SCnn+VxrMB7Lt251ZwJe95ZivLubR2WGm/mCp0FVMd4R3EiUwU6tl7UuENRA3ix1bo5VJiBIVtNX
V+c8b5GhzcfiB8LhJ7rymOQECMoHX/WKwlAHadwvTI+ZGutECdpIjZcrg+maDE49A2ZF/110jUYu
dnbvC0vuFEblNonGKMTif1OO+io+8u3tnoh5pd24/LscH7DzYdRGROitfspmXk4vXBtkR3lRHnzv
fDe39S7pGtkBgagawfe1IjDyzP1r72TWBf339wAHewr8ZhWP+AC0W6FS3qRtCdKNzA5OkXHtJyGX
AerQILWN1we9RoqPVaG6DonL8yoP33UAemBjLN8nYKo2djwh7I18JmokWlHoq7lJI2C3uH1HPC2f
WiZnyzAdmp3Kw7I4y1T7mZoKS/HT8/M/AtKsWJoMAOQED7NArrsGEmjR9kAPTvAZnchkRUXgH1VK
fODKiqOKyVG2d4sbFhT0OqtUHkGvoAAPZAQHeNxulIcShjsI5xBwdvXS8vQmudk10IMNQqaHBvzi
ypoSQ0tlCMwRG3Ulj5kIkEPvDeumjeMSd1J5aV0bkdoHrFDhIIXyYbt1PAK5QxkEepCWFpIOgFgH
TCMpMXBdhTmaMb3y6FRnyzuyRuPnM8eQHZECfJzMgjZkq3VF0cwu9ItJN0SHVbAEXdBSK3zFfswn
WzAAVKu5J6b8VXSJDo9rCsnZg8fHDBPEV4ooFc068mRsxjLFl7IGSSdqxnt40s1CnCUUGJJ2nkaQ
fNhMGgfMSMCWFDznu/3IHcZc8pPkJY8TaUi2hFl+yLOcZ7Qk9/a088ye3qs3KjMhwIQ1LuCBHyHt
xGByEw1kFcNTxWDlGs4WELMNKY6KOxnkeE3hoxoes9KOaIltofwGGGwnm5IFaPVhYLHY4WxT4fco
/8I0yt9RqvJarbqn6SMWnPCzYyl5YUP+oBfaLZj3GVCyA6VwCTlyVtm5AIY5+AzX0uzGWF3sMTgg
tJWpCVVJqzoW4aHtRkl/rarv/aon6arOY/i/nTrOPozx3gXI1TTE3pToL5ZOmQwzjzZci85gTyLY
qvbFtuwB1nvwy22fO/znd4BEH+SSEVymKYrhfwLlEujoBnxMQcyGQJt4LbAG+MRQFW6RImOW1Z5y
vEw6dyQGp/kiYxu8QNgJWnVAZ5ncPzJMQOQZe0hUlh75pDNWlDn3/WRP8AzNOugI6mvJY3kdsCor
RYFH/IQXIk5Posi6w16jmZ0YBSLmELhRLCTofEGXeFT0SpPkMAKwubmeAaV1OvjbmYxe+AGsbhy6
xI/jngIK3/EGizhul2k9ViwtQOm0UA1Q/tRolxdergwUgwZ9Q0vpRNgtsPbqlvowsilBJh9FRg7L
y0GbM37ZpvvS2JDs3y0xKNIFkrK0boVLObRl2liXMg9Ty3W9WGLRb3+qZwULNE+D0vu3ST8XeUBX
HpKQ691p4TjXbhxvUyOe5OP+oNu+PZVhgl0BASGa+WpPk8CxGSdVyC5HD6FUQ++8xNyvO3VTQNi1
eCZPWrYQbtCn6m2pKPYdxL5Dl3zJJW8x9wuVAh9OHPxHu56+oajbVO9xXjWR8uHwEuH7gXTC/O4q
+1QQgh/TtW1x8KIyGfNonwhP1YRpZNtG+kOkSF6SXdSNM06hzENk2KYAKCpKVqSUdQFjQJlcQMjf
bxLI14VD5t4n5KpljWU67UxtX2kldFdbcKwUkfSbO7yK3KWPSCQeTyQImF2UVK7nObsvMs8ysKvU
x0FpPVVMAJ87X5qZRa6ujYuXGrWqDHudAq3tIrKNRmAi1cRrpeqU17kJOTQntoFQamvsjyCOW4/T
IyuYDRixGxrPIXyeiEAHoqBCWiYWaEq4LHS4CWcsATaQ1xoOybPU+S3jFcZu0We6J3utuIf/vxnf
XLYhJPHmHZ2D8oeay73ibUucaxk8PtuLRFgmDTMJPAMsSrS/MXNllU3o+YShDLC7Sp0WZhpvFebO
IV7rV7fX7az1ZXhaZxyilkKLQJ3jVqk4MiAa4zGa7NpjF7udDg7uKTYt/1z6616pK3Vd9sPoNOK8
0QmRxTu0eUS+VbYGA1AmnaCSMQfgH7FncriL6sIj4Ara8rKG/FcnrCBqOgqEd5poDrxtrytJm2ph
XOvsUVJLcC8334f5T2UsqQYkFwpAm+VE5WMw4nAmsGaZHDx+jUjziM9zqMgOCdu+1IzfiojR84jU
CUXicz2lZKix6Hstm6e3qNISlh5quo+qLKql0qP/Z5gOvP6OLn1XvhAfyhXPzrJk0r1o52HDfLlv
K6vj3q2myHHjNIytQwY3e5lEaC2qfiWT8DEnqtYJOY0Ks0gLjaBjFBalMD+xMof3QE5tBJwmCaW1
41iFE/sqWcvTmpDQ6PPdGp4pwgyS6tTjygfcVbQoCoa4Armi7BWC9Zr/YFHGddnQLNRD2ZX4/sOo
dg3nchcGUejK1tuOkw2cT3hjo7l3z9moZnIb9MgelHKgUB0vNxv4Wx6W/mmT4kOsgoObzngJ9Bmz
O0hAg+F10Hh9bmXuifNZ43Ndtw8jSVEmboeTMfLZY2dF4ZEI8XRLmgD+WwED1/SPueu/A4BsdpGK
7H8lcFioAXDyHn8AyqO7qsjEXs/+Bu1B7y98pkHV6dcPhYwibQlCuJxAsQ2AxvUi+/ucEqf+zVo+
E0KBtRDGnogoxt7xpfzHQUNqRwgrmJawwCFGXtlfwCqJ1I3x1I8u8IO3J97CndqYynUrzPEnMW10
o7d9YvlWakJ4FmJjLijt5BVYalXr6uqkLwj+bQEbWJtNEGYyHFsEk40kmhocExo03zSlMJggODvT
E7FC61cxjn3MwZYVFmZV1/ArB1WOCTQ56Mq+gAu/o4QcESAEsjpTBW56xgJE6LCT8l2ADILMZ0rS
UK1SsiBEQxkCe9QSzc6y+Ks6KaPh1NNzdP1CswD8r1iVtmcTBWSpsyg1CWhpG500S0Cko5qup/Xu
ynFhsUqdLHkv/o6jnt1eVRqJBeg43p3WaGm9NGQfeER0Il6YVAS4A74Kh6L6vhelgCviuEFc7v+3
6bTzEH8T46YnElQ6rA42wjm/IWT3Mab0exgDiIJrygC4b00jfIfWVH3XAkos1Pm3sSTFwIcQ/E56
p1aadrOPK4TaxeWdRreiaoVdsKkb/zD/uz7JkRPHn1Yg1c6OazWrHJi5aYbtIz6a+Z6Ju2kOpD0c
3LvFU/JKk1Ae20XEN/8Az6tYUJq7rDzS7kd7l6CkYMvkHroZxMS8ElLBzrTpZGP8imJhgFJhCuUu
qdbTl9a6imag28+3u0izcKHSYhHDELO7IVt7sgJjbXFxGWR/ryFhKcnfS2CsGX5em56Ql5m9rzkw
ajPDmzyXc9sN2xgpkhNLhdPUpleIopzIc0FIiTILz5TIl+DpOFWbNrlgD29KYNsgdQ2jN4EjZAWB
VzcxEgjnNJSaeVQMlbGyWBvOnEYYDsjhj2HsRId5KR7yjeoiB35bIVJtBM4kQkJ7lFOaWWoAUM9N
5o5I9mfiC3UVHpsbuxi6rcwu7xqscm2x6bsNY2mTe/gvfob81bFTDrNVtv74YKMjZuiSMiUDJ+Fy
jBi5zomscSyNNhwnkk+0R91JIPKNg4rQmCtyN9D4JEHRa1yt/FiN5aBNtBUxiZYI/8Wg+OJbzFM9
zeEJgZqWhrkHcmArZLLXlJw5+tHXQhNyA/opvwd4+wNcrsaQLbMBKahldeWy3fgNkmlIX2XhZX/b
sWNd8MdctpT+Gs4HkMc1oRnN0+2uiupcGrFbPlg/fIA0wkXi2CFG/bhMReANCanAHXHhzF92IUab
WB5PU28Jf6aYrSVnoSv3oLMazJkX9OMUePhQ3okkexnJq5108rKVq25dLtzXKrQqip9gr5NEgB5E
EqU22fGk6PrZqxdFgY/ua25nOgJrxMaeX6Vo3cAHiuuktdpbGCiFcGLsq4sVW+ZAiex06Iri469P
eapGiqb9aorBSz6z6V9GjNqRF50Us8tjvK1Ot0bYfILN7FMrdJ5nGOru6V+mzeX2u5aMUrDJn77n
P0sRVN+vxIBpGjPVCIk7/j9HkHtx7he8EUyB+AjjIWDoawUw57pa0rA71dXY0yuqLfKAoM2KG7w9
OQnxRJde7d17lxo94EMuucokoWVxVbnRrO0nmc/l1vqphwntyPbXVsKSHj2MYhNcLDfXI2kqRSF7
XY8KTqN4CUeZuCZG5wM1OoZZBPytsLUwnJbS5G9s9LXSFZkGsnyq90NTDyZn7r9nH4zGz2lWCYe/
CysrK94mLnXsgb1H3y1smdIQ+kdjmLt0aReJDclN/xFLp3gSnZg/8PJ4RF0ysXU8JKs7BEwzoqGs
9+IF6uLlxPIFAKIAzV+jxmJk38ALfh+jRF2Qq6a1YvYCVJ9MgxOZM+q0bDsBWebXwc9WZ25WC2Co
sp4FtfNWUrdnP1HTKUYV8NcWcvnzjZgMY0Wim/TVwsmLg5fv5PiJNUUQO4n9Y/Kqp2AxA67kbqt+
AKG72e5rtCaOVBlbsi0w+47V7fYbnicNFvgOOarQICtEjkJEGPF5KPugYP0GHa62rgQF97fwxOqc
cvV3gVgzc2ZY6Oulx16H4eH7SxCnYTQZKihtevYwMx6zq+TbxjbZIpnIT0tT0/21wdf/HL9cPzYP
In2GmYy5JoayezVkBuSVv7s9YXtqsSwrnKGUznnsG4dKdNa7KGhIat/DuvvBbnJiThv+YdN9qXGq
0qwnTQvQlZxsoxrT9aUZ6k9EmIHRF9CQl5F/kFf50juxiiype2Qh6W6vXn9xv5eBM/Gr0YBDfPtR
atp+SuAsExpeElS/xIrMQk6wivRN9WculZenKYbYDYSNd5x5q+me0B9DDCurn/se8LgtmTlZcYV2
xIdO6OE9QQzD/kul9JQeR5x4hF+6S/R0krnMuSjjLrmlPBEKMVoxEJ+T0Dhbc63rHuDt9UI+fviV
l8Yid4hQQNq8DLDUya/1gk0X9UP8iVb88mIaQUgYlURj+Hs0L3QSACsIU7YKCtkYQWTsHedF3KIO
GHhUaCrZJC/MAX1zCixQ2hFu10SOYR2nz3tiS15z2nr/Cs2NQ91HMv7GxnDKQkhxNKwmZV47Xoly
s0xsIKUk2uz3upF+yIF4uqWvxZRaOI/AfNCNDa/N03Ugh9eBv8cYqDMz0Afv8z6CrZozVCpgPp6h
kfG1VvSjDrGvdNAGWKpXWLyMjiWF9IkuNYQue6aCBbO7GTFtuaGMGAITGWu1l19ZIb6+/iCLIVL5
eKcjlj6Da/QENEDfGysGTZmdeo0MlakiR3gQLA6WtrG8n/t8QXn1nO9MeBGt7to0jvuxBw+J9Bos
TaOqwFRib2D99a/hyunZruH4WVKZPfNrQbcComUxw+dwLmH0QzINvkiuaw9O2POqY+En50G+8u4p
yKqQl6xhj3XhhBEQqgoW92ByVGVENYo/0G//63vCFATY1qh0FSwO4LaMEY8po7kl0GHLiGdO865d
BiJPUmUHL3CC284IqcUSaYA2Stfmhvj+mNyGpf+8U3FKsq/2/5punBOL25VZlFgdaUGR5qOGpwc+
mrgZRWo8osYpIBRfb7UEaeKLpdNNo6+UstqWK16WUY35UqqjyoRgNUUJnv/XmZUmbiUjEhlp7nw9
bH/jjlHXantb1Yxm7hG9E+oQCJhMix++RDp1pY4joSymxMJl0ZywOxj7W6m9a9joL/M5rPl95Ua8
ynxwbZ7rt1nXS+vJ6RORSlqGuaW59QClxVDx7CsFuHthljitv20j6GIFWnbnTxYW3IWKMz3l/+WJ
AnKLbqL/a2gDB0YuRj5AYGKeBqYDlJxtoNX8wHsZjEdIcAIjJYubIIut27zgrOv9zxTpzbTh9YEy
SYmmfuKsRcvVbTFO0tzBVTHIp/+kkkwJIIPBQFLc6NPygxrw6I87OzYyun/l0yhfoVxV0elUST4E
NkgY2XeYIIzwPD1DHK877wNa7rxLMcpTsqT2smbuKnxuhNAR75KQ0NzPzM/AlL4KhPrlpRAexyt3
H+zS5PR05C2JHUUmL3GBhodj2oiQyIt/6HhIBoxa9QV2Y9YDzup+HLtjtzpjvuRkLMmxIUB5QUER
UaGy0Iy7ge3OkhMdOtSBlFxVStLd2/9uzHH0oZ5BrLMj0dnHr2Gj2NgrSCV+tO6z7ujXYoE60ipU
XG3iTCccjQuwr89NAW7GC6LKUpPqVs2pRXvZxLf0Fltsa7zhzXsVXOTgRxBInpPptYFzIGjV1roH
TXD5X7SVDWQmLOUdxqMmP1ltFMiBDvVPBCyCJbkHKLuM19k18DOIUQuQuzb/j0iQfSS88TXWYf8L
Zkje+yNGixmm9lPcOT+DO0qa7C8iazBUVyRYPvUCeI7WIGa65T5fa8HmZqPwmgk87mDnXdWSJSdu
29ScH8426KSM7dcotGcAixzeLBFxMA8Vq04fzPgGTKbcSzPFNfpkWaIL1J2aZDqh1Hz+fFA5kGnJ
OjZJCKgbtiVj5Ys6Oj30HZB7dFHCQyiC6uSk/xe8pqj2LPiFDyx2ZisJOTCPol5OpVNxfuVBsotR
jQUa5nwhsQFPg9jAjhYG7XOJUWR0qscGmtqX3Qj5N+CQIRsw7BxHfQ7cW3ZVTc5Ctc/Doh8GmMtA
2J2Gr3MPqq6V1hOZTVhm8ItwEyKfZ90ewIr10kMNDd8oWWgUEYTQ4LDcB1uBkzAIbzmddp3UkmJ7
X+3+ZG2z5pBYIqKABpgfGLHE0cLA+WuM3jmm7kVyU9Fyfar1sGjKqPBCttmtptrpgYsu6yMA+DU7
FFntnUhM/NsaDYwnK5CxE3iwJBT0OCUQr/3tB90VCAjhBsqxKu5W0Vws+eTSKJDh+rQNoCowXmrT
DqfR/Me901PlwI96zissTFv8f3mYj/37FXtRMta9ZGO2Th/BD9QmB/HdzXxK5fwMLuITzAf66mGx
BGsQ9WuCUBcSOTjD4v24GO94q4/xUPL04RxXmBUVM/a/AaaREYuSPC6Uu7VH5ipRqJwMvPb6UDjv
33cBpJoZaM5b1dVjqxGBwMhNm+xuDO+3zLqqL/5KTvcSzLbBbQGdU7F+mO/TJvr1k1p+Ullhzhkr
7+F9QPUuSgPPauh9PRy5zFIDL/U0jH4LkPQreTat0AUCgpp5Rfk8Dp1RL+ZDLxpPKIb95pHlqRRM
J4oPI6wSGr4PUe7YTJgJNDJ4wj4IT1MV5wiMRg8faBX4RKKIGXpeXANmVKVa/N3cH4HR6rwZy4IY
6qJkps740HWsHI358TyKNQw+mFVQCQpyeEUnVBvnwA1dNgbRYdpTQCc3d7ICXmBDpjuBv4sKwWjD
5JjaxI12gqKxc7QfD+aKOirH8/zYM6iGBSwWDEmHx/+TSlnE8PQZ11LO44mPhf+7yvaQ+MEK0fA6
ZjS6aEVZpk40DvctO0TLHnFonSS1XkXmy90zNVOaig+xjPCLgf/9vsSAFlghL74T9VxaIXeaG1L9
Vt0ZBEqpPBDRKrWmSAx/ubsqqB2p/xSU38N2zy97pl1Jx/tyj2/ay2d/8iLLVYrHebmcHzDui6xv
y+Zut4+m8BQLXumrYSkJhxas8Jr9TQlbAcZt85dg6ieuDJr9wlSUFcu7XRzPokV4hyOPLZhOME/U
f4cB7rQgAkk58d7SrUZpGEgtYeaj2bEeq1cdU+kobSGx7Zg3O6Bmes8gBTXuH5wQFM+bd3aDIWTW
ngUCeU/eMHlprbC6N4Ela+MJHzfW5NTJS4Tmib03sVaAl6ycINftsz5ZzW7JIZqkvT7UT0CEuM+C
/aYXuKxLamMb5sSI4+FASQAGqj8rVujSw52yqqsWMzboWn2DzIDn8RaLslcGM3fS2n1t7vsaMHr8
YGuvBzLK5mLXNfSdgnyVguDP1Dw6hDBxufZtplovJBxUnVj4nrRgs1pAKVW9dxIsBTxT7L3DD4dj
cCb7OUi4uHrtycRx+5YnijXhL/xIt/p5FBYBh4COxmVmHYL+YMk1TsRie3tTF/OhU2D3orcUTMaa
E+mHjzuf1EYQduYw+SFNAPbQEmI+wcDM407rL1zTFIef5SLSJIzSPJ7J67R/XyC7ZRgmIxqIdvsM
BQ0pIHcuLiYBeGZ03chDYQj47GNWLrr9TBva11InJ/0vkZtwuMiLVJ2kYnqKS/VSr4Zoi+B8QOEm
qq1e2cszF8Vtq74TYidZyJbRh8EGqliUrQmOLfgS6+oBKV/SPOcnwXt2xJEOKhgLQ8m+2PcglO79
fkhuMunqLOEkrXN2jJ1aEP32/COSdSN8RQr9hj8SNIz7K93D9FXF4n55sKOtK+3nqZCVLHAeVETB
Fl6sQAL+BO/mh6lt/Xv8Lxs/0vtlkfPEW3DAonva69jeyiKJ3Ba/ykwmaSMt1sFEo5+lGTS3uwez
JJ6PB1JQG4ZVVtXlsG+9CISARzcuhXit14ETe5xMR0jX1Fvlqvqz7sfgJUZBJs6lGqr3cm+xq6wM
S3b0lX08QfQ+UxPK5eYLxv0Sj/OFHrXrn6w+SRpXUtoHiNQEnPNVhlOJU5BoGO0n2AGMY/5crwW9
rLVYbeVyuh5B6SJU9Z5VKBBd56TY02gGsYucKuZllzsTt3pqTmjYmZoCOvukqV6J1K4JIzguk2/C
G8IvYzy+XRu3Tk1EZTdpbgD7VE5t+lBiF2mmmKG5cSeT1ALqE6wLPXIUkeICkTbZFjyie4vvNAFR
uttzPjmSNqFAOUbJonJUtqrofqp1UJ0KYxKHIbADap6qpktXSea/V5kOeNbTnsOXQ32DUOx719Vb
d1tWoDIw3upd164qyRwe7d4K0+T1jMSPaa9wgbiuOU+k+K1ad4rwoHcaw4fZPRDZPelITdqXCmo0
zZ2oZSV/BmrPDx63Qc6FVfW60UGIWKs08nw6pXw0Ht+V/j3Rk17sCgmNbg/C3e2qr56ZciAIDFnb
DBid7HdA5fdVkiJi3dSpIMT+FzFD/9A1v4b5pxp4rjzx/iorPoCD++zGARaHbQVBSU6Kxy0YWb5U
gdfA9kBbLFOuTOYbleuSRryKWoT4O/OvQc5Sn+/l+ugEhZIicfz9w8XEalXUyDRukJdA5ec9ffkW
fiotXRDbyEbRzWOXwT+OuE+KxaC/SvyugsVBrHeDGfZ26G5yfdYq4hhFh9L4zfOeLwaaEW3O/273
eOLYILccds+GzBzKFbbsj7BRx+m++1SRfV6p6vHtl6s/5phS6XalQHpyn8pJJoVAQBO/7sjz3FcE
QxILzkXs6YpXyqO3ySbWqLETdfZRLbSV9PZ02oAZ/AG//d+8v1GAnrdFyafO81FFVPioaItZtuZn
oHpfYRIgoXmMHTFDTCOftIDgBCR3/CPnYt9gxUkNupdF9l4mpJmojLna8mUV54Qkmy/JxO1icIpv
TW3rpxOCaAbtoubWQjbrZRzYG9C7FY+eqRX8eWcafslk3eizO+0FPuMNJ6L6Bou6as1p/8rbfF1H
olsFDreoz4lsilfxDu0tHtAzqYUQcATdeP2Vnu7Ix8i1qUM+qYpPSa8WTujvGlrQh1+jhZ3Ng4/f
ZknIkzq6fkvlX12TKwW5/b7eleKDWY4Slti3N4ZgBzozAqDKz22CxiiCLiAPBWNXGwxvZe7GqaUp
O0fcZPEhAXOF9tNygU8+Gwlrghpf61sab7vGC3ClihdWfopsB3qxUSpXiAuNAsb7b2jmlHdsnPvi
vC9Q8AKH50H3yBER6IlTs4BghcNWnsSFhcFZzelglbVGuFGt2EUn6xafrzKz3uccVf+FOCckrocr
0CBxqrtlhhAFM6m8TBXowH+DRAUDpBegdRZnCzBXOvk1feCx+G9YINmKTZ+dVoFaMUB+CgDQYhaJ
gL9R17t45ABhlzvqWZxDSc8fU+mEvRFbZdm3QvfQ8Aw8EMVuJYHNtZZvpsSvXZ9VC4oZKdG4iY/x
ZShMPI3qLimMB1kHngIoeyJbSZtf+J2KLkklptKnt+2daOOSFZfPPkr+6GJt9qzGEicB9UYUY0dj
PKTZBkKWLhpuBVq2YaYX7V0cwS/oZG3zfRzq2WaXuYdUxg0tbkkNmq+atgiqaY4LdcWpHNP4WXWJ
u1/4lIbyaV6Y7KrnNJPdtWxVw0YLAxdjTuIzKtAkWZQ1dK6dfwrIXWXVJFqsqFzVSW1O0HrWJJb4
DT6EO01EwQydRKeEZFKpqgeTCDd3P5vf+M5O09C05OMRSjnNW/08iznFwtAttVHTy8GXY5KhVxvu
8Wj9ZLz/myOPrme+NnuY2N8uhKcH1I5u/96MBjFg3dYlRO+bhu23yZJWixgDU3KVYHX0KhTg+eyK
tjg8mTEoa0jfa4dVZR6KtoKGP93Zyl2hDXunKcDQZTe9VPn59W6vx9Rk2pUULYkM2HaFWMuq07Ff
YkAcn7uRAW0wltImoAHTPaLi04QonPC3w00jDjR40JWfOUFLRK44ffsi5H63hh/LzF1/jVePJjXl
Z64iIxtwHCh1W49aKztIovdAm3QW4ZqSUcmu72a+jGlnHfM05RPlIkaepBEidLb8n7AKosGO2Jc7
wNq3MIaG3S4x4/Nvu/b+GvcJYugkju7H4t1KVzuF24VeJfIhCaoC0F47Oc7tj+aWQ3Pu/fp0DTDN
btQWKJCSvqVZ2UgmGowQbY+5jtEDvPhoULZVeTOWAspnxPG5mbpn6MqyhpcMBoLIX9iJ7Yiw9QOR
PT287ju+EcNcFcV1miS0rlG9MCOSe6BUW6S6YeDtKRbUu3gVsP83rYn0CUscwRbbB47zu189X9RU
uX7xYgqXh4ZSnxp549w9NJXFz7N3aqdqJ1HRf2KIFrPW/LWJKbisRU1s9vlGKuJxXdqcfJuYDltE
xVrHeTvL+KuFgtQPGMXwNKFd+MWOjl9gG7eb+tmPaBv7Ke6y5UL9SlTIvZDERB4RI5rOmL1eZAfJ
dDz16c5krowEPh8JMvPwTnx0swFzk4cdZ7seMUHemsJdZjYhuPWruHkK3ixeA5TEFaBExbfo6SNM
ciau9Np+latttC4suJBNHTw/mE6TR2esHkyytAovN9QUwvdbdZlNi1XXg2GQMOgIJrruTYxBJXOF
RXutXzQqvAGq8UHEhUqr0pLg9xQU2xXj+QMAFysr9cCys1m7uQ5vOWacl5J80bivS/vY+rYZFeAw
qxmrrSf4DZegDN+mJ9YA9dG4i/I1gQ2ygPMVTvy+X2SWEEYCgggfPIYeqY97BQUf3zL48gVly/WO
1y9tBV0c3AnLPFheoYPOjQVi1Tu8UzfLzSgM1xPcEOFCBAVGpAgT/MA/Dr+zO65QvX/SAyjaBp0K
ePencXNwMocU6aRkZczr0myz95qf+0z1ih1tiILs9o0XCPZE3kArdVW2gYxww8SJ24SxBZ5sGxjK
m6sZ7bXFxmFbBeXcsUC9tNt7xEKwczO+k/sSj86hHXMq9wgpwwSoC+CwJoWsC2Zff51hgawvZIuL
2M7ZxgsQKOqXo2aCYCJCQ812uW35nrK5ea+54luid363IcWPa5KQHdYIALeb4ma7XxMFmHqiptkc
0ES7UGdXYy0iOiolhbzqDL9ybjgmfsf+QFuDjEL1if0cv60d6GvNjQgzuPq17IMl6etfeOBLEYO2
JgKnRBADdhFzpBBYrJsrnVWWC/WMWaKRIfJXztJrr9bF/nslrOv2A/NNsj5KUqY+HJHdZhmcMA3G
Z4g0Biu6otOdkBiXM5sIZiCL8qL/FVoRiO6DGuMwcuHnFqSQ1It3NEFyJXqUzNcRPQnEH29JgAKn
Sfu0JZnoMjxUz9mPFMPgCWf7qisMH2c7WV2jgKgRRKqxNCc6c37/kruBWMMA+mY/5ukLrLp6tjAH
E/IBIV2ZCZs90X3Mk00a2jU3yg9W0jzK5dBhe8s+RgcaK4DOc4z0YfbA/LA0/cFZ7aR3hBP7fLZT
Mtw2HWVPYpia4hObpl2ZkLu1y0kJNIhnr7b3nZgO+pSn5Ni5wQrEHL37NXkoXlbBK0TEEIVkCRho
trLc3wv2PDK+CXHpjYc3ziLTQZ0VcFcJjHb19urFfpxdY4+mSTJI1JBYKvXm9IbXNaU8GtuRlSm3
JGHg2q4fL7C+CFSToavOWiJylSSaJlb5bklSO2zVXbDQJtYghhTvS3cVaaibVci+jqI2PznJnfEm
beORJaLX/WGU9QBins5z7sriXkh1FFUh9QfmZiLslz+pU3yjryhrpVpJ0Q0ZV0xvHsKcdJLO92Jl
UFRqk59TbWx60Dc/+MvESw7hKP+XNbU6IH04QrYL12NCCEhgk8tzzy8nxmE6XTwS+Ea+FdnR8sq0
nZFFGVKDIc9FSTFmJfTo/4e+BvLsKRxK9CnjrREizfUXWMoWqIZIAI4dDTSiVBJbfN9VhXhdSNKS
yuGekqQaeJ5+hs4pGVjLvEBE/SHCMVeGIpgIPBA/8F6x+EeeK2YsS8CADISaP26h6d5yBLN8NaSw
w0R9ixcgtPyZVYnArCW0D9QZQtd/u2g5S+tOwed/DY00hu3iDGQtgNTWOJduyBFbyYkLel0DmAoq
+nEFrJah1jgxK6Rxuxuc25IRm91Li7oOesi4XFdBZkHDTrknbvAk1zfq3m7wFo3yNBA2rJ82pZ4v
xWeWSZdlQgiHVHWhznBiWDXqZDMroJfCL63FkuRUrUKFTaaksdCjXOqOcDFFFv5w07mgbVlLzjbj
R0r98fn5Qi+jNy1o7agCDj5Up8ckSQw765FLu7Tp0PSPLJnhkHQME2OxOfl6uJ1L0BOvBlXnkx05
SuKhvgiG7Ui3ozX0pd1v4FeQkZ5WtXCtWBKDm1AbubnrzjGDElWKgZYr3W/5HHich3pIUMCVl0RX
SUJocTFrYWWhmTWAPPOpac2bh+ZX/gu3kbRxADjPRinrdWmW1djxnLYgNk+cNOcb6/uN2APmlbGQ
cpGP1IxnAGn2JvDp7dFiAg+qA/rOEJcEFTeqbaN5hK9FT5Wqr6CuwS3BIPwM3gARlCwUMkBl8N2W
ckCUWNKDz7fItoyhdXgEGSn5eBK1Rm81Os6/VWq7FT3WpKI3nxAevca2kTgrutecBWKAFk/S77gd
OgqbGTM2WjGIaR5bFLhr2Lgc/hSwfk+1FADElw9kz2nwGOu9KBX62wGAd90Rjz/wZpctAsc/6xEo
Wh0+z7re7GofyRc3A9FqMDoo8hPqcJSWtqKJYR4E6N8NJlHgUvejN9ldXpwRmH7f13EsfDR+q5zS
dDtGA+vk+Yw0/ZHqt2lBBAiDodIkVgd2jVgjvd6fMer2kR35iA6ajbEywtZKDVpWRjGXyrRyI10B
f1lyGHLR1HDfxnnig1bXJCmDlljJi4FVRCDnyOaftF7X0Tue8m8bSTWRtTm5h+eAtCNuxySX7hrB
eTaEY9iUitg5F7hcavG2+9JCBXiNXhw87odAqM4Ip6w82ZXV6HBwTaAdYiTLfiBRLcFu/wVgQccQ
UIu6UxT308xD0KIPubnTEPlmdEp+8UKAdt0tGfneoikjHOnZpRoeK0PAHePAoFW+O6ioCGEroM9y
sf2CvdtGlSoZS71YZF65ISIfbhN+KanoeD09PPErjSX43epNX8VYPst1hFxmQ2xMGIVR6yIXNSmo
u8LDeIT/9wZwF7J0egtXtxWKQZvEKd8NEvoJmsOF1Y9VvNvEX9bG0TrXz5Sn6z5taxMY9vi+Lqn/
5J90Qen8k2adbr46KF4SUxu5kndIx1+lCEQCsBX5S5oUMdzsJsQuWHcGDE3VLh7pSR4Yemm7JCCO
n7L8ZYxWZDPpcT76SKh7G4f3o4EVp3OBek6qaUXg/RiMhq+FLPSvngm12KBQ3JuWVsnX1FWiSbil
faGAZW+XqFKXF8i51OO/UPczOb2QYT5j3uVGGOTzBRSHHrFKJlrlzvuKR7vnlTc2BR/i965I6I9Q
bTcVFZenVSDdufYVtsgLTJ3gnDTCwi2SAIZRLrR3llKxB92Nfi2/ucQNteENKCRt+CpOSeOZDM5L
y1jTne9oOs1J5PrIs+1Hc9qJxTR/wkYfsl6490FPPnZ+ZaqqTjKNMDoiEgs85N5MM1cd+DXU3xQA
P8/gCPAxB9Y5xS2CKg6yR7DF9HsnTj4vP2vWIFYeGkzvJ+GLnXfNpdhDIrXeJAYSAA6J4syTl+hl
YcVGFlMYlM9qUz5urue79sJe2b9WrxL/7sY7AThuZ12mMA9exqIlQcSQxe7AQ1QWmFDmL35N02yv
+9fdLWniVfiEcGGwbTnSigsb7JFDuqnlgtSkU/Oea0XH6NpBDe/tJf7QoJRKZOKMuNCPg2ufjpb7
FKbZ678Cd4sE+N+1RBy9LYx8tmoxVFZBRrWpDnADsiRuVF9Y7PMZPEIPSp/AC8k3X1xLrJIT+8hG
Ut7iSLPOhWiIdtSYcTbzWXky4xEds1/emKH9WOqtDndR2uM6hmQv8EDrFUwP1V7JJXoZsG/pi/wG
IZnuDLGtS239xdp/9CfwCscKwUXpO3GzgRykfeb1mLc9JCn6Dr1l82vxlMlYB7aWULS3s1A67buv
3vXw5QxQUB60MULv+fRzWoU88hbHqX13PdwztV+/MTihM/kX/8dR3QhGPrbn+4TGTVyWgXTNUO2J
b5n0iz5d0oChfwsOn0RF4OY/dFf9STzIm3XS3k7dZF5diNdGAc1cCoAk2fp9qIswAFGbfwiao/l3
bdV5OEQW0LZKtfUCTyQA/FOSJbVdBKPSMHJsulaaKkCec+v4121GpGWgf8O5e3jTiKiIgx0CH9iX
9xwpynMydxgcgbDtcWVCebB56OFfY8jEnWzpQqPcb3fA040bdhIksv3mva+nlY9pfF30bx368mky
ahyvzI3GiYNmQlrpHMmMC8FEfXPN5rBnhfIkk3eTnXtpgRGGwbGeyyuX9aB9A5jklce187U1+JQA
el3S4sXiKeLPJW0qxwkYuhdQGftrArDMXAesZLZVjI7CtLC71nEewml7oqsXJ4Zq8KmfI8t+0dlK
OpaWWFXGIuojwII0LKXdy6ZWccvCHrgJWfkGGdaIX6YE0myujHivscLwoCEO5rDHCoaQFFIO6Hgr
k26ExqCZXv29GW5H2dNGcFIWKE8fI6adyop8oSxOxL54/5Hmu4fuoH/DOPG+uK1Nf43u1g979Qo+
gnoVvy1lzH1EsNQFjq0xOfToyzeVzwXwfxhnIw9pUQUXawbeDG0eV+1xQs0o4Y/URXJxtNuDLJUj
3LnkcyOZsZI1sPwoVF1lfFHtZevtnGwbExpsJy2TpcXUDpwsUt2drh4EeFO3dZcqMcjO70K8xnJ6
m3+Qmx+Q33yVDSLGz9/lXzkSBilvGx+ireBFWJC6IJ+DO0GQ2gFkuezdr09/6NdKy9wIU9rwcvgF
ZnrOUWfdDpbfnvpymIQABd8K1sNLMkG4+Q10Kr+FBbI/+hgnFWSkK939ShA5nfmcH6Uc8MZ+GYNv
y3u7mAT7xi5MO17RELWPAQSQJMGuMQlGGM+fn85tdURAhkGicYGtUrSS9uMEOxLgX24gsrLdu1b6
pIAQoaYSdWKRkI2RbLFYlfmr+sEHC5raofuQGtWG23uYzCaHNMW9/oICY01V3LxQJox3nyVMIgeu
DGeFTM19+qCVqQRGavhTErgNJkwWxDhdqO2Als6HrRH3Ytru1l5Jn8TxBRipjYGWhSPhUOAWxc5b
xIdI/fC4BN0bJY9z4gSCP+5kcX33wMsqPnA98azY8LxW/BTF+9c2kxDQ+K7d/CybCc5bHQkDdE+Y
SuoECWM/m34A6OK1/muIwNzVv1IRV2imebca6vCmzYye6K1uWDVSW2yk8mA0schL2FhvGzA73+BS
1Pi1bUU6dnU0luIdaeI3yE8+wWXfeDh8vKFx+HryWuUGNDgHb4yeTWMiNrHPVeiR4K1GZRBQw3Gt
ynJeWxHKziho9N7M2IzRyff7ZnBgwJktWR2+7RqFUovG/w37sdHMb4vw/RO3/UBNGMjaHWTmOmtZ
5DVLyXjKCoEAwPc9Luyn95qd2CcNK7VTvJ9LSfCp3MJBIEUm7kPxJXzzc6eW9B5APddyoLJUqYWX
AFNTPQ6wYHIzeTllcQU8MMoPS4pN3ubhfTPBuOOnrFOmKwzH0QMyPfGEXpPQfOq5++3g7mSLaCPo
wIYccns9OEovSezGmvOKMDy0NcXCgdcUQiF6DTklWh/dP6l5EdHptLVZMqquC+ukFimCLdRwLSwP
7qblyZEaBKADVXfRG/CdDX41nyM1nN62g/bKrWRRYWFUM1IRp8dgBvb7RiEJGLiYqufgLe+fl86o
PVDD7CIZbd1tXun18apIKH/KutyySGwwRpSKtVwBmpGg0UNrUqCGbG868EBMptwQTvwb9nM9uPPE
36A12Tv7EYSv6e8qsW8zsdlLHYLyAKgC5wy/3xnYgcFV4ODUBjoHue7vhNSx+U5e9dC5GYKqAFSU
dsqzkFZd/Q7uNJQmwy5mjGLIbd9PWcYS8ElaRxHTFXKAeHjW9/bAN9JkR2U4dy7eIkhxh9OvZnP/
pxAal3Lxjseu5ceMPWKRZrRkI1dlqRqSH93BoKFmktrsSPQFIYgefsd1greA9qnKpeUkaZivwjMS
bKuwNkAyyP4eX1FUCiEGbb9jHFT8LUkDArsX0RdwJArx41Xs9XjsXD/AgdwUC1D+zCdaZ70DRcTH
/ztqcTn+3hS8jyAptEIYdUWkeZwqs8fKY6WERBJ/PQh4hnjMJfKHam3wEYK2vr9g3dtWGlE5Enbe
kRi+x5UowZnJo7ExyMrunJaiiilBbgEuFpqUtNan20cwg3E128YnpXk3hqBMgt5fd0dEWbwF426w
QsqMaWOyr3ufhogmv9WggERoDnwev7FbmVh5/B247siNZikllSpaeIvK7tmpX2n3JwL23d/jOT15
qv1xhN7Fo4a9ozyhV+o99jHm235AFBQ/M+MJq4mGVMChlHTh9+iMFh9pstgDbqgRMxmoCP7sLDCt
M6ocI21ekbp/c+Vg3iLhYkkNcDTP13cIq5nglDIIYjlDXIP/sIxUWYmOjVQeT7FC/zIDPm0zq9zO
6dus8WiY0uN2R2B1rqRaZfd3Ybrb1Pe5xIqkfu9MKx46/R2UlAZ5wKZXVmfwkeLRIFprwjzDNNK9
zSYf8xr1n2bjd0HEaJ1yZ240AHbnaJHuTWNx9TEN/LxGl5qPbcij4iBH4cjxmqbLoSvCn0oi9AjZ
c5Bqivluiysc06BFezzOcN/TyksPJHWaSIQ/dRqE5gMlBfFZkv1prz8svL1bFYNLeh4U38truuSn
smaSlk942MDVQOnUH+v8c8u/u65mCRmkzSZO2UTNeW/uJw+sbX/fnEdc/zICYq/zYgJkt9OsiVV/
yRTUNXGQfKoLi1KsjZTor6aOH9ZG3/ER5pz6HAtD1NhnAqOEjMKlw6tdYrzv/+YM1cnQcTW76AuH
ZSCySyAsYvpddXC9I65+Yl0WxcGUJimPPRyQ5si8zU9Y7mRwlmFgndETs6ZK5/FqYwt83zjW9eSA
fFfNWkhVnu4daMXeJyRc/t204aB7HWI99W5NKszHMavB4+dELw767yZpn2nRxj12JdTG5AiweWt8
vlCrjqLBHYmKZHUQUKvJ8NuNVdBY8DBH8JAcKt7zCtYkZbazKUH0o/pBzD1+j6y9B8mYdw4YVzRC
aEgmyHoRJHCYdFB2l9ARKg+fZ5OSuKo3I5zkDRCGbmFdntr5w0fW6ogTVRdUtclV2eWlY0oWo9UV
RmO2FxbVwY+admjSD1bJuaD3WQdcesmdgUfsV13SdT93pYlEKH6ruewrubCihtBAGAArXLfe0JY7
prwYaqfqRfb/SrUWNiTNHfIGliwolSITW2bBp/R4/5wzwBPjqXvWrQYT8TGHYzd2/Pu+S3LafJJl
T5mx7ACs5b2Csc9gXfNzdul1wq9mdDrnArTTIk6SXdO92mDdnebahfELOyf/xp14MuysYO7xCGch
bHsT5BYijrU7Fps6F5DTCRlUIsGH+ZJbW11M64aHNwW/OccBpMOqFg63PNpHt8ZWhRRJallng+UO
R9TsmpibHfaY1eywxYxExz9nBbUxNn2ofbm2mdgTFFSOJi5aqAFnH8xFzoxm/ezNVrA81qQPNXhP
Xhqj3pKKQbpiK+NW5lT3olUgKkLscy8Td49axl6WEj5cW5baI8jqiqjegXWa6BnwV2LulBEC543B
2NgGz6PgFdQngpo94yvVlfWRvr5XvL3Bho1jy7rrOOKj5SWh1AaiQXGgFRJ6hFYvZGcksXKGaWQm
Q1lesaXa2UBk6gKLOWsA7ac1oCS7/juPIcFsUHHq2tC/7PMSPRaOYtA7p5AxMfIREhjOp76oZzRu
C7UJSpWFJTIKWGJM3J0i8agjivEavVM9ig6bOBCVCsiV8gXihiPxd3Yy40EOBuTWeNNFiq8m9Bgn
d17ey08vn0Mtg0T17lEfvNKvWqrL9wPTdxNgC6Q+K5ehSM22o1vzzsZewqmaho83Jl+gZrVbPxbx
gZ+JXWMqhsUzqNp4qiirRMXO+9oaWoeNgd8hSuIyQbHrp+qZ7JlFNiq+XTjmO1FDl51mpgK2ZOa3
sadThJEmUlTtSdk4vIdVl7RMa2bEUXDuo7dA6lbARzma4utH6v+OF1UQmx0N1yyEZ2BPMb9J5bIH
eTXM3IlFhxrSy/2GQLS3WfeVCG8WjfAiaZmoxRGpa2hElt/l4gvzfppBLgGpS8YnDEUKgFuYwByL
bULHHGFzMdCnE2WaX4fdbqpB9BmspkHBfc8ZAzcXGN8ThZ6xFBiipxkMurFTXkYI4KOnzUljcWZz
jQTqOhra6bacqFTd8bTf9YC8ndejVcFH6/GxXpJK3FI4txfIuOOfhMogLSbZXadPX6m0FLbG7xlY
e2AI+Qlf9GBYxD+CXooHJODZ7BxeGcHx2umLf0qZ5c7Ilw/REyAIAGCfR8NJAwPFI5d/rIy3qmJm
Z9+MmnsT44WqmohtFFEg/MuYsinhJhvRgT3nwZVFV4FgCSLFB1q2hFLCdoDnI/JFpD69XEnRIGcE
5xDwC5tQG2bFuv0PLhLWVDQYbLfdlxtfe2mKAXWOaO7O9RhEPuBdbF+G4CUuYVVPBlAymuiQIj7j
aQxKbbrv/Hr3uCjSkccK2MdbT/qkI0sviCsC2Cq7xRQIZsRS6y7WDvZqBZV/abkol75VAtSoSkMl
P4s4OUx8i9ouDLZOtDcXj1DNFHWhdjo5BcIcsU5uq75/YAhhNhgMqLWjDovr56ApMRIm76HcGWdq
TmeQp3U6eJvn6uGRm6sD63uFCKXYklfGD94myfQxf177H3dd43uoJnvTMl4yiouGS2+0K+24XKD0
nVy1Dr9wgLXPvqbNLE449psws4W38zQcxtrlX9GpQWDSxKZTbrY4i0bYSR8iiazK9TGmDMJf9FC2
M/oCGcUNv90Qmbca4dMr4q6JRkAhrKQ4zFXekSXSMbhcIccREk0rV2ylMugNJI8wXH0U6yIWgVVS
3UBXyOWcX6xJqoFCWzlrgEg0wpn3OlG9Hk8SdljE3mQiGQ+73UhXw8qnY9HZ9/Hb15FyIO9SMKSC
3cK+FKEnBVRQRzA/V4cdUXAt8Ir1GS2jNR13Qya3d9FJnK4hxRRvumfEwOsO9hiutCW1a0nu5XD9
2J9LEbuJfuO86nFtJoW5BuiObJC76HDcfSDE8su/1VRlhIE4ZuOGi8VCsFh/Inv9FBexfFeVy0oQ
9kwN5zVxhCbx/58F6BwP9yYi/5Tpl1TlBHVvJuNpH2zE1lOvfziV5BGtHgh2M6QlVIcC5oBBkPXT
F51skt9xjMa/6lmJSIvAdaJqGfeXQRGVAymS82oBi9dtS0FWDWHkBIdC6oBwzrR3PZt3NHo0nCgb
jtCrFm4Mwo0JUCmCIwZDtz8HI6Q4y8kLIZad/JCQAeJ1i87m49Mq+weyzc8v/icX1JSycNMpzbWA
ynnQGA3DeuS/u/RizJGktHZsh6J7iAf3A8G4Xt6pNmw1MabxmeCbgREDO3oHgnLEHzzyUrrn93HZ
bBZX1B9T+Ge7ykfC8YCijXx16xhn3JUx5RulyGvlSPwqoN+ba/UdzTL315I+ZWkOjvWsTCz2W/0f
QkXnp+HbXnvNcNPTVo9xiVkQaisFgAuBqi5loKzRC1cG1HP1V0yqWTC4DfEhNmsvrZG0IZjBG2Xb
f2gnzUdilphhocvBkNAgihdzRzIp7B+cafd4l0qhEjOtuiLf8fJKrsy7x0rMKczb95dCMn2SMNpi
R+q06h6NovqPr0aWUMBrizaXpdFd1Wg2x1vegDZJ6vIOTnaROjaVrJt7hw3ywPbWTQDHmZgz9lGr
UmcUPIRz7rurryqFYAMjPgzw3jhrfUMzbIxoDfwl5W9tGBsKdxDdDIxE5PFjCBUxSlV7riH4IiZX
MEoi5BqAEl6vJM7MzTvUX5MGNc+l/8teKGh+aF2A8+dJ2m5TNbR78N2Nr+F+hn/r3p1Yg7Os3MxB
9UZZceeUhjZ3QuBYNdHDAFD50e19LGuxl5USzDRRoXKTGyoR9hSEhtFilxZgHTMRNpUYXHLqdkAo
2N5eyRETDlEbj+p7bYqPsYNDYxnzRgh7NllT6bHGzVv0ZZUARryhjOlhS9OYEWrTmB7WJsROXwdL
uiUt5+mY/qCYPDbVzmluOg8d0SkehTp9lzF53skZ+LAh7EQ7XAwUBqPT8ioy7VNAOA4GsZHG4IEP
dEZ3D6+l9yCWNKxy7BEBRSX7Q6AHR7ewGzBqKzS6NIzUMDOjEzKyHrdw21smH7H0cDjxW1/gr8x8
vScmfFJG4XV/P3ifGVj6xBTOb9jVxcyrfHk9h8wh7hUDthaoV1QpoL34mbVlEM4snHfKJWpjWb9i
nv7oNQnQ+wtbtYtHPUbE70SJIquZxisUOeEflCDShlHpE78LNcQbCv9lB0mSsbKBHy+7Pnt3L5rn
HmAh9UjP9rAlOy7w1/0yOzI7301HstKdCuWyt5AQAOqTM973F+3y66lvOUAfO6IGwnzS2B/EOfSA
LtBKtDIWR6Hod3Gwom76b4vgSHGwrttadnbYHBoWCmtPA9wOj+XafXRAT0lJ1Rd7q1eX/3vF6dot
4yc+nA8W2OU3mwPU4zkAiuaJL41VSSMCqUvmvCejdUzt8mY8mbCQm7+IVgr3GoLKZHWFfEK/iAHa
AgjSw2QOWagZhMAR5xQg3anfZiC8YSAbZTREeBjou2spnCRbHcvp/7U+y/p55Qc1G28Xev4Hrp/+
EkF60WCwVOB0qBQMPdRbEDufA44EhEOvrKK+mRMumvADmMTiHIBwC42YSk8UPGXB73M+EnpC4iKG
rE889sjp5hiIq7iZ5xwmQ+Ref1RSKA3REGzU6SEazdv32tGc9ATu1Zewd4sY5qDI/oi9q46Ukxbf
hor3jSeDw74f+kSYmj7fCXuD1VfURmr0eOb/h/ZqqJNT8e9M4gF2/nnvqZ5y05UuD1B64KHio686
G949K6H4VQYJmEcu7PjnOCBLff6MyQCcgYVwaN8iDuFDnIEikf6achjWq99v1baAA99KYGZyxjcs
ne/gpf2M+byIXwy82+SxR8OSrlLRNKjL/OKR9EKJNy1ue1gx//bOi/dOe5lxqXxa0kjnrJdU2Wfv
5YUZiTnuOlH4ExKbl6IQuVRzt3ez2o5+oRdw4EVRAfZZilVBdb5z3KAaFIKPVywzdLjx5lqiBNWV
mKBuZWtp14yA7Bbo+ZhRD8veBDa4nxFFpW/XD+zzpa7ORJIN1wG1v1spoI4h3TqnA7J/KMmm8voL
/Dlinorrjhke8BPsZLL345zUKgdEpvCwtJl0QFk1ltHTrc4Rcub1EANN7AZOlb4bk/cUYHy+Fve8
vblbmvitzWck7qNP4pW+kY2+RR81jX4/7KpVV484VVS7ukzTvXsvOrl0K5+eZr8rujdiWg8evzx/
W+M6unuRhg0oR5OF3psZ7P+DxDJM/j08ib/haPIUpF7vNXBr4tnG2tI/r2Hz535v8I61qkiFALy8
Tv9gPPTQugd5YLfN+H3j2Q8A3EgvQKY6U7PzCGQk5ompEwtg0BllLr/rKmfOPP0RJVXPp21cdUnS
fnurFxQWrqAQr4HvjOv1ZwMcXudCGwssku4=
`pragma protect end_protected
