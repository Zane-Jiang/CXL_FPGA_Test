// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
EwIrtyuoxnoTyZC3KSZ/Zd5HuDp40v9rz4ROZx6OyWzMADMYALTF3bPjvzMCynI1
xJsFg+AJidWwZJ5eBxI3qMsrl0zln36Jd9ZhEzTd6T81hWtOwtoQCSO29Ob6KXqi
tPN1AvlOnWC3fWpjneSr5cEjmnrFKs7PpVzOQUDN6b4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 217824 )
`pragma protect data_block
XAWXMJpz7146ePK+6iYyaekUqiexXaObKY/NXP6MR2TWIKgUugO71byxYeMBYvzq
Oe3I8OHcEMidtstG7cqOpqAmrAjUUdL7Bq0b5+3d2r/4Wz9CkmtQq4DhsrGrFUgl
oOUR4YCpxMbamzI6wAfwHZKHywPgWS8JrFuu0WlmykVsFRYQllUTTsOITuK6Y2F5
XT+o+zT1KP0PGRw4xXxfZ8tFhwGvwPvzir79+TuWIXAXJ6rwpNGvAnvPlua+Fou4
3oAp42QPLbyYO7Gq3Wqd46aaHSIXy0qGVfc5iZo5O8bwdNEWm0db1Jjrgl/WUfeJ
QPPO2uIBqL3Li0ipGVVgJblO8GnWA7dGMjhvNWo0mBKvEgXNBiJLmmw9ZGfHKQnC
ThfJe1xGgbCUqUwDQxqvOKxkEy8Dr3NEB2vw3p76DoHIVeUdotZXKef8bOFkK39f
IhNk3r0o+qi2r6YzGHQG+/PTxIjhP749XK1WQBqOncnoRFMc+D5qkghOkAnkgaFp
qzImzv2BoAr6cLPwa2cTipcxSs1XuFrhhR8SIVFfRfGHY3d5+b6gXg3sdrZzdFNa
gtzkMxx1ymIrMnarw0xlochxn62FlHNTnQSNllehizi7qhppmSyGwJg2tiokV0D2
hX1VoE/OQ8NneXiD7O91PMKXlnMluxZXKNnkVU9kUUFW7Og4G8CDx1u8f7xrH+ly
dZsZMo7h6ExS+50a/ypFrNQcugfXUMT4+Lul7/UZtXLt6AKE96iNUnD1xQ20ykm4
cOB+gTD+sMLzbJrjtfNqIYSXmvROhc2npLcrDHWkOb/GhtnW8lJ9pqp6AwKHQCkH
oJ/8Swc2biXvYYF+YU+rJTQzHM83MovCLWC6a87CS7nTCZp63Fi2GuQQ11RTPSri
/mdnDUPHMoPizGKOzOB81MrDjFObvSX2YkUra8D4UXZkJpwX4rujmM7L72ljGMZt
1+Qv9LSekYgwIbYpxg3lmAWGbpgRy0OBXLRpscPQuv5IjWNDjCuw2h1A+5rAxcTr
CbpDDDXIvxtR7g8Snr2tt0nKjSwm099DX15gzTJfXQia8ZM8XGJC4vj5myDPD5je
nxNwLftBI2aTx8MFq1hRK6YC5l5hohJX4eBewvH8wxmPdSttExam51J4hPSrdYo4
iV07WUcLpYYFoYpr9WDF2KTImT6CRXF0S2T6bMeiIlhkidMNXoBIGnic9Y8Dxm5h
6fuv/cyTgaS7hAJhtKrKuNDTwnWGzks/Wl4s080NHTFRneLUMLspuf7bxe6KpCNl
9jUylLQXrHETCuQUWRpzy5AXycak0okVIjUFScdpnZeq9hE5SlutwpuNBOOfDXkc
LbvluB4flDekFwJfPVUM1BA4q4NX0yBuN19ngV7Vwj4bRy6R3ztpjLmZyRTJLmPM
HvggVW4X711EQKfzUbRvVGU6e/tc4MbmiNdExW3mBQ7UIpruJdKzELFMMY8olZwP
5mmipZt53u1IJmAIQpUxn2TPfjGHp6ASqOhgkwyEGrI1TUAwgbhfhg6mlGHPwz4z
kVlEVuYOKrEDNoHeiNNuRxcLHA1r4utcQv5Wko4RELrt+1y7qBuuWMXe+BaMSxwj
5lvOQebrEym5yiRJ45KJdpow/0o0MzgKg2t16OVDrY31kMyrioaFhS62GegfPOe2
vj2LaMI6VDt+pNKmdG+pjs5imGqy6htyxkR3Jjb0LkuxL5k70ul6sKZaqaZrnR5X
cfaGQegx8u9ZqTdkKXZb+8HmyXMRi9+rqmwk1s8E+zSHr1MXFZTjzOvs4qAykXV3
CNeLpU/Y4bbCUGpt8R5EVA9zsHil1sPx+YDmESRzs4zQ45k0VJsqeAYZ1GeYdrcG
t4mqfmHxqABSLijiNM3RNG8jZVgyO64bVl3ssuaBJ6pn6Wg7FSspvlUgMlKWWdZx
mE1dQqxWtAw2oM8ECwfgr/Ddlyx7WUc1lYVMUkTIwCcLbY4yS/mfo+M+osUqJ7Uu
1fUNcJWQMQL3IfPtllgBr9pjkGkeiDj6gBeQALNXLH0Z21p2h3FqMF9xSvV6BxrL
pTty6/mWJDzi+bn6oWLHSwgBlzjMB751XVwJPriTb90gCjCw/S7KPSYdKx51FK2Y
dzOkJXcvnO6xxB1nkX9lNQBQFcxJVNyRbsAKSptKd6O+FXMGMhI6ulw+5YdL3vYB
KMYQngFIL4hWEfc736UsS1wM04iEGjatzG6gFAUWdxnRQANvPstCcdBiNoW/wH1H
JMDsUtZcQCi0s+IpxwMLCX53bPBsxmuwwjsJlOshMnzqU3Mm0NHbt9iGibdXRSiy
UFkXm+3kG2jyLL1YNxorbjgWDBMK+NDLBeUsQ3HIGst8Zg0/Stpx3LHRq87PE3EE
zNrwVfWNbx7A4v+eWGul6xNlosiHW10x6tLpBnnubBZyhVJxeN2nsuProyUjg+vo
xoR4I5PUwlp84YkIKxvlpOgxupyO2zNjqgrkpNsPAgzbVTdiOV+M0xlqSnyy1EC2
EO+9/2BU2DcuOBycpXUZU+DB/ubvPUcMGObKdSTfTy0se19afZaFBXlNZ1Y+g5Ks
mpR0cWccAyF6Ct5QlfC1sDuKZ+S/rqgXkxzoGbxFZaVHdiIQwkg71unqaHvPUBkv
btvrZweJxGMIZX6FNtKaiCQV0UXarOguf8TSJW2uOeBVUuYwGzP/F7crJc1WF51s
++CZRK7bnG2ptTJighMItw8cZwW5jE2ldSlkp840GBZeel7aMFCUkusjmsWEYU9W
F956UklRhtHx4tX7VZ1+5ni/6onFd+Z1XPQJWa3GAJCQWuYM8vD7Y7wGF0LoiPcP
xHUnZANZZJpvtvgpOec5xE6vNLJTGvDlDAsrZ2MGqjvD7wopGdDFs/8/iHj42HXk
F3UFBWsiAQ0qm4oaTex/FuXtBrn5Lz964E/WSp015Gw1p7MApe/jjGNOswFKhb0N
ttbQl6Lg0zhr0WceiSt3MklyZ5YwZKwgOcph9R9g9buNLON0+uNh8A+9jzsHX4EI
BQEs6x0ck2f3UG8WxdhC9LS8ML9luUN8mFEAQY+NpDb7UYsxUxL8KMfqDWY+Kdso
W1AZ1M+GYoZAeRhVAYDxNlXdv9XKHgZMoQAKf9s+lvZ8ejZK6i9YHFNEc+fpKpbP
O/9DgXzP8Mcvxmqbis1RCiwJ0VI3cFPjl3MPVNyggVcPhB8P0h2lH6E2/yxxuPr7
GCY+BPb6+ypfqNeZYuAkjIwJGyWAsArPzrrQ9i6QdP5rDqp9JdVQoeNOUKAbPukf
TEjPe+rF18bHKapUKi1KynJVcM7j0qlkFTxGaVmLit6QyI5dz84Zp4GTgSbmsuVC
0ZlkSkETp4jj1DKEfaDCzLvUvtK3UIKevaxIiGgV9j0oEMxgr8kj/9hC/hnCuQyk
ZCmGKAH4aJdjxIq4sZOscG5BPbhDXsGPQN8HxzmwgFG0ndHvZFMeG5Jt9yYVShK7
jVlwcSdH0TPZfQfE1jeaaBtKMZOn3m6ZXK+FnqMt6BF3/4wvrtCm3XNJ5kl2GvSJ
Gs0OB08cWJT8bSGVNpFY3xFDRXfPX2qDI1nr1q6wqRYuL52pFI9s7vJDC/NmwAL9
L/pjiwuxm0xgf/MB16dcB717x/eNjuFhXxca6rA8M9yZrk24j+SW+16B+xyExSyW
q5XYHp5oM2PgaeS3UYVCzB7Eg8XWuEG8ddX4R1kYWoXfuS7dXpZdzzcaAEGp1/PM
CG4/QAf3wsBA1Tqjv3Uo8EKMJxJJkKf9VL7eOs4LtKESXbTUQeycucUhyH78WNoh
G5s2H3+IUMd8CTbwjX6Vr1O873Q/Kh9LSKN3jag1GBE0hqUzuu6pam1VsdgvRqsP
u7gR0FoIelbPL7l9reIGNGEbdsqkjkgiSk2XT08zWCvGGqlPQjrfSLVv2noZQ7O+
n4OW8m/DKIAYu4ySItTg8Lhef2kROZaC3nuJZaZfrXvYxnhKpUpgUq9IVnfCn4TP
0x43cVYCWyDMF/WMHVFE3gnV3qUX27KDowKvxAEY8q2gx4t8hSroxiRgBMWRQ3vl
ZZ206KIfWyyQ/Tjc7H/+r9ax0OiRPUjx/I0gsY7LBdArmR8rtUVWCCRDoRBLcWza
wQKGUGZE7S95VSdM5S44/2zzQ669NtCjgXHmINJk69q+zrR4cEQ8cASYi5djkqBp
xHjAB6dXJ76pHLMztl4huT/jEmbjZCdBCIqvwp7ro5wMVNxw1ay/qxhYWA7GM3Tb
r79rQ21r+jUttQ0OZ/k/MzpcMMTir+r6nf0nzP3hd7v9FNzL40rIUJSfKc9RGemU
ClBAaLhii9xKtPV3mcYeiZWbVkUeUjwzwqrm4unvH9qTZmQsAu3FUOqeJPclq4PB
45dxRPmKqxLUAQ7ntIPqM+z/PK+QdC/wCevyVk4gHHbk4ega8kJvESX31jeVWwK0
jc7I0UQoNG9jUbcFfYmP49JHVT620rlZXfAbVFpvxuow96Pmx3OoYBWO24Heslwq
amO1XPwknPzPuxpIQ7Bh3zRZY5aDhydCl63owhCFcxJRflGCywpw5MR/w6JxsQy4
tvFT6VNUgY38wmhgKOUkZZq4dpupMX0/b9pdepWSEwx9lVrB/Z07+9UXgny32DK/
RyKUGMfU/xVzMi7PLPYiwml2y//PbJ802qpzKq/YMM/hmSs1o5nZ/0aFIlhN+F6A
iZoZ00kgpeMmbPcxcZvvbhJYWDsG5xYkHOKxxHvb0qW64hUv+pFwOWooOsBbdvKa
3+BcNEAK9b1H5/Uzf2cia6/KOexlFWZ/4DvEzpN4Y960cRzmmEgKMHobj4p3vOkF
3ygidCaxIc0DnFymYCJnV1GN2kWklzE3SLJ5TbpITxl+L0Wf1jMJ8D8DyBpptMr7
Z9GwS9WaMuKaFqS2PpZvAQLchY2uvaFYaqDj3f/4kLxIInfR8307OqHywPOEcC/t
56g+zowP1EhqIRf2stKmwnaXKm+uGg107l/sTDXVlD41SfbwvttsyE8jVSlugMlQ
VJ5/TDpp1DnF0oHXCbQ5GhEeL9mM7BU+9ZeystLGXCjBaPROqONHtAZ7NtrwHcmy
YyOsCYrkmZS1xq2A6pi6hLw6MZ9EcMKl8JQDNMuWE9e6cbbzbSGb2JxyJ0SJfZQ2
zCtGcm8P+dKbTWQ7f/w47zgmHJic3Uhb9LpMwDZi7EhRw1v2/uChQgoXEi0IabGa
v/G4WdC/ftwN2rYUbRr1p7qyL6hYfvPzf7feAM8xXnQEdL9+TiajnGTgVtBvjaEc
4jpfWz6AUFHBxQq3fsuSjPLTL25FCGiQH/kzRErgd/KE2Uwhwi3OD+gc9MmYwszo
2I2CAWB97480t2t7M2iJ6l06uqHSNhJCO9dDJdmV6YGHjXe5FC8t1Lgn7o23LPfs
NdcTuArfbr8q4KCvXVwpRHa0yRjVuRzUYpPG7Hu8vU9ct7B/iqYKkHR1Deryh/Zh
6Lr+VB5pkKaNZ61MG5N/nqgyzsvzHA/pp+ylQGpJlsmXc36CH93kQh9AQTGGRPtX
Bl6b+ygK8tx1jE7pHEJlQ9Xnu7D4SL1rfDIG62JkhQchRbmSrrB5L6CuXW4ByAqS
GEOaoXlPuSQTQhzeCCwGzAh2H3vKziVropAP28Vmw+nd01DrmLRTZkneTSuBD21+
kM7rlGYTSc3QIMR4cG0Yh9USg3YUzq45ydTzVYVGZcuJzlZLyGHIqUgWqz3bZwr0
38ZLdYyyC4PBxq0g78wDcdrYqg+VN+f+6Nbp8LqJqUmLGA870HaDwk5R0JyX5Xrh
khPab4jaYz1uhPeCwGhQjJP//cg6VyH6a0+s1UMz//fsxm0/nuL0OK7+24zbhLch
8tyGiQg5pnJdapIX7zv1673ZyMVEXqZ3GEsssZnGK3lBvr/aPX/TmQa0L0rXhwKS
OecU+iO/MEHu/dIFIo15BZJI5wWuTyJUVv1BHhhuDXAiFYbD1rh1SpkeY2C00YES
PjNBFmfZtntjHDmJcoIRBTWbzlY0wx1KZ3uA0MGHd6JddE25zGsag8rf7XFVHWMB
2bVfy9IEbi9FXMelEryMejEyyIu+HGOHRfh3caDtlQH/Xb+YCGYalTKyqVCMhTgI
nF/u4bjFo/QAzHQmKSb16q6dhMbtxzC2V631dAB8M//3LvyFo3R+dJDp0jU/4TJv
DARd/053GzwYt0ROpOvPKUNpUey0kfb/Np9c+O27BTFpjDwG8y5GlZEA2jVqASOK
VAA1xtkChlMHRIUCGqdkYZAH/03mb8AfLYWuJ13C7ClsgaQFwpH7WNK/JGpMkz5h
ow/vummdGpdLjxYKHZ8R8HtTpWesXtr1E8YHmihzhxVGeqdqMz0U6UT+1RZF+O6n
vdutkI7XXKydsrV1DWt6WuTR/OLTJQU4z++k33clthEHijWgWSI9Cuq1SXndlbAY
EHbKR3a3yhzrep01jgCPRZVlkazCUvpXWMffyfOxopLWqHeeodlOYpEREryn3Q7/
dzBHCERwgHoEJBDUCuoRKo2rogybXg1ujg0FGpdX0h9mnM4vtpSFN3QET/xh2kvj
GFAFRi+QkbUGOQI2liBE7HmDxkffZ2gIFlqPla3yZ8HtyLJDspWE6ToRimoqBUjg
GI4kqmOP2KA3my6k86ttl8Dnc/nP/PO+HgPBBpvAsSRO7z/Ys8BEjJm0VgAED20+
ZXL7tWa+nBgH5sAlEqPz7gPu5QG4DUYeg8/aoPg/pDTPCi30mNNNO1wCzko6acbv
b3HmpgV6KD9WiDzWwxoE276KbLiy1JHtrNVCsUSOKsOjVR+qjWl8A3i9c15jPf6d
4koYLKN3hRq5f6sb3t1n87WSvZZD/2Un0U8w7b+y5GW6bYEvFs3OLyRFsalKx9VB
29Ae4nsXnVgWosn8IoB6kBSh/qDmChpNlGcsWXcjWIMyOVWBMPutF+aIL2bMYYrF
aaV1M0yOQAlfReR+Sg/OXNDx2x7bex5drNQnoKzgg9JEALQ2V9UCdaRb67rnWAOu
rg+RnRXDxA4KX6T3bdcdl0VZGMJaclnr5+frajTvNNqX6B/66Fu49aiKkrjd1RIt
sZSyeUbf3/1JwUaSIerJ60sAndcQO5ULV7baOzc2iCuwL+ZLto25d8/MJm/WKflh
KHm/3Qogu2/+WMT6yM43lZw4fmVZXBaRqp6Ev4j+ahEke+MOTHuwmsS7OFR9OkMC
157QfB+u9wkX0ZscDxMeio9UP8o/0vK52WljnSa8b4D8H3uW6FAokZ6tj7jbbV2b
K16McXzJRLLryUlNyXPKhFLsdJPI2Rb2kjfsUbYjbcN+zlnTQsZ1tLhCoPc5cM9f
22DJHz77ZGp9qEvDNf0ZVBQ5uCcd/blXxgF4nkcKc+h/iqtuj5mxxfMRg7DoTH0C
F4RAoFiaQPviiEdWqVHXA0bLtcIYPl6GKgMSFgFv3JVEllQHx84pJ+hU1JRavF/3
zRXuPKHt5riW4ZuUnycDSjTKMnOQnkkjWYrhFDVoEIS9sHH+xGfdqrkSbGFEIKGG
P4yXNgmIndJJyGlCaOynOw2WUU5eVYf+yJH0giYW6Yah+J9O9D84PhsXLvXr1r4b
qZjr+nTSg05wWCdZ/VWaHIwnfFbPfoeMyos3v6BEw0pw8svZ+1AkMueHb3J6+id/
gYbmcAGsdsd9+69Z+qYt3Z+uzeOXu+R3PFrDAUBqzaeK4pwabhrZplSU3ihMBkC/
I0z1LxATtlOGBM0GlVFtK1ya4jGfGxDBemIOF0kffms0Afp5FLUJW/bWyFVVZymi
rEK8YRVh3cXfTvzTANzJVO29MOiQJwDeXakbXa5cxp78PIGCAppYFfygzVjUa380
EPscGwTaUkY8EOnqniIa5At7FK+aU6kbkynF7O0IBgyy4HarhUCvB+kRAxIT3fpx
+xsrLklqCLZjZ1hWoUjt3hO5DYhegpxWreXLb+gIXBCSkr7RSc5TcdkB2R29OBaK
1PO9T4Kht4ZvSnhb4lozgHhfHw2L7UW7rz3qMTu7HFuZSu2okMh9BHfnZLR5gWQ2
CmmufBjfPmX3u174lugwVB3limCZpE0oFpXDqlONWQ80/6eBfnQzfhSE+3YBKoWs
G3j5hX5xoMYT5Gc/YtulidhomGV1XQ9OV+s3+Ra35lOuobdp/Ux8JHrWShojjHu1
vyf2qAh6k+fG4iz4jdEN7LfYw78I6dJVZ/txlS+f8SOgkJiErzxlN+5ZzoRLD416
Kf7dTuNNPBZVbLtCASQ7LHZKd6NhpYuCfCGSt9TAemfg/FTrYMJzW9ptvFLkz01+
myic8Qa+IM8aSCiWJiJbeiCtEq1Em3uMU3v56S6dlyr72PFpvFujF0B0O8wKWImw
N5sAQ/g7MT07rHz4424D6cryDMo2xuxXR7Q0UUObs6JHu2Xq84TeoyWqxU5+SZeo
uD6hmrFM55HpwC4ple/CyWtraupTAXARyQ/M0qgeNIOTo/pwf5Gj7sKMEEYEmv6q
B25fwWJIiAQsAQ1oZ09YUYF+j5jJN6nkPI6TqVOHpp6WMrWRAwzMp7VHG8Z71KaZ
L4NXcFFUK8QnIHdL5sgkO+8Z6bHz/bekrg+hVTiAGlI7g/dvw7RdgU8LTJH3r1sy
3e12WPyTmuyg/y4sA7NsZElKCiLQ1B5dCdrXow8xNYrIoPtyeVyWjJ7qB+HSZnN9
eKJKpt3mx+bCeP4UGgb8FGvkZ/9QI+ZCFi+E8Xmten+y80B/XymWP32xUpHBacpI
HxORkGWZcvV/r+n3OLw75wfUT2HdbPpBux0B7iwwt4jHoev3iBoh+nIH8u+HKOFd
baj+NMjBvME5/lCZTM+RVNx9P4c2MBqB/KORFxIlftpml8no0T/+v0LzjynmYJKh
NaTTfijdGVtOHxrmk1WbGxAXrowyOcNnqdFP5NudNpSHbMHNjxat6c3oRTvg9GSM
X+ExQWDkTVn1YHiKr7ZeYHpGtrXlt6rFwCVdktsb9y7TiF+lLTIEr6YigwNQ5/XN
6WBz4kQEEk+f5h33if/OAdChypxcCGPSwV/KwDvutQ+mZe63pAGh1ZdM7DlI6Wr/
Vz7KTnnKBzKyML9sEZOEELUhQyazf6x6aIxZ7hwTC0Iv5UwgH0TOftbt8Zz7iHZD
Q3kQe5bilzukjVrlbtlZezyCY2OhZE9eCRj201ZpPfAVMOycNbZKp5ZZ8ziSTTy7
TNPz5XgVfwCq1j48PBR+H+rYXhpDrDCS/sEz3vfYB+y10YrWfI8Vk8Tr2vwmfouN
1yEsk0namehXnMz28dlbCkrHPatb40j7zbhHtjvw/D/4myKOzo433nDIBzoJgslY
npev5WxDNfYtmEdThb5Ns4XqPNPBPzjMGvgtVfKglypGRsboSgbLtHdKSMdBsotj
519j4gIxHkKDlSGe0/0CyjPeW/KnYq8Q6Euy8sC3ACZuWyk4RIskrVdA86x3XWU0
aIhMfHobzAgZb3bc7a/BXJhFWnQibxpPodKN/z3pLl8WE4f6vZPPk6x1zxNTEIQw
zJ5semawpbW1L70SZNbLx6jWH00fI/RuG7WBEBrKntATBNqechfe7sLVYH+0UmQ2
zZJWiEM2kK0QbVw6ewtNHodPESg48Fezq0hizMas7RxveLw4Jrw6bub0DCY4XySH
PzNCMFoPbveD3QWZpArumKZbCryiRm/rn1fFJxXBK4U3uTy4570kbc3FMe3g8XWr
IOM2BVfNQT1/Xf265Xv3HlWPlD6alNjbWuYX3IMf16UfwGR7JJ9x6wrqc5Tv9Qik
ryWFXhzOaN2YscJpoLxu2Oa1jVOVZPOU+O2ZlU2OmPvnM91YUA/eFoQliO3wGAqE
sxGGrApQienPNi3uP3NmSmraf4egQRGRPNcwRUrMID2jgf3AMvarVMhDbFhW754d
iDEoFzVLkhdJIBw8pPsQSPq5X5JRubVRa3wvCPfWhIx6E5G5X+YT9U3gkJX37dqP
ZCy/UkiiWUXHYcwI9dANC6hb7strg3QtcxZfMsqXnegDS6Dihl5EVer+5awlrACG
kN8BIUrkQ2f2SbB6eFdxjOn0eW7ItqRZeyB+Dj46S/KczzYaHY1qYEe01amCNJBr
LnHXiF452iUM14QlyZNd5TeE1j2A1QejUPj6wJQEoX8RJj3wjFxm1BSrdGNqHZDW
zvw05KofPyB7dJTlERJsxPRhUEjvNlcjrsvEMBZE2Wpwaw6c9GduYPfFBEe83hyf
XKSqZMzJYkYu87I5YMnZQw8jIdl+2VIsiPXH/0uh2eDYXyMwI+y1GhT+a8iCRnM+
JgKjNfrWZ6P4iuibzxcz1K/Kom/ClurtVB5XMH7ON+gdOELxUzAo2wkNAm+FUr/+
Tf3TBMspObuJ3XLL0REhFcHhsaVmgumrN989NG+x5tPiOgcKtumtUjCc8FDLX5YB
yiSqitqtBIoO+TO+aM442V6lC8TQzPC12OttFl7rRe/3ZRqH6t1ZVmu+PDLvAkSi
7tuDUzFhryvUo+yZjRqnQhTvflJgqiqoNwMAvDdiGE2Kdwfd2S9CSmSSCjCYHCJY
t0dmwrdiwdSZdcyqmzKIoeRWMCdYJKEXQ2GXry9qO5+T5HzALrdhOMK7wyPHYQ7/
GJ1G8IJyILmCORYSIM4Qg86PMj9hp0sSSZBfOvpTiZ2feChxmOM15f8WTS5njlwb
XPYXZ5Z1iS3aXiy+lJQKuIgCKBBQQMhx728talK9lXoZN1kep1RFFudLi2GQ8hHb
C2Lqo5/n5O+iqq2lg3TfwOsoELyarbSuMyfxLI29KDpKDXYIxMebCSkQ6UzyMq6f
CoTXwSdJffK7YCu01Dp49yoM5KgpO9TD+z2eYvjRvEGWVYNefdDg70mmmQ9Bk5n5
qbOmIutjTwpUhN6S2Mzt4c3sCsazAE+B82C6qIRV9FO14RPrJn/+WgmKuRI2bG7o
Pyr5yk+iAFiigv2Sb31dbdeasKbpgyzevzmJp9eScRPC32vJdGqsbG7cxq9Hzpxc
nDILBjq2K3Op/UdWQnpHM/1v7fl6eaB8DiRiPVkGGxUIfRzXVx6MN9Jb33Tgde23
K8f0j7i3zOEoDYQeS1RLK/lZOF0xiyQxL4IswBYlS1eWhlIjyRUnGKYyACBgSUsx
J76P70QzKo0an1d5hnSJN/tL+QxKPTWABVmbDTnHGRAsREatNGis8NAjS2dse4PQ
F3A7hUTyx+d6HfKd/5s/tFNVuP7WlYRoMY64YbthbGYXSMVHqzvdYNt97v+kh0Cj
Sp1UHhF4FpP+6xe4JpFMtivvt/KWTQACejRQD2/jKv9+2Fnyh8lnuLbi7ijv2yXC
+Pv9RL0BxZILsukOdjdzRP7IiZX9iNfoUM788VWxW7ViHq6r5wMINJZmvbjvks8Z
lMrRyUW5Wptb6IJOTnR9J6BF5NukGJ5XmJyJhfIvpJPS/e065NKlA/zypmOL62ae
MfzrRiBJ6G0c1eCedNDcCN8hj1wTc/vq247OOd4iEzzLAuG8/NjrEscRLHEa7xqA
t0RBJvM2LthHBo7DXGlDG2mImjoycXMBTd1txAR5doTKX9jS6fA5izsk0Qg7VMae
ogVRipXehEkV6xBpDEW6+xH+5e/2b7GtgWiNKQQH5FANqu388SUeBz5aaj9nlBl8
fvVuikF4iWD3xI5P25Ro7EGY5DH32k8E1Ti1akJiiwl+rxJoW2qmDkHBUYSej6jO
MBpD6xSy18twZMxkTts91/85GHJAYA5fxl7HL151Jw718uafimO1ddDcLyLI8Lgs
EG/bEfuHuMQ+bt1IktQgw9wzPI3Wn5e3YpcevXtHu9xploDwtPsqu7mI164/uTHX
vKbjtOUd2705kHSDH/Pu9h6ghH3URZ7pgoLwnx089vCEn5lBpOMhSs48b7atcWjO
8buWDoN36Xgj6UAysNWJbYbcL8r8MdH9bW5h/9Nmrqv2TZFIJyMfgHiz4nBIQmiY
M2E32Pg14fHUfEI4P35j87waaOBbEnlBxskCpMlug3UsShTuaKu8ciV+piTAPNrU
4QU8pj7hlqVAy1Kzcpz1vhGdnnt5FTCvhT7CGcbsORcIHuBtOCSdLlWNUEztcLPN
ym2XiCEvh09sBGtCyUtPkMfZQGGYFHzmMyO0wFWgXaqjDcjGGBaYKHjaJzeEAjpt
E6nlGmoAr1n/nggNmwBQhyQnC/63TQogO+ODUUigiscYQXHAhqFr6kyE277N0a+l
qjPAshcnD4cjPJ9wYEDVX0LDKH5t1ypspfyJvhx550TWKK9c8mdCiHy5Pxm77Qcp
/2B3axN5iZGajeu6FX3J3nNbVXClql9q4ec7nDuHqgqILRX1xl4vP0DwrOmUC8cL
tzBr7NGiSEgJAzfLl8b0GERPFCn1N/XoNanzMcEc8YiTEAQTwvJ2MciCmsUuqlFj
eg6hGWkLoej0YWpIcyqvpPut/WcDR0Tj5dGEsWPZe0GTpRKeQ16djojLamrLKP9c
lILEK1zuiUZLA6bhhFkAxcTaB4ZOawVMxb3YI/Vpn8pXzg/MddY6XgZUavF5/RW1
490GdXD+Yv1pf+8i1E3+fMyRcjfod869+UTW/vnY0myE5U8RsWqv5kZsOpxBBYC7
EHs1UD5Ozntru28L4czpCHvERGGzKelO2QWcXdhN/jFXuNfW6vhp5oI1p0h/H6rP
VM2R6JqAqluxEEWvHq2wMjFmb5NvTb/wIcGYtSXaWLDTyYgpx7GBCvXm2LYLXDei
DIKN/sjTI4a/UHoG4cyKq0gDcM0qKhIRQfVl0jJsXReW+rEAlCwWI9s1XfBg67fR
RlTtLxjT0W9D03u+QdNmB9OqyHP+JuuMzI1fv7S+GbwBRXt1HtHvfMjAdDvdrov/
FbR8CuLiH0rxhAYk5h4h/v1vv0uXZiWO0MTmFbH2nxifkj7KbcR2yxAYHlgIj9Ye
R9VEJuSVyVA81JclWD/EejeWbC57YZ5eGcUZ9NZmradZbqd3RHMWKlTJi5Mqz4FI
vXIQNgOVHqQVXrQLLgClYamUCnJpKySHQJ0BW2gPh8TUbSfIViqyi7dQcSh8v9xy
UYLpcI0JwXf9/uCz+PCTD3Hli1TyRg+q3X3BX9AIRRS383piuxdPw2iEz48baG9V
G2S3YkGXzfSJuxAQIQtRyDbSxE7slQidekY6kHj9IDzGKE6bAXh68N41sC4EIzkF
vUlPHlI6ISEDBP3MHhNFrI5cPBIJCSFIVFKhk/P/LK4QHTiC1ICh986yY68jKfwW
O0y3Ixz+rFFpPxcKddhtSaUk85jZ8v4twZmo05hEkASmKeOHZ9SMZYpurSjuOhTU
XUjd1sBODAD85igsvwLuS6EZZHvVFuNgntKs1tfxRLOUyhMAZMCAFGXWLfolLlEN
/WcCnb+BtZjO7gxU/kqhhsYSNR8SG3aQ/ozgng2RUcik8iK7FbS97Tvc1+6iTdAX
Am9QCbpTXmgBRrIJNyzOqsjS4OBRLm+LL57NvyyuUqXjVpsXtAxK/1C7AA2KtaYS
Ny9ENn/2ClEWDr5bPcVgewxTmajrsri0aoboMOoILYgQEBKiOiqciVQcEVWCx9fT
ebQaTbrO6LI8OVKd9mH0vGuEzXDNKLz7WeMPnDf/IXoifhgILnOT5KwhkqZTMos8
lELYUW2QcWg2RaihQW0tbaNo5REMe00Zu0j0nQnyTgxi+49fRDg3mBNrYukK7cvZ
KzjYDv0v1Ph05ZkCMoemZ6akD7F7z6yPYa0ykIPTFVMUtmRFhEVKqUME6OUUcBkS
5m8ZD0YFPRX54b0ArgZeLEajWiCfNrOXvKNV0OrSOJFDFikvDGSFdkIfDTtooPmZ
LQZe8UpqzWWazIUZsU4WBeyhAYkZph9X8HPiuhuiInZcwO08Va4b1Frie04pHm1N
MW6yLKCF7saADEryp6FAShGwuC8yXlNnKy+9F94COh/luRCob3hZ5qkj+8Ca4K1k
rTxDu+aKt4cxWDDB1+S4kUsGQua9vLkSsfn9cQS1hCo0VKL3RrASPoxyJwpXbJpa
npAfXo6nhKg3iKBxhSQVF6ljXW95vokRwkDbTzurRqJ8j68XbYhAD84ix7qJ1HNT
d9aHyXrFRKArOazCTmj0chfH6vvA9SwTUn4cBDbX4vy/2i1ihAmT2BNwztMDI4jw
lA183Amw5DSoe/Fs2s66ZEJ7V/aNl28xOKIf5Su3FZILtBtEKC5kWHo7c3gwcpii
aDdIUInqlq0sgT5uic+EHi4+mGuBHx6F6R6/PT4vq+X4TDI/jQUP9pi/mUEk3jtH
15iiIKSQmChpty3F5DPhLf03vBFdCxZP9o7YOyoBIZcrdYJ6deK7JyDZ1sK7ksQ1
sqRWzLwkWdDLPFn/eqqmkmo/b16YTj5RfgL+ehHlMNZvhXJN0JlaWIB6UBB6viGe
WFdfdwociXXU4aiPCi6aYHbkpv6siYNBcSCMlyip6O2J+WYy2R/E2p3HdP1oCapn
AAvDQSKljSAf45RHQiC1pL0w+A0bXLYGan9x9yC12KeQgI3GNWEhW2iDf9AqLrU8
d2qcRrXj+668+DkWKPucAuynbvDGHNLGTy+2sOeDsu5JpG+fraC5czch83b2INi8
SZd5kFqRdlIR1cJOvIE4d8qRr8fsgBoCk9fDGndd+1KlfXXh5YCCLChzUfLoF4ra
D8UqVVub6k5n+mG9EjvOX0HYc9gPDayW78KO7xZYYknfcQtwGMmTe0hWEVchy9Y2
altNk2/gGCJExW5q9/phlA3optx3Ag65Wn2ntqriQTk34WaTqHbuIKLqOFcmIv8t
iCUlaFzVcYrJya6L+/aTo0PpH35Vk99zPu7zMMy17Pv4eUVWAk2dDGuLtkNlaqey
Jabsquh/vYjOoWKQPwaxhexVpRTloJ9grTBvoqpDZE5PF7bng+vknTkZLiCrMpXg
L52Z2etdkAuu22oe5SrQS/L9jlvYfiA6nUeIzzHXVAgQLikYUa2ETCXF6MANU2MR
eWZoZpVl0oUaNwSejpIKp3jcn+B83mKF4w/NM6r1TeyQJAxoeZDsot53X50jazfB
GfxcQh6akNY7P3ATqu+Hw8I2dybhJ74MSDjVU9SNrb8ff3CTo8+vQUPiWg3mcQ1T
YyZsDr+FtD4ac5wQ5pexF+p2IMvBHXflTVRQae/sjSc3derQRZmnESXhSHOEjPFo
AQy/uOfxMqdqBURqpZXrCtQlJklxDdVsB51e6r7EXx+F1qrQLaNXy/8Dtkcr9Asq
G54S33mxqJK2+tnOa/YtGAD0iO+UJlvIqWx0LUt8zf74GVXN1KPxh5jqfymyYvtw
cQvMuJEC36Hg/TnfBIk6N1Z5IIG9adUPizElIdf7LgKeGaShG1lvwjFw+JWamqz3
/QAbMSLvetdGMnJrecsh72/lqpI72aOcRb/hlTHEW3oZBqSDdZtlW8cteQN9pEuH
4RQLduDHjLUpQLk1Bl8I8SH0gpAaYYdEPFdyXivA0VezYmPvvQoxMV8mvwJkbcAR
E0zHgmIDk+Gmz9hcThjvDBvQT3UsMMGPKK6EBOFGLU+YZ2meiYNBtrJgl+SbuiQt
P9d6r1nOqZ5xOC2gVd5F97SeU1g73NjYHkd+FC3r7c0LZutD/pKBe4TQIoTulAvj
zewbMJ7qhGIMDA3jjmUjXO/Q9deaDrwldI66O+diKjaysuNPYwSCKxfkvl9fcLXn
WZRCu9U+RLOXQKYpXVPMD58Z0nFWW1YWjTfkbqBWmGZsNExUSUzJgmgDKg0yEPJS
aVUuRyN1ZfwiRrKfRawFcofXdopERgMihXl8Sdq3W19K3SF/sfvKxdFqMqBTo+uq
/2NoPW2Sm5QuISKsJSTDX994hruaGNHFYfEIF5jX5K4gOUSwSQyJ9UbVVWUHr2eb
ctHgmGOiZ+heaNEqoFY3Alx8jpAqrfnfeyGP1V5pz9T0YHaRu3o+xizDc+XaX8O3
jAIF+YL2loaYQwxnHA1tHfJ5kW56MhvbomojPnyit/DVtONkeiMkIEEmKc16AxKf
68GSLK5rPS4+Z3XUTLdVJ4kbdaKIWCBc0lbPhHhCfnxRVZycAdLKRaa89s8FbgY0
OSPkoqxP4ji6O+8S5D9YzyyN3Toq68KA1m48EvX+RUQt1Ng3gyupGfz9FMUj5uJt
bh63p2O6gXUcWLQ8eHh1Mr26Z1Dr6MUSZmz3yfEaGT9faCQ03Pdar92PJqgfQLqu
9X8c8rtiKwXUi+R+4n7WF4A9HfMbNBjrFK94UfRXht4OmpNxn6nBrw8C091l5E7V
KWkmLviYPsL9t9dUD2ajujxzRLR4t6VivETgt467f2VQtrTkiHDxO9O8feNdUdr1
wKzBXeoxKIsXLT2Iz08TMmVjgtMuT9gsIo0g2Ko9XaV1eD/fAvY9Ez//2qdoqKbx
F3b09ZPwHXKBPjd/NSe5OQv5NKEU5MLeaDxO6zj9Uow54JODjcNEfI9Xg4ZDsov6
p4wF9z9miWyFPVtXEQsaZyblAB+hV/ZpXVzExI0C9bPJxvIZ5OK0uQDuGdeYPB3n
uekNJshJmBOuo6a0qNgdvsHSKBoU8EHuxOBmY7Bi9blz3CDUR90VF7x4d8yLjEEY
3amcJ/joxTTLjwkysKt3YOwV1H0IZl1qR4m0ZZ9S1YfLbDiFbPUpHa8YUgv7S7DF
cjPTOs7K58A4raZFDBUSb5ceZJlNMwKlfiZ2jkUPhQ+cvEe2Xjg9gjVYBYJZ0417
ulDoE+JW7S0FuPtFA3d70Yov9vMKIvxMbqiZC3L4lLIiyhRnP0JayYGCwQd7WfnI
O26uVDyJXgJ0AfBN1gHKgt6cuFjf/QXN/cUc9A+HX8oPI3CesqFUHsEDL4BpweDT
A6HRCz3PVPXrhKm0f75NU0Gsf8zVkWIw2WcbBa1e8x5G/Rx0ywcLHy33U5E3YdZq
7MCE/++PcuwvxI3vy7JRGj7q0kE3gUAVPSLRivuXGmzzEcRH8i/aXhLB2WD4N3A7
9bTRHVek4o1KGp9/uy3Q57acZdD4pA/70hnLvmipIOmzzpVR5VcGCN36NcsuByly
tYjkdb3nxPZnWzjMLR1KtdQ87zjBF7whGv99yJHRu3cmlpZf8Cub24dhymdGIPBT
Rbqg6Eck/7XJUQ3dTzwmYN750pn0o3wcIAyTtBQhqx9w7jjD06/fFfQorrppcQdt
lJ0idWKyMr1SoXp4HaU77ymeKuWwra4lDSVyUTAtAsf80amPfvvhSu/T73TruEJ8
JrFpKJivmMKsJ5taiSiEfRAdKPCICx0JT7nVko4QXpZAxyVnhaD/B4Q6QDxeh4A+
RbX8pvKXLOtp5rFJu2dcA3a9tFlhppP0sq+ikIieCeuKIcg/M85VJIqcxv0P1m1U
nVDoW1vnOB8II5hi18AO3qZS5VHOsVYlnaypWsVnBt+OAdzTI2SjmHWMh/nH4IaC
ceDaheZkH7fkBsvkdCOpNjIFiIWUNQ/iiSU1+ahiOd+lmmysIILuK0bILtrVw/Bg
A8YsBY9ZMDDUJiR9sQ3Mch0jRKpeSNYomZAXI0mPvXzTHwy/Z+g8KW8hsMRnLCnx
dlRXewlgQOtGSByz8YNED/4QL2WOJ8+yYKGdrJHqai5kb9J661gVpN7Af6U/KPP/
8hIn4j6mjMoS7Df1dfvwU3ZO0YOS7on3ZT0ztZAcFSIzsmMPeIgcAUhcgxUOPiSE
O+4q3KbRf4fYvmBDWmVLmhkqvT+DiTa3L6hxbf4k6P482p+dm7Wbzh2bSFuoFXdL
LXlTEGBKDk6yW3UECShmBfqb7ZWDiNMGJrnDWohCl+HevNMERhZmI5wSxgqlUDtM
djeh+HxAWc5HcliI8pK1h5VsLGIu3iyk2hUp7tbZLzgyoeVxzEXybwx6EK3tYkiI
GvCpb6XPEcW7smFfEBNpCmWvhEjSsj1Vhs/E+weNkK4vOgorkd3nQzjmiEYk4eTO
s4nZijDwiXtwCC/b8ARF07bzALHiyAd25eILlRo19TP0+ya7cpdeaQOP9Lk91UpE
LX6mWQdPBkoGYEceHK9kruXhgceCtuwtepb1Oz1DtxdgD+TTTGuDPrf4yCIO8+kf
wXKKbBh7ZZrrNC3aLNr04nmp6P/GupPiQOFA4SxjLvDs5gofwJOcUePIB11FlS+0
igr8UsiUfjf3dDN9M2Dnqr4XVydEBuVgu0pd/oFwqzo7VjZDCVSqv4jZWGauDS3Z
miaiYzVqrgQjzcbKgd8a35H6KZE7Zn6XSFUOlMQwg6Filt9pIZTCRrSGnUxpxcUU
85AK/TiIlTOTMQ763MO9Vnh5Kf5u8zCmXahAuIrQJqCOAZRT33hCWU9Xh/BCKaYM
Edhc7RPRDKF6gHyQPYiyU3DKUWaPu6pqKfrxw7RfDfwvKo9lNiUOfm1cATFdlf+S
9u5l9Vsh2N/gxrsWk4Q6er6K0PIX5aKyfJ6gA1mCUQ8d8rwSHzlLXu1vJCar0QV+
BknLivYJRiDbw+cILqFfTUkzbCBfW1rdxeDrLivp5g3mBeZcE1zVdObMh2i7BeAQ
MTOteYfWRtQZGbAVDcDKRYpf8IRWhnhF6s3f2sYGxl4I9O775Q2zJUTo5GtmYJMI
M3e10JMAsJeWfwQsaolSvQnRV7Hj1con2ZRkwQewvnslGy+UHZXqGhDKZIQ8SDba
RG5Ef0I7AHnvzDyOg1ouwQgS4uw3FjD6D3HvnZfqbLMmtOimP9dTPvyOwwfnzHnU
0zegnIQeDyKkdl05oGXsqXRcfHVgw5KKHzLG+PPjyNYOfSDlKJZnh7Hvm4mSHbv0
oay/8ETAxsPfj/TCn3s9xlSOEOZU6su/8tTNQlu+qNMw+6NoaFJj547rfT5Y9OVn
qkRCbBOPb8r5eN2BbaQJhoeLFyW9DrMfrM5t96/y9sbBw/pgyfsqNgo44ikTQlJA
mdxYkry975XqfFkOX/VUQHU7+sHdyFtJqfJOZ8HL39AI5vwTrRbASReAUt3HzDpE
ck7Hym4Ay0b0o9JgnonTJMDbVLnq4doFcOc0eFMPDbQ5Oj5/d0wXT+Z8OsUt4oM0
L6FYsFn0ai33n+2QXrlOcv+1bVWQYvtjrPrGE6FTHhbx88c/tPJEaHkz7fBW0J+b
Hpq+kN4ax/NE3TDgKP8qBUGmvyYzxEDO+byVu6zj38unpjToJbBWIChfmmz6a1Xm
lUw0Ar1/hY/DN/1XNQeRnyqoiWOjy5YeDP1dOnJgmFwWY1YiaVBgkvEHeTFfD3m8
JXgbQdrmBVpdWDad8m6kcWZXeBw+5lvvGfatt2oGpECwqQGOOXeHYWHn4gmmp4LW
wNjnTGEZLbwzhZPNBOCW8yH/kFyam/DWtkfQu1mLGr16vh8HKPyuQMPJA0CRGraP
K+bJ25chllU8KHDbG+wFcdhPjbNBhP+iXBtPUnH+HIFCH1a7DvScZ/Cd0BPqHKc1
ZlyuGAUzR+EayzW6d1fYAs/1AvFOQsPdo/hFFsZcZC+EBesPrDo3oxIFnJzDzj1f
ZcIUg6YVeMqkUtm+3eHwIgDa9MMn5yopZQH+95r8Z49LLzZS/5swJR9e0D2EYsbN
emeFA0TzcPcw7Rj31CkRW1YD3/K99Tc74Upi/vEni5zoxh1E8gBKYn/n6jA2V7li
akvrJGojdjjIo0ntyZB8Dd0l9rjLmwlHxV5QsGdysXAsHiZS/JTxT+UgysOI7wmg
OtqtSS0JoDGxhV5A29vKsxsOwrdPp4EtebBKb2uw/KHOBx+luuov3HrVe8kwfOU4
Qn/umm21ZUFHATcV9sc4peYNnX0FsC9Rmz0bJqHfZs94JmP4NZAloNiEIeS1lV4b
hm5aLnt/orIQAs2tRhLaSwK5g2P518qgZTq9UnzvAWhODpiULCfE5iZIcbwAUErp
zZEVfKAFYtURW+Lv1wZQd+QjkbwyCmNDgA4cukxKqc5s7ZCmmCwlugjfUFlo0Hlf
xzaCloxCKxJOjYBMbQw6ofxo1q8bDCTy/fRqntgiN+esDCJvaV5QEM7XYC0GxK8d
RPcUqo/H5bsdelLT1Y7c2tYjYkY8OGWK+mDQIg5dTQVLdixpn47Ybdf6SDCjgoA6
moVCnawIEBjdoDVJ2ByJmNMa6i4on7Li/Fc4Njp6JuaSD3yPXwR8o4QC1LtE71GL
KNyTNmCILzU7PSdCvCMQDBA67S9grdg6UblNgw9xMK8GADRwgfTLFscvHxhMGD43
NbYvGCYlSJkuCRcRPyt8sm6VO7wY67ErS2d5F0kMKaLHdC+YgNGlDuDazshfKkfv
kBKU3eGfmd/8uFTIxXqDSsKFxQJRJdJLLus8kua9aDzZM548EevksaLenXw9Lx6k
vSvsbAP2aThPp8Gz5Dgx9gDgFf7swQJm1XNWvZAeE4La5+rPm7U63YtXFjg3aBkW
MeujQwIN1BrfAa/z4A+fCfgC5ILxBjwqCiQroi+Uzn1BVRUx6oGT/mhGOz6w2nYr
F84YKod9eZRvKh7V9kaa2VE8jEkQ4acDAM074qfgV0AT7vjazPFNW5HGq1joXmaQ
lZ0SqZi3fpmi/Yr6IZvUMPSByJlIZVXUU2x6qBSZGglqMARqTbcM8X0AWrlDvF/B
sucNsqn3I/7v5dlEFKkmt5OXP27a4JRtX6eFKbJFV8+okZYsLJB48JejMrCuZMKo
6FUJ0D60lzhEZfb52WF/WBSmQEgCgdVuF8h5ROJWFxEo9Q8qm5jfZbYVdeyEvEFn
IF7+KgclfCRa3iqb+TSJ1YHIdf90Ytn/80P3yKImGIfJjcQAOOjtLY+Vm9vPb9mD
KPmRmMkfeO+tT27U+duBsO/NH+mi9BNT+EGyheSDzZTL+f2F5cX0TN4b4bNHyHcJ
iCUrtCvt4eczVrJrkcaU8IiJ3V4r7oiWHFAKjkCFqL0Rnc2pDjURDTOiEZD/cAbY
QksOJ/CrD2Rg22GorvB5peDoD/rHnM0/28QbRTQZ3pINPzR97wJyW8hWwzRhpAhK
YnzHV2e3meraNB/sCNFMWUyuQF1nPeaPfk9Z7pQghJ5pS0YpoGi/mRhwLhZhHJXA
QpiyddqeNgzHeGf8kWIPLmCh0zjXq88dJa5mVJxZj7OSA1p96qbIM+c3UvqLTL8A
ZheyIiuBe08yxG2nd1VoLWLLuZE6mJnOdPaFdYDhJkEGl4Q2EjAKRwodUv7riWrg
bEQRH4311PCGIzARShuligQJPGm505+myyr1YW6M/F8TmDuJf3swpAyJ9UcVwAq4
QRg0VO9NuSpPolIDuR8Ynb37rumOvNwb2G0OzbiQVWAiCqbQTIF2DyaO8dMIrm7+
+NpMQj5Q2mXLntzr7tuRntyn0mmLHaIQSxsvuBgJ1uMJZudrCkvhsozh0vYZzkjS
kZ4j7/vqTyngUjnxjKqnSYGm1ZssOkKLbSHnEwXCBM9/Qj/7j/twhnF4KNlmj/R7
B84KjkQgZP0kD9kGmGpTskd4jsuuwKWPtrqSaOoCZiijjRzGfwS1oR6YI4IX1v2o
rSG2KupxoWlVksdjrQ3WX2iIm0m3/zM4M/HUwRoXyVV9s/SWH4h1IQTvPx3sFisq
MKi9ZNXbgWu8f0qzRTFXUFt7uPxy+GzcR3j8Vok71JQwIwiik7Emtp3m1kiU+g8Z
3ZIAHRMwCFxtmVpHPIb1dk2daZgtKEoRCuHB9K565GaU4s06//2IOI+zx3kMRTZa
NZvQoB+/tA6W2D/+I3f9hsLn/szVpWrspquSwc3ZAu1Lyq8xR7oAiYhjHcKGnUFg
Yy5fF69EFy3B9TiMgcWKG1t5LWpG5GxZsLXgYOQwMOVBjvZ67OboN1GzQM2BPslM
q2+50R+YJRRHY5kzuG5Y9FI6VCFrLy9o9dekCLf3sEy7UVWYtoSz7phej5b0x9Lc
81yTu3f/PRjWOuzHxMC4edG5+974k4rFsSJYMubSjr2UXBuic1wQl70ewbpdQ6hZ
hJFBdTZ+wEVvaIhsAH705gifmVMgq45CisVSNK1BuzFpXAVBJqVsKtuvWDy2WZ9G
HMippr7TZSRwNhFC4WYtXua3MI6HZTyLGy+C+36XExj7lqDz28d9iwKhAGLFMyio
AVgv/lr/0CXTHgObEV8N8DlFGp9enn9W4iJsi0WyWScuX0l0l//kjxV1taqihmqW
HqyKPqPCjJ9q1Kxu0cytzOalPXNB25btpQXBTKwPizRpzyhYa4qwS4ilBgSkHXK8
wfZORWZnMuWMPrRx2M3R1W5OuVtI+McyHGpdedMf+Zk7S4925q1QEgvl8RbNWTi8
NLk9nD5kQ/u/fwGdsDpPLS6tlbuGggVC1E6c6urrwLX/wH0kCmOla1WFaocQrMSm
OhuRIyv2690ocvVtKe3aMvOUpai7z8d9Y8jjt+HfJDr7+ElQe0XcdfxeddaP8C+Y
aM4OGKPPLnALjo8AmQCQiFll0sm17H89jdLruwoVtKWkZTc9lOgDr6ZI754Kdrau
D1l0FNV34GW5Ujl5McWQKILM5mQTT+Mcl2bX6irNwePtSG9Z9BtQ8v4girZEKbj1
CTReBJda/d3QOGMjH6PUbLvGp23akM5dbVTtUfXp/7y8hk6HRBzTrdcGH17HWLOc
CzpooulO4aVSp0Ci+RuwPxvd9fx2GkutfM4H7VNQynpIU4INXlqkJ5a55RWxgACE
d0KZSzARNJAVpYS3gg/2WY0hE+hE9nG5HfAdyufzXQibYdgO5w5UNPMr9LqRCuTZ
wQUskJB8nbKvZNBxTCrRBjLKTpuuz0ViPu2ULUugIbEWvADx1cIQmoNuI0vHakEr
hlyS7OiGIWPJT1Sb8aZJrDTts61KjmJK7Ys2t9mZs9AaWQXj4ztAT1qTm4Tt2rU7
myV0ph2Y6NpbASntZCA5Rl4VBWU2la5swzQrny1/HpbelsCR0oB4M6gCXBiDXM5s
CHJ7noJ/X2XfhjVOMJAqVhPYoYwsQObJAdaOHBaNmcTH5hioAylweznMX+RUtH4X
1X1n1cp0P8lMPmPqohGfBfSbJNCxU5eJ/1J9KJOYvw2G29Yutc4ypLz97fdqjDIz
OjNYo6VTFkIuG5uxhc8fB1OsVx0CQwt5lF3ix9e/FxEz1bRdSU/0ZTaHNZCKzee7
NhHbODsaZOws3f3G+qZu94TB83IygxrtbY7+GXWzsSSKwQpmHuSJGhsaG2Sbj0iF
UojIYCfCWEo/RITqd7ddw5r6lRmAB0OOAyrdb9HRW2p2uz+LCh0oij2ePbk9VWV5
Bpurx529k6SqbSVC6C9dVwm0xdfTYXR9EjI5OowovvpnY6mHb6GA6EZz1PHvYnLl
XywwK2X+qdP2vOFT9YdMYlxa8mJA8sG90WLqmD7qMKqEOKlzRPPZZd6stVKW0Wkc
OX4hFexPv8f5JC3gK9FwNWqFL09iAl70Y2YGWUFtfUE27vuueUxbB4yPZLAKBmXv
NwJXnYP9UfocJlhdhH7y+12JVAKoS0UHYBveErnyD5qVnyJkSdQ/ZRNhDdOD8P5w
gw1jrVdInsJ+uev4/kdEwkojh5n2K2miNlSjrx1Gl1xGqWtXCR1TusKt+PEN6+Mv
9zvxy1ruWnpGrQtpWF1sgoICtcEp7TqV2RsneiDATIpTyR5U/Lv2w2hhw/SfRcFE
yV4WYTiILA53brIVHT6Bh8uWMdEsaMLXWQT0x9lzFYzLZEliDUn3g8oE/jBzY3Y8
+rpmFcAX+8248ePn/JGA/AhTBzoVHAbQmj5KDgztyunbVL4g8teD9PWqsTnyorUw
EXURoPf1AlhdSjUNwO2KUOLnE+/NoZ511LTfpojxF5h6DXeV8uFYHZuEbNEuNdru
n+F0yeEq9XqQ+3C5GW6YrZZcHCZNKM6MfoNTFd+fASzTIsnols8mkQF5pP0kGO6+
ylGVEjREX8RK4LGQ8Fk8q7YT1GsXjupticxCIxVrHGULCeabUh7mM4HRMJh3f8gl
bMNU/mkethW30ywX4vtb7pyqJxesswifURfOHjOHigI2CjBtDHHI1tLx8i2LfgoK
JKmXLNLfGPb9hmUBfKeQjIbsnwBNHhcwTIHAnuwOo3ewzFOy6sFFqZceaaSbJ9L0
LPP1voH8XvY5Jm5ohv7s/T4XpvrhQAF1nffHWeXSr7AbimdvxzudmmnUh9CwVBRQ
0BwTe99fwgyiKNQmfHLFkL6zILXrOUZwruRUlTIRajN3ZiHZPwNAyOySsGBDS9MF
Fta9NltWBJe+/XrIHxjHG/oBri01PvWNES2ahgn3VNxZQnHLEgu/sB8i/LVR2mTi
KkFKHr9r7m3xaHT+aXzZImVA3z6s+3eAgYZB1+lwfwxJrkyfoSNrWYBlb4WMo68C
Y0DJtGd+Q9AAM6Hju5U7etCnsR0MhUkijq7Zszk9lIrSMb13to0x5UChnomP3SwP
IDvU5q/YAjnu4V9tZLWojd4l+PSGPozJR8grwtjA44LwSD2WA/HHXs+lJ/x/Kcf9
4gp8n09EfXMrrB+7IdoBMz0ofbwYsOR1Kni+poJYnU9GtfNGmq6hKWkQ1YNHRc9A
TyXFgSjsFG3R8/AbhO+3FLeA+f9kYfwNrli8e+L1lGITwNgkTNM/Zc0ifzSwmqxa
n2PujG9ZORV3CNQzoOqcvEzusccc3Df2OWZzLv4P+cpZ5EJVq6BDsL1iIfvDwl3Q
E7nUZeXLrSQNCqvl3nDBU2edB/k1R/c8a1vtwHjWlwX18wY9MQYZ4wXKXXRW3jCA
CGzVxa9frQNNpb+y2Do0qaWEvxXV8W/REMIZnoBed05+UW2+n/dfO2rdCi/QKn/B
n9zL4DuhEN9lVkecR2cGrhm/Vsl2XbHK+8yXp0ZrF3jVxv7zkbADWfwAN1Q+J45Q
RGaZKonCCgX49lLsmNiBK4kcP1cXsw6hHJaWnr3abO4RhLIv5T2EgVjGERDKeFQU
62Z/9ZjzU/iaZ5eEL5RqDsswyzcnfrAa0osH2uneBVaeRs40tj8OEhvRQlsulRmk
+ZIkh4vbQ1TnzqL54nu3U/v0VHG2pQqg/v/cCh5CpXB7WJMkfzrE0xOhhucLkHIq
xXBxBHqarUj7UgK6KB0hQp2GH7JJck8tvR9TOT6TeSLib50GnflCfwLW2PCYSKex
aCCmfxwNGE0nNd65jgEEJCPL56aAKReEx1odwQD+6FTyMbxmUaU71rzWbIBPB7J/
AQ1HGkhgsAtOAkRpts/+4kKTBpBwssFGqTDYhKeEAjC4fQHhxejEPkB8jQ0AL5p8
9uBXqnBgxEVoeBcxtB0QHz5PY4Jj3z/6v+feh+1YXnFPRj8Xcqq8zFxnCjrnMM8r
usKLkKa1bVWqBTgo1scf40XiCoM/JbrzsQ/ZTZ2n8ZWnBcDCnTd//77Mza3cU5qh
Pqi2to2IISNpoRP7QbggwgBMo5EAxAmmYqQJgecvJogpkygBixFapfJkyFs6Yz3d
abt50jdWcqCkCKytUAeaOu+CavojmfBlN3ypar7Z7qDCgzmrxrYzKbIEeTTcoqWH
fKZCL8seUSUEefWz2/1PVU6D38jsHWUqfIK0JeVq6qfYfan6N77/qOg9Gfh5wAvH
d8aXqcT8z20g08xdu5hEun+i2VkD34/gDYGSMkpwvSQaw5AAXYnVzy4DCzcNDFqv
bHCdpHLQ1MDVv1r0GV/hApK2fOCitlBgvpr3FNUE3Dgf/z0SScJU+1AcpnczzTjw
x/c7KzUNzohpgMCIm8hbVmc6U3o4d2ZWgEpasNjLmY2z21IOEG3B4ypfXWXFa8Rg
dkZHX5MTAPuJ3+P59+0TXsXr8zoK46Qk0DQhiOucJJebWDoxXDP6McSlrV5wD0MC
lFgRUhQQXzDwlBiRJKaG2jioWu9U/djIP8HsKP1QhhlvETNuMVJzLWNi+ss3mUEL
/+v+rsBqEtQRFAY0WhOlpCDtRZe5JySaN12iE5MulbLBKnsrXUyqKA49EyQCICSN
qVI84l2qvLKTqG4WmSauNIIvy2EKSaHbmDBOjN12CTNUggTK1TYArGLSxo6QXnn2
H4ppqIDHBUSk0xB6nhq8OeQ3vhU06H7sa1HueIXVb0ZsRt0rKqQOg0M+Yct+zWDU
wLnB6oYvbsjzAzhCJ5PzYAq93fr+lKURwiOIE1Mxvk1oW2XMP9gJ5H2hIbhsOVr0
EgmsTvB+CerC2xbenptWoUmy6z8TRRDmUjxJRRXbjZlNMw3d1Cvb996bonfVQF3L
9Q/HNlOu3sW+2b5PWPSny/hghvFjwM+uvC0YJp3lTy4fMMbwkZ4Go/3HeWjBYMDw
7KT7Ev3vJKJvrNl6iSFyjyTsh9Xelomxf3cSAwUo55f2oYRdsiG6I5DEG7ZRWALP
msQpVSALXIF7jTRoAiWXUKVu+VcQ0iMudfKXV/+A65fDrAa+r63/SFNuusOLdYOU
d7rkYOWfm7jMJ1g1S6OPltSqrm0BGFoF3Q9Q6IWQu6dDayxyj8L25iIxaRGDE2mn
D60MpQ3GQUIQ7ZbJ1F28yedJ93ycN7GKrlFmVU2y8RwI3jSw452CJ7dpfgH6G0aW
yJ79bygKH/3XCp53oTshCk9FJwvyhPWArcsh5PYeUhE7nPYqW5UAspfOyrRs5dOJ
OV331t8nPOK/UUK9yPNKRWYRTjhX/O8i3Cu1BxFcSc15eCO+B004NbC7Km+s2o9V
W0q5EXREMwVm4mg2V2psrsg/e+sOV0UeTpEXer+qaYr6pG3QSo8XsrSd4fRJ1+LW
irfCdMctNGZ+gW4iqVKdIImMpAvsDzD2qlCyk049NZy4H5o0/651kxx/U3kUTOBY
e8QWtKr/80KlmQXNQ9+qiXlhtiS8E+ABB1aqrzkW8gIP9wzzBQ/oacyNgwgkL7+d
LO/KF/vJvgXx+gW50IwjXfK++9oOseT1HeuCLB6sMGbUSC2dWuLSiPzUzb1rO9JH
opv+sZOL3+1moqbjNalfZjINrHOgM5NQSrsXyEWrhMiDhqjcTViXKxCWQiw+K8hW
P1dJ4oFS8qN2Ta+F+zjA5f8bVIWsVaswj/3VjMdDpoXI/EQYyFBbiq2xZrh9xbIf
1rDhsz/Ztv2Fi5PZIY4MQ2Tm3U8L6EwrnI8CXD9lhnoH0+2gpIb411y+eQZNCwwf
Sr1DOXqAUlg+hqTxDVJ6cQWYCxt46wuKVa/YZJIVeCQMxtG0fZXjcfqHa25qmy9n
kLpHPZgSToJmKGWSsZw/OyqFiPl9ZVe4CLY8tI7nvdsnqD2w+oPSJPSlIqzok6Wx
hP8KrWWR42rqi7sQE2KopTYALyBmt+nBneKYbif0pMzNvIJqUsDj4Sqg+opXZL53
OnnJxXj8H/cSs0I9yxGBxmv26miUNohF2bVtahc5xh+660Va054mT58PqLCLVgEI
EMboeCp2nMZnbnDYcaZwcCtABIIPVXwywwZu0rL4y33RyhSGnzZeWW+UXyUYBWAy
nEQdslM2sQlsXCmck83F/E9x2sqS+etg4aRDYpreryCvFLcLB8rUs7Cy+cP31+hD
/SFiHr2hAQrJ4TB31FPx76Nc2XiSAo6BlsSkA7Xe/56WgaXmUUkIsLNxNOOWTZ5j
73XRinWWHR9dIoC6ge03mh0cJM/Sad5VAiP7tZW+iwanFNPSSrPD/HOaYswGuMMP
58GkaE57GD99Z0ZLrpuc+H5waTVS7Hb/HJT6AHYOEFPIsHdBz/HWHrVmKg+BsGdM
3o5Xokj9oUFV9XyAxewFRg7O3aVnMaCJmCChipStY9y48fUlezHhFi3HYC3A7i1S
m/ituVMRU744gx0P1ERTpfJBIIEyxu/k/8DPS1SQsnBSyaZZUn3yz+q9xKYrwZ7z
BuyPeyJGz/B0QjVHoYLwLV+9rho3+qlIGkcjcEFwbsO9VHvTXQK6Oj7qcbM/cMoU
CqkQVbbqPYTzpsolvgO8iQ0lxrUBx6mxZPha93E2L1SWTafSMMP6WX0/ZpOU1VmI
3fW15MtMd26I07r/DudyjgwF5THbguyy8vwMvzspL1snxxTFjkiPeb5KOJla435m
s8PR3rCSAVbGMUMQkvnoeOjPYtkRKY+DkC/+wSP/nwBVnCKFbc8ex3hMfcrrFanm
NcaaI0FlPU7ASLjNk1sggQMMOZJgvmnv/OcnJwf/167aBbREKIDVYdvZxN2C0EEf
kDgNyfYqM3RVBd70lKMKKLCO/f6ehyiKtfHZG0yajNb7I59K7CTrrnbEddOQOx39
nHecPOKbniZ9bflSbnwGZB7sn7CLaRhLdt8dkmBa8myXAyZCaTZYDqkurSZKnpUx
uq2F2M+sC8RhA6Nm+N6cBFY6Cdoj3/IEYvjx/7crek+wjHyvfXIEyZk8mARG5gF/
VUTNXBdGpdEyWWbmba9OFLZ+3N2Xrj4MafA/bymrtcujvUmV0evP8hEltwgWSnNu
7dZ/ngiSm9+CXzU6AcIGCclKoBoaqJKIHEn2CaOwAFPm2D8EtqoyULMyhJRcsrxt
NfiaBeKyBqGDqVvUIiBrpq1PPqF6POwQP1hVYnL5PkFC9r+H8ZLDVoJljm3toqMI
Z0+hTgDIOsU8Mo96Sz888hksF5aLRlK0do1BdiC8gfPm8i/en0sFaQdPMwPm2w0K
Ywt0oFpNlTcUcEIlljJKpg/yd69a3g6EgRIubKjWMnu5i8o36YISPI5yu8aFxtrw
CDln1KJxL4lJxOHP6H4S2FQPokzrTeB5bYiFKQjNenp+lXCWLwVOKKDdiPwOmJXA
gDy89vV26eg+3e9ppb5r+wfz1f3Gp9tia4Wk5uIYwuJ5m5V6npvpBRXKPsumEvKF
ZTYnAO7ZXnQz5RqkMNM4pezuNnXobZWfacpRmmjisE5SsfEhvRzilWBEOywtYLgE
sI7pZ7GdsrMjqQrRVIDlzAAN1HFoTCRZDBSnUHYx99CPfOOw2uYC/lOP16g0yIHV
ds4Yc7k71MTitPcbncL0a+8KsHrYfOm5Upn58ickyaxetGOboz54Z/5HhNeg6Grt
oEMUNIE76bM5q6Rq3gmj44y7xdEUVLvfPGS2Q0MERhRuNOVUHyBJACuq+SdRrHhN
5MLDoh4HCNWpl2YupfybSgrceVbqzI0z93lYWo9+rMDWc3eBa5WXHyv6/zB6Sbkg
Jo//meHv9O4tZdIpTnZzLRTmbtBeW8quZuAbfLJNwmB4iERDZdVFjePugjaSqoyq
7rxH+tERb0S9jZ3xGhAClqwrN1XUsUeYxFQj5cPdZpdTD0sVI6RDCdG4vR7ELjf1
eq3kSawKEMgOpWuPWH9Xsx5+0cVLoLR7w19Mu76cWtwgwS5oIrEUHhGYVQl8LYMu
RBZJ40TI7O1nvHvOzoWyJL1eAq9PtcYjhblpBuF1YQNoXf4enLjfnej1sTABLs/e
pqjRAYQASuw1saxsB7gInJGKcchXDC7K+b3cNVlxuPnIVWvzdJRh+uGFn8Dl2STI
Am+NoJsnwaahMKek8EIqiFISgwPxQ9jR/VML4gjBrOXXc24QurjZTdMurdMGc5hE
OJI9awnq9N9nnoTEYHG3pVBJj53eeUfietQ/0yx/ocZjouF5dG5LqdwiYC59lqPv
rZ4OSrAfVX3Zlv7OfMadB7eo+DwhknwDS/8CKGzmX8RLOA6kNl6mRUUj//VSc8M4
EikykqHV6K0RL339iE+if+OTxJu4XwuqKchnS8SWMjJFJ+s8wGAWjwlrQE8ogrQd
N9RgNrF/nNJNso43VDjfSm2eWscU8YKKm0axVFRTWHNLLHVaWRn/914auDjzAlJa
cMjsWmvNuyYvgfxeSygHnwywJwdzCg8ioyDhigQ3CE7iocPfTm9+X8VcD0F7Wpcd
pkXcq7WFmUmy4AKjDbTvfqO1MYdsVqOSWoGpQ327ys9ghupAXq8gzkF36mmG04Bt
V4FYomXwxTO0G+Ky5xn7G1FSrGepPxYRqd7z5bXEF7AoQUDL84Cpm6hLXE+Q105p
tbQkBCgIytPR+6TdDgx0wY2cd14fhVw8r4A2XsPOcM/HRl/HdmJeqd/rAG5rqayb
SRpeORIuXRmweRegVCWeiA+aFdnBSd66Zlxd0pJqI8PPApgMTmoQCpXBLWGRj098
58DgtzomwNHCQNhUZyopWCuaMbHv2lPFUjLXHLk8uOGjL6EjY3U3y9OkrJlSY8mG
dfNoU67dcHx1S53bG6eY9PE4O6e5W/beLQ8hsjFiOWbMowChGjfkYDbpgnzXahBH
6oGgETKI8SjQr2xnVmpql6Cz2ZzhP1YB7sN/Qcdeb6SGkTCTFEUqRpR/HXjPkcEG
tADezrOZJSy408LbBlTX2aEeQ0qeUj6tpmROOfhFW/jjIbpdb82kw2y9yFHuM0sQ
lz9xyhaBJlFVymi+8Wwz01RXO3PQP5L+3Lt0aFPYi/FGUp0MW6INv5GQ0fxZyGo3
tBXndI0/paDPmnDJpb0nM213FddoTm7XHRLoJil8ENdU8ZBfdG58J+enAFbw7159
HBXKOgsOJmlUgkAwDAQF7cyUzJ/K9IuWugyQ+a+Tbdpi909Tj6cuGchg2kNo6Cu5
90ahqS0xsxKOC3ScctbDdk4LJPxV7uAdNImo9qNYOf0UIq6COUEf4kw9RBVgrRhT
kHxWGTG8qW915fLpX9X8BlCAbSdRzi1wxxQDjc3FkAQgD1lPejodvUAjzRde3v44
RpdyXliNjICyAT2erpC4gNlEuVjuIPBiSspPu5pV515omJOmvfZYPG3ZBszcXXsq
utg4+nFiVfUgRivTo3Aq4Y42K/480DiSo8e72QIny6HniY+Vc0S7KkoYqT+oe7oH
OKbwbOGt+oDjUR2quKJRhJf5rvXT4LPskLhrXDLxPzNd+BUQec1ZkWyLzBwtqpPw
07geDqjOXZBshYiJIxy8lLZE+4mgjb9rJsLoGt5Y04D8dfzePCOLb7m7b5Em9Aw+
ckrOjeEhsdJprKZ1a1/m4m+CuN8+gZzyTNXqdMt/ouo3nCuO2zek6n8c8vRLZLso
2dZbe+7YWOlSKoDh2AJUR4Sefc4OcuPMMyb7dqXrFI3cY5PRXX5pQYzF0/W9uNiJ
bpCU+CAchcktU6ljUhUxQbsd1lLLa4biuMeivVsU9mqYgh2iWLzDwWxyDQag6CC9
C6MgvZY1xpmecfp+ALakJVQh+LhhvqTANKMOYJJlWXvaHNNRAAHhxNFkSvnDQlwK
DrxkAkdF6i/YZNoXFKKKTVi3EpFWc4QNypSB7mF7MWNKmH2PBTg/rVNm0H0qfLkl
bhDUtoIn2FRAHNWPIqODQubr+HXHqGBvhc/ZvvPqkQzGWA/KqNjN1Z9k5aH8KksM
3VUWI+cERT3pS6hvbTMYmLFYvyhGoCmQLrZbPN7M6KE/Q34ahhRtMOAfjBOrJs/T
Kz/6edYVrWQI1SrooB9cObN1Bu+05ykSBLPtsxb3sFc16BsdKPAvWXWoNwC/c2J/
owJg1ImEdyDuNvRSQpvucV4YDhGlVY/+ffWax16eVI3vA1oYjn8HsXuij4h0v3rA
o+KDO1G45vsnFAS0FJSp0y857E8uxjfU3k7cMzjMaxaYNq5ZJWxM3yTNO9xedIAp
1s9zxXAQdzU28HeDaPG9Z4RLm6gZwOQtTH+Yr6LTpSHwev+qNUIvK1j0fPivNz+g
YwkD3M1eA3w+csNLRARjIKoHQbr3evo1idwvcSmn0d5xU4vA48sZGH190kPcHd54
doqnXSiHoqezsQoScNByjgMz/facCpHATPPKLNVTmRkBN7yXrq/iEIA6eaeAJ09o
WdFYHTo211POP3dm3okC0vNVTnQaGKBgVLiCy8LtEwPkbxloNq8uMqGRXDFGQXhy
IcylMJIBGAW6mi1iGv6rXojT8vhIG+cmQP4IKGa13sD3ASRVHCoQkl1TC5xY7E6e
jXdeukvjtkXpBk3kYSd72AKgF2MRzwUJddi8tsRSr33ViVSWNgYkEmlAySvg/LUg
CePJTZ6UxcDmNXi7hLbyKgF7KwEALo2ekfTm60y38PRTsLzy4+J87d+1aF3c6dZH
R1IpUE1lQs5oafN2dLb/3oQjJUjMvzuznSzYDfYz5XueKv4uYFYP0swAmCfvwKsd
qQDtJ0aBzuRojg3oS1BWI3WkamM3mfdLOn3sOS3dlbQHPLlz91GSmwNqrYNyAmIh
Q6nMJ+ZqF4hq76V6X1eyEOd0TRC31Py0yNH91enIki6IkjyjQwRGwqaOGJJYTUPT
OWVwwzu5yrujeImacyVwLYhdDWJ5j+nDVxqy0K/EwCOnX8aaPu9/791sYrpWuGlM
5AOS9FlD2WWajousadOJeuRYEojXIJ31IdNA/K/x4gxU5lZJ/4fh2hhPH/lWhaOY
f8YA6O8f0EaIWPklaPiBAoSb3c/rPJLq6xRJgsgGgvguQMaSKXAfau4ljBcNx4TV
a2DnsryPpQvU0dSifTI7QTveB78d/EHEdgg4rq9J2WhnC3LyuMlfFJWRYHJk/RxV
elrMEk6QAwiuhrF107QdcLTVSKbhxePqP6BFYaZ7dbmC60ybw5WWFtQ9wCy8xnrG
ydymRR88XqVTz6FRgh5QZg3T79NXiCeOYs9GEorJNplNEpW2QGMwpjPe2ywSE/0j
pT8nXvevbFnUxbbaouF3PkpYq7OCPNpAinOmrh70loH6pGMTIsN5Pik+EYdDq8R+
MVKeMxztpxTJ6D/tVfCd9AzUXgYjbot5KxiPlKRcATjCr/4uMm8FVmCyaHunb6+X
IdopNgacJrZ4yI8O+wtAAT6ua4XHA/MQdNG0QQDMSDJ54JwLQ+qyiuUqZEu+tDa1
fc2Q8y+57E7cZRw+fHCvcFwK/Z3mtxPKvp0Q9wwFr36KvDSX/vSedax2yGgDuHtD
W0x77di+XpWOYc7FPuRQF6cdC1dExgjFND4cD2IzYN/Zcj9lAwbPhh+9jcNsNBDM
LLrAsq4+azsNKtqL2VEf+TUxN5jIqB9cbbApTVYE3MG6OkdY+4QfOIypYA9QBu/6
2aHFitdKwlwGwDEuZd10qCctSBzyIHaWysedxGvz5hIgYR5EqIuyT/VcRE04dhbA
DbNOqwDKnNVOJnF4VnAErHU0hHXrh3pHJsCxrhK9Ari21nlRtFmi6Qy9Re9iH/Ua
HWghMjsMY+iYxeX3XUSwo5c8HDMITuMxaC4urGxAXebnUpYWOQpMwa84GRWR7d0y
YiKIcEfmOYlOOpvmviMoItneSUqf/ftdBddIFgO3YqW1kAaehGlyP1eGkeAIv1z4
BMDOG1RJaRiwVx9LgAimVhQAT5nXZNdwWk6k2linYxnIcNlo25cou+huA8ZQ+nM0
30A5NYhaQQuB8L+PPatbIQrbdMrHe6oAZjGhk7Tis1QMj6CO0uhUqceKj98zwtzA
kcue4HKvZWXxwK8PCbRx6nJ3NaP9HUw0t3TzgZHbkM1t603phcJRzGLGgV3pYfsh
1ZSLfu5G3z4Phptepyyw/V3zgPXBahUKgCJ8tLfW7uk+WwjdpPVsymGAGRFXSPni
zwSeAgHcJLSeG0UrI3tqOFyhPOEpPXjg1OEIqAjw8EcsUr260KrXMoX18f50IUmr
Sx03CitVXuZo/Ax1ePIaA2ZHO3ytTY+RfGjcCYc6XUKRyxAY7ml6wws5xixTTXEb
m19bEtBgsgYjAq43jQfHrkTDqs09m0/wCbxPY0zGUf1jEmLaXLoh1uStw70mK762
2xwVhx9510T0PoUDc8CJmDm/JadCT67ae+usCwwiBmzMMcVGO3XajD3RfQAT6HuF
lfVbRWrlAvl3G/DzD5dBrcSGZy67g2hSmFC8+HatlJYmdOrnTL+YtHuIaGex24GS
Rxx+OVNaqEX/5E/N30cfa2hAKrEyYn3yyJfNJo1qCm8ZKw6tbcxIuBlrkNxxrfEH
uXPqBKnYoP+vYq6vIYoBXuLjur/um2tiM99JiKC2ptpIrx6rt2aDrFM22LkuE0xk
7gWQR0/GpmJ0WDXKQO6BdkfLbSYCR86hrmFQCaFl07XytUAQb+RAdxEw0zpS59Xw
uuSx8rr0b1oGOk3FYAzUqeneczlbKgRJJB50vWZC9TfoBYFqR8gmSRoPbV6F781+
+mCbQlC6Lg2tOR9jnfTRg0ftVS/GSvO11HFh/OHGppYjxOISKmVOXzRNBtGHmI0O
dhsmmgTySnM7X0FZzzLMjkNQ/l0A0Pwlg74HPdTiFNPLQueGmRZz6FBwl4GpBzjR
1lBGWAr+7mllk/SU26AbuO7bja3dRZYPBlWEhwOe6EEjlZyQ/q+NnRphCdJoyLLN
JC8CRZSMQG21fGDhLl3OShizM4lTlVMeg79eTV8B0cXBomu4qsVkDu4CN7aTRkoV
oQiyK+PkOX1T2lQSurB3SesBAqcisFIV/KKYLIMn1/XI4zkQ4879TJCum5WndKPk
3FgZXKNK9YmHy9SkAQC4FH7aXtig6lQpV//RM85CU+qYCHY2hPzuVsdBal4hSN5b
5qSjkHe/0nxj5RmkDXSIyI+L3/dzZq+k57aFGKNfN/zJ4Qsbj8dgeqbV81WuLEHD
g9cbYblUL92SFhcbJOENT9r1QmCfrypBRwL+pQdoDETv3ajva5RA2poW/b5A2pYw
zi/PgpcELEWUWJ8QfQPI8w6DzLmWPyloii9eiHxV6FohOe2Y6rLhkgQuIBPOrgF0
3oLkwa/UnM6+mHM1fzZiXQuMh8RmOOrWnR06yBM2RHwoP1cRNOK+zZuEe/JcAPQQ
MfY2mxW2CB7KNtCPr8F/qPY7B/GhIPPz6UEUO7BVhTtMtntsLHBnigwIhxBq3pJC
xkxO/ZPEn4P1IeQwFIls++Gu6F52W7lsrAhJh3CJi7dY7Tx2XNWtqGDh+PtJJrB+
aQFRvQ62ey7/Zz+YaKGqOgR4gAKVSa/Zvz81tJet5WOETzJnuWKlslfLmdtSrOG8
sCtRTlagnk+79Razfyc+SGve5QEh/aTkNMRjnUs+OeeTZmD4Av5KRGXZPRWP8UGb
+/SBQRjxfqziNpXMtV9RWjUFkg/K4VcoO5F5RLQNjvHs32eJQcp9CriAYIKvZEIE
fjzkxag+P9EN4H5RUYl8EBGbPOqVHYH6WNYAKWmMFT6cMz4qJ6ULl0OJFEgSYBQd
OYah0152muIjjYqpWCrrNv9YRYXBe1Cd5MOsmJvW/mwJxIiR24nNr6aGUTpOgpsV
jvERBGYctSYy+lwakme/lM+Xny0UKJz4PBNtmPGJKsN0Ee+TSLoQvG1JeUOF9VWf
DX0QEMgakzzq078jl0hPiWu6jo5o1Fnq+SZ09ejJu0vkqeVKc6QtzRVnx9K+0UAv
sJVb5iKbBkqrj/gpOx8ykqwlfKDSp+9fPMNSH3B3/ypWlXIWJgck/wFS9E6895on
gr011ywYpsZqxxotXpKD+eWtXnGYgR/Fo2JPEBqwVRYh3RdUnPCqnIbkLwNWzlFW
L9tUmGDiZQ5dBtYSi1lRtCjnkNstrqqsVm+faOABclYB4SNRKhqD6ZQHlJCeAvZR
6qXxxt1VmMVRuU9fhE1BnMp2OBU/8vPrw8Nt4LwXkzZWTO4JROjjsp2hPQwACFQW
rkdtn8+DiVj0QSGYciIw0WpYb+2zdlrbdilifnpx8NO/5nDtLvbqU6jIGruRYQc+
xE8firMUrarQLA68uorM/2lLpxImF15PBwoi8+H52KnCdukfZHrfSAjyRy+jpvKj
2k7d/zrFmIGXvhZMfIcK4J1YMi3qmwFIysqsPOVdhgNFUx19HShFpCsYVLRQ0NaX
laDz6chEeogKxR6yT+E2qX8VDa8Lgn9lvnNubltjCh1a8GvBic4m0JSHX//X/scy
btyEgZeVdTA4uMbScJ9OKXPi0IYZ7vgf7kwLS0PSB6N46WTFgrPa2XLBEF7kh/mE
26dioOwFPmt8UxZfRWqOHR0NQRFMBgsv/9KMR34Su9FjWnSdFDTFyjGZuSmxmVCn
UduCJZ471HBoRy0x9Ty87bblyjKY6s9Vo6rZPOSq8soZXgzpgm2x1+wkWbvf6rNk
QeNGY4cX9REh2I0r6LXGuJtXmPP0fMaps9Uzgq4zQLh1NfIi8fl8Gy6Qh6nwY0Gf
bz87emVvmmFKFJBNyHdVoTM5XJr4/QDVWVZSI4ZYpB0MaXf6jCB128QA7dTnRpyG
f9J2zK+m5MxK/k3oPHi5ye6tOkFJ2A02kXVKYIc9qqDmT2YCshrPh5HO3ENThHS1
Gb7kkzIxMcIlCDN1ZJKbhP1BmBUECghHjTBM4n351e5uB5w7XSLmayhMVcyBKn0q
jwMWpViXEZKK+bBdqxLISu3CQ1PyL7OD/G6shtkW35XA49jbvfVOWE374yFOKIiY
VH6fTgsK20mQIYOblqjgW0BiPTMjNPMb5OPuAPGUoqpqZCSK537eIzCvzJSTGSVw
LNIXSpOVoTcY8F7ou0oD4+h+Lr18dWHtn3ea5uz7aTiQzD1aVCPiz6AQ5yFed6Le
UgbMWs5FxzcGneEuN/5VIe1URYCPGhkIqFp7/Iw7AzXTD/1/qgtBylTU2YAszUk0
oJwKWBZzHS8Ywb8ebPUnbQkneaugglTAHwfSM+/riOrYSEWw39dA6CkZbp3lypQG
A/AldVrOzvKCGyTVKGbAbE4fLj+UjjG0zlLQHaiDpBO3sJM9+sSQRTk8cKS5L1zY
VH6LC4yLG6+UEmvpmNEY7vMXwbMRP3dOwnwtj9ljHeRdxbzBsQeXslRZK8SHv2b8
6gzfOzDPDemApWirnPqTpkOQlWPr5Vy1SFFUvOZLsr83ATHeacO2+6SGiul4ag1X
RwTmYZZkUQv9MguCWyEY3r6xbdDH8RVbMIy+eGgs62KHHs5nNijnujsrRBYwteFl
xxG4TFhaAIYD08ENMReMx8nQFaL0M7BYam2uqEGJfqyMkVY3p9Bdi1kZ+CCKgeGW
vFfnDrNh12jt0apNCI57ts2eIB9uh2OJ8TzeAyx1/4XRs2lSLac9ab9Is/gUyXKb
MdBWngzSBFU4Mv/x8W3q5jLMczAwuj+p+lW2Q+yQkjAPqwKY9bjw0Ty4VEjBmvE6
M6gkOWrEtXxueHo7C+JXJXYctpuAqVMNaCvgiYXLQxgUgy8dLzvgROTFvpKVIrir
P0EbOYzqtCVNyBY4iGueOnDDSEn6nmfE2leMjWoQVIM7rawRggQbpl2DrAhwHv8C
rpIC6srUVh4tbnUg/IfeiSSgwcRHuNGn8xlTz5KHE8zrEQkobsn59i1etzKZ9G+k
4vNWTFg/k65cwpUW4pa0cL7lwnSSedrBaM8VnsTr7ZkdRmdMD5VkbwXlZqJ3bsB/
K9up0jJ3Tv4b3qf7dGcy9n/WlH0bW1r5bAtxsAralNdThxhY2seG2i2Ka+V9IrBA
yWhwrPpJR3Cu9OrwHbl6AdAoKQ3QijD2O4pIy4wSr2fEWYTslQLEDBu4HGRRoXxu
yxwmGQKsDebV5/bC5sUkUP9y2Ncj26vuw5upIwVqc9USb9okJ1BvUkAJeeG48Uxh
llJzEIPdKBbS+sONxHWk7Cgvw9KFLcMRr/bQHGp3a023Vb7T5brbCQdXtC+qUsqQ
75VIjukRFkCJ96FmmaZev9mWbgnGQ+3AhaWqDiVcjzENVCesh1Qo7U0OtZ152pgi
WV5fSNRyBn+hOv46lrM+PPSmZGXFI3reBIdVPe5q3Xw7N2Wq6kgzFyqVhq9owX1h
3dgubCZG6RKJtKa8YaQDJ7aKRBYcMosa+6WNSomeX8tT06RZvVgqJ1dvvLaHDKX3
3/X1Y8oaTUJd10ePrpoxDPs4yMqAFFR54SPKNenpNpGQiH9oic/rvkDkl+XN3ViV
fhd6VFbdu61bBH9gKP4XhQV65B8D2oyXcbYWSZhEciTHsnJ+Ev6t5e4zXUdaQERO
NiW1QAi93HRm+2xyHQgT2/her/gw5J7b+DVa2Gf66oo/+njrjKcVknHh4oEFVs3J
eQCVPvpvvAYhWbhaL4c3UGwMtBuzUXn9yKISbdKmbiDdb2XqGeQFNeAG4y0Lw35p
feh9Q3CuifUiSxkKkIuNB8+/GUnnabWe2rogOFDIFKqcv/FG1smSK8d7Yz5/eS2N
L/zx34B7EQwcGU9m27QnHHY57Gt3Sh2Ms3Tc5pq8Xh03ZIVfyC0DjvueV1m98760
JHLCi2ORSxk1nM1+1vMQcveYob4RjHVuVjMv80MLA+1HD1U/f6F+mht0bsk5dk4j
S+Ma8P2gTSedoEbU8gWwS5MwArIeBWZ2pTN5pQd+XOnudZxcGEyA3VUcts0XRhsU
ZQJ7X7+lj12pgszg/T6jONW/S9BPWzdqoKKlI9MU/1AUkfSCeVaAGtnLpuDP1wuN
bngHvVwgF5gCs5omHef2PJOGbqDbOf+7pMTK9KkA37nUvjcQ3ra/nUiBvkXBu3/x
0Go0Psm1iCjzGhUJMulYloUqbOCQk+/Oy+pqUVUREoLQYiAvdNaxn6Yzj3WJcbm+
BviLe8Yi2ssrvHTSFe5p3evD+wtrkZNf2gLVSaXdo4Nc/bp5FrhB/QB3gbsDZimQ
fujNFdVBd576SCKZxg8nxHXGiFT3PVSkB5Bbg+K3uKJ/cwnE7d1H+V0ioMX/6Kcl
JfkGV9ePS/SSkJPxTN8QaG9JLIJEu2QbJPCHsGWgI7CM8GZzy8kuRCl6zf/yzRsr
mvSndsrZLcRKeY+tCWeGPdZSjV+BksR3G63RntxofYKdsCxl1/n0HW1vMr5WSoyX
rO8EZoGAmtKwmuiEt3DXgFCO8i1vcUDg1xiU8/2ARKQxzD8t872/67P3XbxnzPvh
BTdJm340Bf6dWX8mahp+U2etZkELAf4vCzXIwrc6LeivfT0WohUY9blcby6YxUjm
1tyBSvW+XrNybPETClQFpJAJb3oEjxQahjg8NGjzX807qHN2ZKApNLqTFn8EZ3hm
t9ftLfesiXOxYFd8iYzXmO/4nA2PUwuhkQSZ/goEgCFimF7PljjoFsKkqWoeIp1o
Y/YTOF4ZQIna1KNu3/YP7gQYotWJRgvKNZOkBBuOUTgAggVB+gkGWxB2Vz2AwXUx
cuHECn3+9XSRPKnppaeKUPcAt9ier+NOrJWxPMsWRnYX6hg9sRCYxLvIvuVylXXt
dYuzVZhboVI94NP8wdn4hzslfoxSJmmN1j3GLf+v1HtRGraJt3aJlhgsU/0toG4V
Z5iHudwicXTcMW+4h2TTBv1nrdRSnEA8jQDO6CwF/g5yeqUYwkKiLhLkTg+fK/Wj
b7CIjMYLf3SwPi1Vzn7rJShuOhThfWIMnmsrS1QOa+DCFOQZzxD85U2NsOMw1sJw
01TbPh+MaBx6uB/QAVp7GG8RXKKgkHeo2Jf8cCWVWZw4iLNMok5XprNheDw4BuVb
bKjdCqukWPduFIZsaVFp7eQQyKu5s70EsHvwui1c19AmMiPKHTrWF8h7KMf6FzlU
O+0yyce9oy8sWf/fKnbeo0XDqxOwRpwTPZnwly1yRPXnbLhaJRhtSCLHJtY8n1xZ
Hluud/8spN3516+ojN4aSrTBNtiUs5Orq/0uJmPIPGi5wUe08fxoU3Op6xrpKQgs
gv96r4keb43KheBJ0C3AgdpYQyU9no86XBI9PYgk2R9qJ5bJBoPIMdpk/4QU4/gK
jeXjKBsLudEzMRJhXNMkPPqdgWOi/lQ1QVNoQd5ieUCrnjL3o2UOrIhed0VVrnmg
QP1QDv6MqvV2BTWcL/xltq6YieT4NE8tnPhD4j9aG3WS8ATnm5zwd/ALvh/mVLFS
mynCfHSaD7+kuiLkTB4JNHYKeq4dmwN+kS6Pis1gaX9m6jtyU/4pbpG7Myxg4OWa
rEcdLoUrEQsKK7rNgZdmeboKrrTd80fWzvxV96hj4Dxov5fX9UNpUByDnf/WtSZ+
9eyNIyxQzRkE5GotYSrAqRUUFFF30Npo2qKKUuhVR2luthcWBHpVW8cYX8FwBbWQ
X5wPlkpY3sr5XPZsUik1DaIJGsioc1uCfMn/mOIs1dRBwNxenTzAqUvfB0CkKTST
O2Qpdm6sYxjJSLJNEPtEoUpvqrNVoT7uz6f4CyEuVsp2tIfuvlAmBN10hcdRnD6E
4Wq7TRjmoIbSJlN/KEFCtGf4cSt/+aW/WBDhrsxIbbyJKEKkq5OepiXBdWB575bo
7GjQ14Z8iUB0ZwtRzl+BavJCw9xENApZ4U+MHgX51VEafHvF2sRKjrT+IfTyG1Kh
Sid+3vwILGjjNZUZZFXaNThHPRXzFwHtDBwYp4MMQNKfpSO2LN5L2gd43JSLRi32
D8eUlY2N8OdOpFgzfGgKnAMnjKZUDzmK15vYQNW/La6bxv/jzq2gWmFpWaMmk3Oi
HdYJ35Mn519iopgG5HhfUadIzGGKzHeguEg2N5wCbvowDK0s+tMaYySZRNDxRCtJ
tvv5uL2q6ykTWSycsDjz7XPNtjMtvrkUU41PCNEuqPPCqslHguD4Phk0WKG9BoFW
jPvKVqLyBvls4dMGGsQdcaBFyz5s/ZbCK8Jd7l+Iia1KwsY2DZerC4UTMcJ5UU2Y
2mOtl0maRvHGT4+WvXjfokGrAH2cYPrytqdz7iPsCpInxkUaGwPfVBUCx04KqoLk
nSMhi4lGfpDvMVmHiPLzg5xy7S1rfyXqMBON8/D9Wdg1LwagL5WkEBg6KwoTLihN
vB9kGgtQqoe1Il2x32zxuJem2xugCzMwlnEM/WOWF+gT45kA2witebiq9eyvyN3q
dh+RfU/LSlBz4qXnLRF9XXtqBu9e5/TkU16t0k0t4qmWfFWY7vJyC77dOwcapjWn
txdOL5NY4JVZu8s0A8yLl5kE/efEMV8iAssuRfXqURH/WsF6LCAFGQk42rrKwuEF
sKk7asVN7+sClaAFZK2v16EnPyqkRbUlQcV+GUximkZw+I8WP7cJkhc5OCnl9SfW
USGdsV9xQQf3RgL9QoJqQOCDeshdkZLcickcjiMfojYcutcxldb2uGI1VkPFqlZS
nfBqjQbcPfHVG/lL5nyCpLBMyIMo4y0AXI5PLCwaT56qfjDCSDLOWMqCKhfOTFOh
O7Gf49XAK4WKa9t7mRo9Et9uMYxCTW6Kw3v4tb4cddAvBvN+eWk0yYdtNcAphv4w
I8hda0eSRZXViAOjYcejkUnHExv5LdU0HTrBaBwT2KlT4yRFabJ6Cj7FuwFn1IWl
f1kiFmKpGIaR5EX8q8/y4PlkdXzPOPvVb6joxcU3UGkEwXfGOYs74IyA8VATig4X
r8oc9XhmW1QTbw49R3WQ+5APHzNJ+HH0OWqkwmXN2Ohh+YtY9jVw14QKtKmKICJc
Imu7l7Wu1LFV8xW3YoQYeOJmUWoX6nVeagQy6RX+iCVTWUBZrNrJV7ktXeHutuvO
52t+QJruXpZWhAlQNI7xeVJIoEr5EwKpTVLqe2og+u1SJJUbF1KvcYguQHc0RZtq
lG0Z9VyWfRM/bUzB/N33en1xlvhhdJzZvZOdVCOHFWl3Bk+jWcTUkhxsay+ZoOKc
Tysm0k6heXWFWnS1NefKfbOGHsW9evwQrwesQpFmGQ+ncKXdLa0RpX2ueIlbwpkn
CoXFNBfVX2BdOaSljtuEUfhDotQD2t6lzGvcOnWDslI5Yu75MQqH+pdM0UkBkQc8
sONGc2/+2QyZ4GQjMHeuBJuUGNNa8UPjh3QLOEH794CSBJaG9k21rM+29xXIqVch
5Im4gtm7Bq6d1VqVYFdA+GA5H+NvOjZ1VhKbrdeiJ4W/ybOARGUBPOzQdIFzbpv0
1p5dt08jpP0rUo6HsjhMhAbpFWwKbt9uS48SFIwuJm2ONn4VvJvtDAmZknGvWsLA
CvC4Vy/Q0yWs0errYyQp2XbkOWFA1dv/mD02k+lwd56P/ntUQlcZQZ1TWJaPV7Tw
y5lpVeE1vgmAXYRI6c1762VvL9vA5rcbYsg7iXWrDpyPfQG/2k+NszualE3iv8e0
whIlDEMKNR2btKE+WxpeM+a8BNaeXulDcPY24iCj5YE74ZFw+oS+TX6heOjL7cSV
6Vex7UQuMehiyqoWzMbmjSJq/27jcvhsYMpTFxNGEBUQ6TjBFgA0vxVIOhAF/D8Z
sfivkhCo6CiSVTNj+8/ZU/fFR7SGb8vtvW/gntEwoIz7n/hoTAijttakiusg0CXL
TM6+wteU9LYovFtYBwEmfJaWLZcMX3sYGZ5urwsCrX8yYNcUnNSrn+U5vD2+2y/b
Wi0X7lO7Ll2Wu2TvbvEBApO3M4GRT6UATBW7kZij9gPCfT+u9Uxj/9ot/uWvYGbA
XGr1zP6c9BMyv7T+xY3UDTokCenAgqf+3gl0TcJrsUQB6OasT6FgtPr9jBbWSk6k
Zk6Fi4M5XB/Nuv4unD/CrEVv4ZyKmGV8AFT2mdMCV6I7UDBGm6jfFuzX/5B7mJ+h
g6VrtkbqDMFFkhSwWCNqjCdOAjrEDwhUO+CuCP8XXAhWPgYWK4n77SJ8ucpyAC9o
LTogMHcLlnIG2w6kUxTFPVrsqLZUFgLaPP+1fE45kS5xWqWvfJn0/U2QuZLLfKcq
KYTFPD6T83qtKWw3TvSa6MhBrjAtB3Y81rk38i4M6Ur/kmAbllwXXgIMiBRCD7Hu
0L/ukMWxRmDgxTUhwhugdKU1lXD8cTaEJV+BvJ9pYTvFKEBPCsrX3xwbs17Zx4vf
JiOIXJ3R/NtsOIWi58At+ajFrgGS6FozKJ2edUBr60P5VNYYTuQOIk3ezYMuIG0r
Y1LxNnvwPEw9FctMZcIRhkL+H1uZG8D7kbO26Y+uFJMLbsHUh5tnjFZltXQ1ZabQ
7nuCG4tyOy36fY4rvRq/ehHOk63HfLRzNQLMteEmnhA57ELMrVqVt6l6MB56enzc
hKWhLgZgB7SBVM/T4ZjTMZ6wVjvbWScGZu8abvDOgTCor5oG0AekpP+jktTOd+3P
3JJ2ZnH6L0gnznbKZ4r51mUvBod7rEzCd+MaisrOO58wn68SciRa38mZ0AGUoj6A
8bThz3GSZwIQnBFTpfp/amIa43zcC48cUx7CrV8h6QrVD+fsHKBS1lwGfBbQjlJ2
RQjOhsJ6rInnt+Ci6Zd2V1hdIoB96QZV2cfMJ7wjHHiwy4kpEnX/KNk40hDm4xBy
9oMXbSNW90w1TsGlVzbiqXpYJNCVoWdyS+PifcL79TX0knpbOIzLTo+LrCP23ddj
VhDcbNriUyPOVTnbim18GA+tLPlR/GFtIDcGGfexyhh5N6CVBWd3U1K6EQexxmmj
P3ADt5QwQu3J2vqMI52EoGBCjmwXNt2IONhZ/VfdvlFhadrYDPd+F8zgPPv2v+Je
riMNyirKeDkucqKdxnVtOBmEhsakDWUS0lpN5EfS3NL3HRt6XjcgRv2mDz2V/KkN
g8+VuTSgDMvC73O1yFppG9Mq4IX877yqcEuCzU1entAsgYu8OmWiE7U9qsocavcu
R05bds8g+TKutFXDl+tw4QcZJFerTnxhu7pDMWT89ZRrVqtLbnUPcpbsi2GxhVwU
Iz+6Qai1C0MhKTqPoZRSNDR8YUvwEvRA9SI7Lxohlr1X3XnzDa8wyTnP7qF9gEYf
jGZUAcb2l6eYbvlbqXEbyuFINo7swDI7OvmWYNFgR1Zqqy8FxJCfwJ0zDqHfRlzC
kYtPJrM9+yCZt+a+pCVe1EudBjhYgQef7dho12CaCoQ/XuEVyyhEN2ch2erYlpb6
23HuqxZL2pJL+IvW4UQciOMnv2lhyoNj30P5ur60hQg2kNim7VGYXVS9bIY5RRHl
nxPwe0ZSQ3Fa4EPo7SZqc/J9nnJuu5r/lz7oQYlFsMdFA/ErZRpXGfHD7/dXb843
qrhR3+yHbesulbkU/WxJfaMYbiLJ5hnckquAHQWJcm9uEfmNFdt5LeC/Wpq5GauH
Mw8QW4KdqTyAgLmwj3QsfjQOGFuDA1c8K59UY5aCz5yWc0n9Iu+3u50We4G3nmTM
aRTXDABX6BZGMiPcYa07upbe4PP+xAG+lMppqJJtEV0Qj4Zu4W58bFsikvpqwASQ
8ai6lMIcL59NgWlJGgpr19YFx8XZetpvcjE5NTZFewwjBERxiTtuGeBYHedVxc6D
X1smTdNQ2LQUoIW4mEnMN7O5zEiTyTibiFkAk60oIE+G5rOEp1XPRqWp3d8LVB2w
hj+SVjUrKaXnDR80YfeEFs48JI6NAYwHj5mPpWEw8pGQpL42fLrYPFP0UZlQZ68t
wPiMjHYAb7h9lMkAhjsO3jCWP4moqI1vNo2rcAzb5VG2Ip5vRKP583gO86NLSihq
2qkXc90OfshNT2mljBoVcfYlRpczh5QLaWgF4Y2M3qe5UbYjtPrku96mJNNrO6/0
yhWUwp1G/9NLLfVXPMRNshQ9M7cLWD03IX8N/DIiQsXMMs3DLNqx9x1VgsBnbPue
ajWuEMfdMEzLU6bYFeW2xE8Mrb1ywBcf2Oi0NdVR2R06mjNnEbSmhxAvApFmIY/f
AdCwXj/C+IZrL0wmrBzNDSFQiL73+LN0sbQAJ3sOXNaTpfe4yxL95MnOvTLQH/+A
2RLtoD/zRackQ85j7loSrwHGXXlHQ8ubfKUUGNL022lPto/RcXqZBdu1e767QF+Q
HJ6wE+QotdRNYnF1QeKvzswMxUWV7Yay+B4EVmNr+VV1BeEM4QQSacp8QpdA7FcM
7tZBDqQHXrVA7zfOM+qpKnkYpBd8Vw8hD4lsx68W+Lz86NkN01PGg35npwv05nOP
Ojd+DORdgIN+O2LAC87HfX9FU3BPvReG2daSeV3QiOkH02o1NKSCIg9kY/cbu+7x
lFK5fwpRcH3ZVosfCUjObVPd50qdQcNylc4CEXNVUBcGgYpKSQ1HmvfjyBpIpn/j
/zIbKYMeWU6QCQ6UaRXVLxucPy351S0/1D63V0UgvRn7hqkyQvc7DwRrd3aet45D
eCOGupeb1OJJwoIxjYAcFy0/6AXJYcrp8Y+Ong4K3Ljy/8tRkuSBTpm3uy1Ghaby
xTwckBjja6xrOT8GF9782JuM1dOPMUSlSa9acY9UlYptVon2gX0Zyfq/J6pJ6Qgq
cK9AmRflAtfYGguuK1gc1YDN+YPq24oAkb/nmF5gCOveDcTvZEj4qnqL7Oe473O/
BAGF2oiKSJf8fwHRL74EaKU3jWO0YTOHnoy3rNLHRxxF0IEb6ozwJSX7jVV2ZlBX
y9l4W4kurDqj0/uDGEwoPVTL6ml0FT4KyU7oR74vhgi8Av2K9933HYK3QfrJ0D6v
i5S3B2mc/ZoukE5/JXcFhBWITwJNm3Rw918q+AcnNUIvgA4vgSANxeLL3qK61/Mi
DQ25HXD+dulKya4DZxRqAxHdWYtaK8GbC0fyaLxZDhXtRWf05JRJPWV1gGsTuHpl
mf5gOmzltPjH/NkxteaQGRxK7dBu9mHhdaIaz4CO3pfbVY8WWoqo5yPvUDMHKYKx
pr4X6CvNKOR2/7SxuT8P1J4E1XToV80XJ1yuYhHqGI5fDkZ1DILx5fi3fokjYGdD
bTdxGHV612Ry19gVgjkgYwLS4s4Cb5PowQRvEpRa2JR6wB6J61K6ryhLwlrFy6lC
eK0AChGuDp3O4ZWwFJUFeMCkvcABBHXAi1x+tWFW8NrhZm8Y4X3PvpiOYMn1+B1G
O0SriYRH7j5gQThrxGzAYj9GV8yWzO1w7KIp8kU4nmdUj+lBuL2fknM3VG+V2DGz
jc+vBENIH5eq1SCXOfoxSXZ5PbOxXz+pTuya/rp+K7PDaINKiCmZmd8erb0QjVXB
wBk+CNicETxujQdqIUoDpS1VoIz5SNHN8DXrJf+PSA1T7dnCncsmtCA9FRJkPomu
WURilKI4afdtp8ddfW80/rztGC/2Y1J05Of7XijFDLYa1MwqloJIGyn6GxxGk4K+
eUJEf5xrnrgzh5sEXBKlShfXDPCKERYvsydsMWLhmKbDX0FG5cifozdjfiYjO++s
ZmK9/bes/aP6Rm21WN/eLRXtgGBZQYvWMbJG61YMwGaSjg+rUIHE0ilIXq3NstfD
4kg0/EIF52Vr1cOx10KN8k2+AMjiaXIxPjCtTLfXj2cEZj42Z9GZ5GGs72rKeEBR
MxHC1kbm6Iq+Qx85QJn5gaTdHytMpYSNXe/nnCtyCON+cie8ssTHPnHca/pNeSr+
Dbia3MBTMVmSYZ9IWwR8AROQ+8WRDCIK4v4LP/YeIYvfkurE4ID1AabpS4ihs9Pu
ANjXF8tQE9mxK/BK9ps6KYRwh5+j2OUP/u0VbaMKgqGCeIowSaRxCBfD6zzRkRpT
H6mcE0mEMpwA/rOqOOGoVdM3l+n334mCdqKUAzrE2UczO8m3gUjBFeRTfcpBMQxo
rAUulQiMIIlKNF2YVVY2B6fArk5iuN/GWiy+9lu/4ebMp2qhyskZNSP8IXc/ED3u
E/ZurzUu83M08UmyF33VeOxjIAF4/uldQYRrjRVvLsXrdqXr/0ZN/ygd03BnhRvL
dm3Kub8J60kGuIrWR9b9nzDoWcwvEgYyFQqfUGYhyzlotrEyryBw6vQSCn9JMUQu
KVOTj2I3t3OG+2HSodwCYNPm8fsuRUk2ywSJGk1v6jqukuz3uK6sBb5zTZ3w7aGl
ndO2CmZ5a6hTHc3UgvyBN4vbkqmEwMGTHxcy+ZGa661V3vx5+Z/PHiegV5ZO+9AK
Vm414lcTj47Z5GAIUpj+CQMFyBnazml8Qdk54JkTiPY2LlR4QQY3j8gK4gezLGba
mWaPZAFNhgjGHRHQzvI0SeYmCwjELGf9oOuFbnM8Yjx1XjINt6RotDh74j4fVmQo
wMf8fMqHxCNwDSswPJG5SXKRWC/T1jOqg2jnlhKc5qRPGGu4AaJSfw2S7jFIdql1
ZzhGEqZme7dvvNB3XqNcw31iF+3YHrBS/+VPMJhxnYTxtVI4vEy7Xy87EiSnDqFf
8+a5PkJ0oJxvGt/yQ4nEigx1vtFc5UPLnx9eYGeEt9SSY2vEghs7Two8QMBJ6UYG
5sX8JmGmL5hoVrQjt7lqJV9cDurnqnkprM6g7q39xeMYM5utDC3KpxmSQDCJg5y8
PKEWpDzRrMf1mNvUmHSBK1zuDhUSBA1cKsDGSSfMyrh3HJZhkds2bS7cbp0zQ96B
UqG5iEq6Lh10FSmW+I3+PVHRH7RBpsUwBeoewesmAxr1hH9uctVVQgWF/IMvl0Wt
wZQmVqjlRILNatb+f/yjMAzmRd2WwV39dyHuXTXln7W62XnVp4b4CQmZ+wNq5nVT
veL96egSFp/G3Z/snBtLKpblTWadpZz7CadtgzAuP/MbQsodHUGAV8sL3nisjHdV
qQvu/wNJaQi0tfxo0UANffcdCHf6aMVF9D3lNg0Npb+9qILTxT8zuFFSrAN5NlSz
LCpLcN9XmBqeAxkj1A/JMexZtpUbsfj5Ay+BZYz2KxHXrcs30cyYbiPtqN2XsS5x
RS1BJdDIsmu+ZwqZbIG8WdpKhoNtOq7JL6T9Um2jy2ZwNnriavG5E/qVl7rikGph
VGA0E7oHaxMGBfP8WbQIhsRQmHmpYteodk9WuXBOMwtcPm0h/eDXHhxKKHe5+dxp
kBdr5MFMXEWIcTgKBBehCiDf9uQafTHF+OD5esZkM4pwheieV1IbwUZ2/vMFxx3z
xyO8ou1ZBgOPTrN2JV6GejJ/nb2yAIslgD1HPALbRMyYmA7qRj5qlL2X6a7gOiv3
WEyWkLg4372l5GfPQvtaZQ2SiINF+I1Ogmc5dZzp7pD25RRCK0UVc9dACsezbTzs
EpFpUfQIQ99CIvGX7YcGk/28XQhGQvV3TLM6J/scwajv9i4v8pGnKZnaXZrIJSCx
ue6OOIE6CCYTNZIx0k+bpen3eGPAy0sG3kQcbm99ZD811fdXv4buLEwV3QFeuXwk
f6TkqfqIT1tEGJPZlCWcrOfN0aI+5Uj0itU67eFwObWSmUJYVdsePmq/6zGU5u/h
mxO+22nFWATHi36D8ZnzoifbGN1IomFtAX9HFajvBRyy7oRvMaExSCPM3x+FfJsW
2NYKArSPG4/SWyEZLJwqrD61YZqonDwM1YGXo9n3iBRsubPi02g2zdnGy2hCg801
kt7D/RchhvTMNTHebqCQfRgaFuvt02NBePG4L1RTjaIG8KibELhvPsXxYTHMsIqX
kj7Nz+bkljrlvID8w5YrXsFxOzWuh3q5qwVcN+XbJ4L/YEfcKdhyIg1vesAYPpie
diIx7/G8Q+fmaYq3K6ArvaG74QtNlyjrhjfs7/nJgthLqkLatNIoFTsiofizRmCA
6p4Ao/L9wHyG7GQkBhUZiSY+4LmWNW0Btt4TnoEpPPOZf/m5cqgDLL2NCsCKHd7R
ngO9XLx4iJvyk/dDcILYxim5Ch8nPQUqcKj68Le2ogCb5CUqXFEbQO26S/1cw7a5
L9WZFuMfbFzVCPnrUFogb0GruUyp7u5I3yPr9Gslu1vjUBy0WQMMsAT60YdKBrvZ
mC+CrnD4LhpzQKSIsrV5BzMR4CvID1/PD3nGywOaYi927z3BGW112RtywkwKvKQl
D0ol++MrOh0aFq92Bk/fjPskFL0bEQh1KkROjaM5l0tKnzOpfhHGXnStQt/NZrSh
OjEpCR9MswkBf0i6R4T0kMQF3sersUz5qSShQcyFIi8ziKfdbTTYP4uhFGCDc6rD
jUPNreGdh7Hs7PB2tfrASaJZmBuV/+qWmLgOuDPxLUuRES9P0IFpTXprBilCG3xo
gbEL+rNPAW+6M8xM6LIEGBvfX3zEZOafBQDEKkB7deAyua2bWhXBIhCoZ/G3EWTm
H33qZfRDpgVcmrvNLCekfESTzEIfvKt/vWXgSUUDMJoAVWCc+AH5iBzg+CsMpfoS
zgFyed7d6poIviO64SeiZ20fFxVH8E+Yzh4dDrjg4e3hReswRza/Ls19Gvm4+D8q
msR5SSO9a9W4EtBZxf7ZJsYhVEeSO3F5dkL7s7TRLgUYFDvYksIFpqx99q5nt7m/
MHzEHRoVdI8Q41Tdbkn5uhxiGXZC1F4bQ4iK+Vr9L6n4PCSz8JkTTvIHEefmgHBS
y9H/5ckaSXMw1A1Ymy+A4PeljRKkaj2A4/GnrItoy6tOgZl3ywrqtlNFGgKbbT0c
qri310WV9SnIyn6UR7DtyRY35Sp9BQuI5CYzEw9LN/rs5KPMSm8EoA9qIBmyW7OL
t6H4xNdYYFD7r+ng9B7uvIXWoMG7fi4+m73eok5BLAPcXDRZwkq7CGEbv6buh1Bg
Dt3sNMi0h0EzvZ49PGGpjk+cbpo6HibWi77a8tK8xOqGpI3e7pufvWXB0yt3LTtH
qujxybTCtceUfOD4X2q08Dex1S2FoFaXOs0duLRqaCckmbe+5GiaCyE/+tK9MPAP
fm/NKZix6M9qeu2oBqbcnDJrQDaPWiq1mYFGNK00yIm7mstZdcPA7JbeoM363L0m
oToLHOuChFWVqHclwly/zSax3Rf+fduDM1H+dGHSp0x/Jtdq4+LUARizzA9Gd0nc
i4vfYhlP/ubPwdJIJzB2plOO8H1JRwG72hdrI4ryxC/w2GsNOh5zqP0PzUvM50Ti
/SlJ65TLh/WNKU3IeasJIFlOtRB/7WapX47Lk/85i9EjwUDgSJKW8uIHrtZfr/rO
kz4eCinUZLfOTDUWfSrq5FPjZ87hmgjkqOrNF/G+DpNkDvjEBIfTVwMrisP/PV2S
iNUk/tTDpNQ9BFSObeE1NDoFBrBvdvUCjTIYWYr8fj4keQsUi2z0Gf8r9BPdMHvU
o+HReKwGIu85yVjeHfxnttopRnPUpYLaTw43+Mjky9zNN2x9WJ7M6w/Y0Sb0NPo4
TEPhmZlxiax2Wmxnd6zDF8ZeTjaHTixS+gpebN0TB7v+W11/HgRQrBmx9fdrOR51
6p8NQLEZP7iErTZL1ihL/KnY2IH1ahsaUDfdDA9QtAUSQrJmnSIOF5hzD/HHOlPl
2hDIvOhnxKCX9ZOQXglan458XeIfM0t4XcvXyog2lrvfWo3hXx3H2PDfrLmlcnuZ
OjcnNsn3m0xRwyVm+nx7HitFYDsgpMycRaHI2TtHFlLwFNMXTkHk5mLeHUXF7lkv
tei8jiKhybq9rpF6LpjQ2kSynJ08xn7qMHS2RuSUCxug7C3Q4OzXdcvQq0rbEqEh
uvJUmnAXHDmProfRjGBNVzcd3fQndiseIUn3QUJ2eH5Wh88wJW9x2gjZrtsDc/DA
0iOPMsgqK7thtCCMD5SWdk325iWA72Ilt1R0WcrPlZlwka8QIlPj7W27JutFWCkg
y2GwyDlHE6uAg/L5vcLK5SwzFmlMbvl5Ayi453TCd7yULsdqZH+A0Ehg6k8IxiIC
tD0MNj83uh3FgZ/fpXudjQa3n9VbIRDpLU8dcw9PQvKVAnuLZcZ1GnozecRHalp7
M500K81QDMohj7qgeKJi/CnpdUmivXx0PGgEkkDs8tT8MeoiiCMvp+KCi8u+o3pq
NBTOcVfW+/rJ9G/5NcCDReLKAJfWK9VXBJ68kZl7m438Fq5DVuf/fKB0et9nyxYE
2g1w4MG3q9bKErKXBWaUvBFFBDPhCumVTXAeJK8zVtjJ6l0wjs9kC6x37yvCoQ1G
YAf6lJoMc8HkcEx8QNxNsVH43hJ7G5xqZgQzAKpDUgTFrZS67N8Yh5kXkGtu4okH
3YM2hmBRsERBMziN3Qnsf3t62WGRwe5vu5ze7BGO6j5ddz+e9PytgZW0jj1fTbVu
jMkvWDJiZmpB0JuBAfJmVxFcb5m0/hclLJ7lICIcASgC0MiR+/r0n/32Gdpwf7EF
IoQfugdWtmzUFSSbsnLJ28Oj5uhcreFidynH50TJ9AS9z85QfjibUzt6tAJJJgJ5
WXb4OXP/nYt3CdaZJt/u1u1XEsNMJsuvZ6ukZ6itELmdVgV/y59UdgEruIbidDda
p794NoaVaq5pHwR0GdQ0dx5aOTm0om7O3VEJKZ+OYwYKM73v4k+YF/6DIOClgKIz
NEgOqEvvjzlSLYSjN5F+9ABJYOj4k5Vki0H8q4nvJ8S1c5tX1oq0vlucrG6J/9EX
Q/j/wB5T6L1excvPNP/kIVaC9OyBmprfut/ONhpt5bIey5kTlug+OFIBnlu/rxP+
z8KAjUYwHUOhzz/3XNbpLxj7q3KS1g5maSDPy3v2Q859ycfO6Ru1er4k/LzpiUxU
+SPd7EU8TSkmZ4NfAxQOWHyInqt1wZVPtL8tq4KTm334iSJnzmFfdTl/edzByW1C
xRJ4Vw2adESRimb61bDhN2zTUP0+jbLveCWT2cXUqP3C8bvW0346uVdnaDkXhBJM
1dBiI4IJx+QNYK3PQuYfnLFwDpYQijjKbAI2puv0Ku7t0NPUIXcRpkK61H5VWs00
OAVAScOqOkB1gi8/iM30ajPuGNYuyGMEK1tVJPiHQmBksG0FJuu0/DVyuQ+1Xt3r
Fb2JmSJPvBMZsrUSwEBj19febbM8EeK0JFSwdvSksFh+OMvXECN2WhKgXcjM+U2u
adq8+J7ijC0QqU7donRIYjZH5T/Z9hpJVaziy+tnNJHPckUND2eWrKwsgViqMNS/
GXuy6z/RUWpsCSOkLKcR51XRe8OLpVfg/kq+MEJ8q+XZ0/VEO/MbO27bdFzqbjym
pP0oWJ2NeCGytIfBsryYICzr7Qfb+dhVRrdHyJAFFyJEOpmmhJfWPEvshvqctkup
34Z7VP1BnDpTiM6pk3EPhJnGzv+ZnLk+Uwko0PZlfIOj/VYIZrysW+vyYu+ZVa17
SiHAr8KCksDMtRlywaFKLYy2N6ehfKqTokr9GVFU1YBpeJlD11rUDudQj949CHCz
u7B3RoN9YjBThQXfw/W1+owWZwgYSkpDmwK3aOy1dBY3pZCoYR/9dmS/031uxgt6
y5BMRGEk2ilOAjgnJrCWvDtjyf2bXP6ZH4cOfzu4qzHsIut4/G4vFyVWlsDhh35X
8xm3enVM8Q3+3eFwtC1KyCSA2/5TXeHH9hus58dpWCacLyofGHJ13MzlPhuBPfdm
k9ppjZoVSopXoizbm6juaUjSMCzVDiwCKpoE+DAgmkoCRakoF0S4tg4b3XX4224A
NMsZxhs6Izrv9I/hhWENjf3/CExi5giyNJ0ZxSdiWm1+q8pEoj8sdjdWF2iugEU+
6nGeYcT6s9NkYzjxZK76sWxIEWOYPziG4bycimHGyHDX8qPU92UJ4ID9HUsjxp6O
OAU71hFjlZSNQ8amUOhQqw8ymKFy0X74W+/HcAzGuIv2iRl5SMDNcvv2M1vd6QbV
9hojuNzJFC5p1rJG5S7eG7tXJf3Z6bhvf+dhOhXEQR+mkD2cHNt5uXYTu2+DCrr4
fpOelgaFFsI5QAhqnhgyMrT4AcWzl3+nyoX4fRiwolrcledoyfttzyE2QX5o+/s9
7G2R9Oi4f3Z6X0ifpoK1ycqWJ85V74wnrm1GpzwK6ayUiPaK1M2F+YlRQGRu4XGW
tidMSv1jgE/MVPeyqsyJGsUmXAXRSiz4D5+Nvx1W6r18MsrcaPvJWb2QhQXpR4/m
tY+0bZSdodrW5Ys9PLRXGULRTA+KehwZdwPiY6mC4B8KFndR6qpx6F+/0xWlQjZK
RZZecTWBwvdbs/QSCqRq6saR7Sa4HKJ6XbSWDxnJEQFzrlEGQITK8+JwL722jiBV
XAfYcNZ0tUtPTlPf1asF/8VTP938djA0+12g+lyGXNbRGU+XdQOwzauhB2kedPwQ
a9iEmV45eI6w2fNIMMGyCpTDHOencXgQ9bJXVog6KD31qNuzJk+Q+1vy/+UB5Yu4
aIK3N00gvC4NtOs6CndORa2jk2WVKcfmmamfJSeCqk13kTMHiDvMVz1pW4a37Sno
M4Lzq5xs22jtxti3yNW1famVSmOMYBwOvwSEl2mhH8pJL4u6ep63LpQs+J0YE/MO
BsIAYk6vPylGue5Rye8Y+dHOzqBITVw+sOXzfG9whzBXQIN+8UIEOMC/7i9KAGcW
xFKq5RlNILIfzkmmF0ukA0vHJbpTFfRAC64+VRY2gYXXn1ESr32Njm3eehOVw+FW
x09AGrswqABXvP0FedjF1qft1lD+hpTFGVAmhtp39V6jkmANr3UwYCdMSIHeX9Dn
i7bFxxcJ2oyeH1ese7slYGdy9D/4b2xmTm/EmsDLj4h9pQXKCnunJOEnOs1dZuYA
DE1RQwPVBel5HaLG/KgZMsVsGCAIhy+aJiVw2yLufLTNHE5T7U4O7khyu84+gJlY
qv/Fs4okA3g39iNKpG3dockAuvv+LSZE7wwzRGrVXTpI41bdxuUkjGJE0Nd8e9OY
YRk87esaUYhfPBBi8payyc5bKT/TSZp7lmhd71yaDBFwnBiROYT7L7e5CrOq6Ggm
SPP1qb2xDE+BAMJTX5HEnWr8nK6fcKftevNy6eeZVEpcMyH39BcCwAxyAVAjj38q
2EWvAq3TF3XhG1OQMf5q6LWcyTJAA62XStcPIbkRL2T1Dr1NeCw4N4gHwcKhqu4t
vRty5ccpn1zICXpYwdUrHS9QUpuzM2TAjsOCTUxXpYJq454NJ7ii+d7xqxNk/2zS
i5iy6d4sLJ6/923W4YptRKEbyXFBf9Gr3N0aaiHJm3cWxDMv+kF+cJjNJcB5rOIM
XnC5p5G+CgyvM1w+6WzG4JyX4YPR0Zf6XRe2RUkwxZ9f9W9LjS5lM2fCCHWLsvV1
jFYTjoYWACUInhUECqFxE/74RbeDSG7dFA8iZAs4EQ/pOMJvRiLDpgQ5nkRlMuZV
ZNx9HlnrpV4DudAw0ZpHLOQCHsSqsOG0eIMQzGafzVcvOKPjJ0Q+MjINQd0QqeDl
CrB6AYHqrCZee+5jSCtL8QFV+Us0UOwKAlTfI2mxVkarTepyGFxDxIn/50cjGfoY
mlsdNZdfZsa7Xw5PaKgvK4vFPz0G57csGM+tY7onfFpuOnriZx2fUWyUxlHBBYIh
y5QFqyWvMeNb/UI0WcCmpBxOGJlrFnngZlaW71xpCCAaErRxNELSmm8wLPe0Tfux
FlR17mmT7LisFt4Szt8rKBK8x9NNNi7wCWqP/2pmjNlZn6xtAo488FKT1/k5hkaV
nGg9JWModmvsdkkN438YxZfHKuzxpSI3jRQlSCNTr/pjDoAQ8ysVyfFrFRTkOn5G
YeYJsMJUUlUvsVIYHywjlnGRUlm+T2QHe19JO7D5SvyXP2A2OtD1wsrLB4DePYDx
I9K7GEsk3gwjlgVhWsSPxaDjE+x0fAm08l80rtfI12LR4i1AuhKMwHppdjsSp3IX
IROSv27jLLRWbgDQvEhkfRao8n8IFHDoeEyESMMyWFTJr1Hxl9vtaJdgW7VrQNBD
4Z3nZEtnYpRX7agTO7f2d2ov+/34r1CuhWLNRgEXOnfx86YKAhV3EIRpkeHVgxhL
CHeMF6+CaKDJN1KwLDPo6FxXPcNmAi5F+9iIZAdYGvgAs8YFck9UCqJfeDNdFQf8
kAYUsGKr18UZkJnWrz5MLeABXLA9o762rpXtZ97pfDPuyB0/1WKMp1QdrQlgvDL1
rudHB6IK7iux8WE5wL24WAKgsU3EDBtb7s6VXmgb93JaT8O0B69nHbeDAR6O2lG1
ccixm9rsUX3/w+zCfHC85pbQ9YdXtQr5OpIsdqO6HEI4mhBOkU21niQ7r3Qt3OWV
Sn32uBjuwC2iM6axERPtzzniiKjAng/lXQQ9XYOQV+7tL3kyTJk0mw631+nweX3X
q2UJ2W4PHjeGsBlTn5YRBpHDOVTaQ7FCSIsxlq4n2neg9FGQIpNk/A0T4O3MtVIo
pl6ugv5uXsYcO9snxoX5C9gz9wvP9NL9To9p2LKI2XaItSR5VNrWBSWGm5/K9191
+T7suD8EpUKbZuplhPrz96ZPwXosLxWbXq5muU2XQxPFEVaWKS5FTK0nVsQZeHC1
riNHCuYpSJ8XLHOVPzhq2nNbvv+CPDyn4lXleNrsR2RPhZhjhyAX8pf0RYYNEVni
vuARAwfqhRIGXkqAFxXmyHEhEC0PijcxQZ3Vq2wlt1wATguPoAXAexntAEIRiccA
p7wgM3rlGtFKNGkNC/OD7cvpCtbLXloa25dG0+0aWe8iAZTTfU06GbuI/2arhcLk
NCEkpTsP8jdDBem/tjCI/BjqT+k/39QTsfkgyRYh+i6Chcqwg4+mcr/b+JvzOcd2
71RR4Ns+7/PHbC1j5Uw1oPmqI+UfpnRu+qhOiq93ogm/FgcUyCygXo7JG1uMfG7v
8jozh1rjXlDUPguZfrPn/qVHX0q9U+2vxngPIkLJHDQuI42XyxlhJ01hkPfs+XI4
ch/0sEME7+V4tGHQefAudptGlmnh9cZSrIinsHwoxYuuA/AY/mO9APy4tz7Htb3f
h5MfLWBEX9vgCFDgtcLubVIdjiptDWKgolHJVBC9dh23aAThBohrM4eC4JCRTUE6
jJfDNHrBk/Luy4IVqlCcfuDhNHXIFVoGeN91M5u62HQggPOorxORqzbGtu4dmMc+
P9NEfoeKuxa60EkC8IoNICiZXdXdvcn6t/BkZ6BYeyI+Pd0mzf9wsqKJi/kvMAw/
70TbmKhnYWeuQUGkbiq6d8Rntl50FKgtJLpjl0D00jnEH5z3KncMB7Rkphb/boV8
Nwf2FxhaWKsc4kgdWuxqcSGgGmZQbs2GjsMUZqd6bCOoxHuPqYVslnzGugJkFUe/
LQsHirBJKdoB/3VjHjcx+iLVp+TCqnZkh/x+iNA21zk8+qPtzjggF1oHX2YbTSxY
P+yaBEs4siBkA4RPkTDahjjaWau7gQRXD/hq1ujmg5e11tkpYTB9ILkLy2u1I0Ut
ljxuOKdsHOxDpAJhlYpSaeV5OrnZnbBWwxXbaps5PhTnex6OGJfKnobwbAlAz8mv
uuaZJknEtqODtb0f7an4muam8UKTosSSUE3ws6lSnWqYeL1PkumtJohWIAFVRhVH
W9iCCJVZEoix7Tp+J+ucfOK8T3Qwr7ZL7cVcjCN0dkNOtU0Yv+gemDwXuBk0t6x6
s/6oHEUAF5HI3jBbFo9wfT4sLoFTjBJQlPqLBlpfOFSB9D7m5ptY0K/flvJGQ48h
4ZEftLCJZCVNULFyVmwS4QGMuqCCZwQsSy2YUP2kctWdf6bUZ26sHRr/dXQLmwQC
m0dE2B/ZVJg7DRg30Ns5PwTEEW50GSGprgulhvhJt5E/qus8INWD/1g/iaGkcxyG
psrxw+OOufSn+GsLZ3Mv7381Bgg6G6Z3Yi9SYRw/wLENSduSWwKSGvjKiSoKwSzu
wBIhjUCYdiTXqtT6GUFQhSFhgqlqYF7wg7Su6+gSczpV6SJTOUVDLMWBSnbqEYV4
Oian35sOm//C7ZH49TKJAJrkKLf8vRti0tffi0L/VNBWWPy4NowEbZyffTvpG29M
GlXOJfRKrJwU8gVstZHm2qiHur5+xsOi88UjX8Q57zilJ+S9ARlHw6HfgY4bXBSk
7K1UNolv6jefXbHpuemPYedDDLwCVDeu2NuJLo3DPbEHB0zqJVs2BFqijpP6xkBf
2xbOKusF65CEnKgd7qQ5JLtqpyzd7VbZCyV4zXA0H8cD9nZ+lEEUPUWwOggsHN4f
R6oogGrCNXqelk6HceSYUD4IbVskub0M79YxvY1vx3j8tV9c5xbY1JoQ5aUdCHjE
oIPrKSAlZYEFZ+oZ0ns+IOztHHURiyCJXcp7kXdgyrthN1B9B1coDIz12Tpz/wPn
9+lLDt00MxiuCeUrhvn1q2bjJSKP5bkohhpWVCodQ/UvliMlaeA77L1tOdm4vpUt
hVVctHYiCcbzOW1zAcMwigd6xqq9Ym2fIxL1+zbMPpak7iTiL+Yk4yxM9KXOACll
xXwfcb5DrWCQoYlOp+IgDJoLU0yPgmmoeJWuK/QTXlXhDlkNbG5FmhOPQ4GoToRI
aFAgMCsocasUl0iTR0uVQ2K7GWFYfrvy78mECOu/sj68rzWM9Bsc7nsuaVw4nn43
bWO4NboiRl9ibvXnq2EsOMdzGLhzDhBYMSuw6OkAuOwHeGjnYeIN9k4a+Dwy4FFQ
AU8ScafpsfruOY5yA0EOSL+iVk0dW6ZCQCQ500PmCaTWa7N0VvoKJbNNOUpdC9Cp
Tm/xas076cM5N6fgPya4/KaDezC7DBiZn08McAB85b+oVd4AGNruGEM6sWG5NPqu
TI0qKDnEtIVl5zKaOqYmpztHeZ9aJaQ7UIS67G27SSlR2MQQd+mCs3pyOuv9Kbgo
Mxnx9XgK0fOqp4Pm3kcStVOncBov9F8TOhPn5YqT06rEiMYCRB4mkKbczD7l6dYU
NlCb/4ThIUiaTnCvnYxI4OuRHHhhzHe/bHtnDxLh667+Eb002QFy1gZUn18Ok6cm
P61aWcKoH9NvmLcA+++9lfyiGg/ZowEgCXR5ZBL5jfZHFI76Hv85x0YiYpKXNbfv
boFiPdkAwadrhut7sJIKXj4BRfbVy9S01r+aF8LJNL9pwxL1Uf2ubvX/UiQ0NIFs
gj4kXUkHBDSkJtrQdIZhkF2b2KDiUPgI2cbiuX7FFRZmE/9NHyy5mUIuqp/KdiGc
S+MFq6L6CX3JffJbAMpMCUmPfTqGFHRYrqUinls5Tv1OWrRAFPvXmvAtEaf/kxfP
fNZYwJPXzsSAZZRgtg61ZBI9i3KJlb7bnmOkxeFhFpbgjjs/Up10721Yb9JGxaIg
4+my6Ghz3wdo5GL5YVX3cTL534sviGlUsl5VwYWgw0IxnodeD2NXXAgMCsixwJXO
5i8QLxfa8QUwuqQ7edqBKJUw8kSsBdKJxk9Jq4V7L8+UGQ9H8I+tnYfEX65vGsi0
qvgrhCHrxX3L6Pyg3v4PMC5lVREphcBU/aNQ69tY3M4JwUfQG8JpWT3dYfMuzmRM
hbSyXQ4vp/bi6SdnddEJ+GFpQxn7PcxnMtzOOhfSUxY6zFb0PoSlXwqliBl5jbo7
vKdhQwhc/kUdqZK++ePAqrTa1Nxc49a1wYGnmNJcuhHq/eoTYj0FBhN+XCr5ZS7W
+iBpfY9JzFKD6q0Xg6LnAOaF/Se5YTsdUMX8rElWicyk2hfBhrWuIl6Tv3WyPvz3
pvcpxgvVySnMonbKs2HZta6XwNYaK+dkyRl4hIvgZvV7dS36Fgg/bGRXd4krXJKe
ZTPWUiWrf1bOxnAHvGpScJ83jiLJWRvqjRvlWWdu92QxTzpZdMb/tsWRoRx9sE58
TWtEfySxjAowtZGZuDCp5CZHDjvy7nNx3WF++SUWXil0nB0Kkl8kw2q5/EBmj6oC
EQbhyKRjJLRZ3/RRMNYZIOYQRKcKO64olGF55pXM2PX8dTrHfncBSeU1w05dGiFb
7pMcgAPqnqjfNOmr72J18a1SnITI3uRZYYB238TxHlvFDBFQ9jOHMehr0UG4OWXO
BchyRaWwf2CEQ1mxsZs9O796cEB1uWFGTu/1tSiJ/TjrBaNnks8AUpiDwOmOEYQD
5AKN9wtp4brRdM3wo8bhktd8Rchx1Y0U4bwS13nOB51fZKQ5KAleOgYOszJr86oY
y1kN1I1bYlFPwEruTtmljwyn0GO2A01LdHMn13u3oh5CRCBR9SLzApxofYzHAz5i
GGSKCmmBcSiL3gDsx0hDacY+rPZ9ElKyJWC2j5YqlN9KyvKhvaQcov2n38s5nGz5
24vY0LBoZnKH8yjHj9MJ+QNpGCKUKAruqSe0Iunj9rKCo9ooGCRP6t9whGJf79Tf
c78x3oNdb9Rwr5m+tsutxzklcEn/dUKdkbhulhOfPUiplmkLuq2dxyASpJjScnj9
PJ1XgcFw3UgiekVlCB937BUFO2xizYp7eu8qzbeMDilG4Kj+beHPIAy1EHutpDRw
/FIyM3sKbPt+heA/3ynREfeQ6X2Tuv1ReIM//ak0W2vGkI6uXxNZW6A3l0Dp6iNT
bX2d12BGJWoqDiGp06LIT16Ml8KIhDX4MsyWLoXB7zNaCPUy0MRZBIbx7LrTpiLa
eBU+RlbXDyXsibPU1JU656jBbwXuPRUCYizs3rOlp9bBEqOIQ/44JE6dbgmJ6yzW
f6Fdt4UIwSNrQrVWFF+zk1CqFI1iue5/XwzPg9jyHbX/ozMzyP6C547VpjSUorrz
zTvZtsOp3/1BbmIanOWRSU/6W1KcQ3eNiGR/mTNyyAk08vja2e0LzC+gUl3+cZ47
ezX8uGwFq67kUcKAg2QgNfsL/4mE7QHvMBc6JqjRBfmKOAHnBblDrpQS9zhoU+Xd
wglXLAJecLmwcfjh2zWDDyEdqEF3uEI0tiZ2Jt3L8/D2DnvkgIlnQSMXCq+gr65K
62QdcAq0FmtjG4E9S4lwibe2Lj+LRSkbWB+Cqb8wy0j+Q9Br9+Hg4hReGYmvAs6N
sP9kM8TYokzqJ4iH37as9MDTH0lpfFcyFBDzVZFanBhHJ09Ylb5GjxIl6vpcOlLR
uZdTRN8sGhCIjwu6wQCPQoKrP9ShaJBA46+nEDVrF9AiqoYDDalhq7ID0dQZ9hgq
dcG4qlbeG+tPv7Pqhk6eKFxVeYfRQpp6bvVXisB+HqVSeQzmr5edP2yK9jxOHMgm
EU89fxl7mDt/NA6xurjHc/D+nf/YLy9AZCKQ6dTW8LEOB/oAkSdS/9UFeI+QGlWd
ppLCi3O8HrgVIPmz5sEE1qa4Vf7rXjswGh9HboigJMeQH5W2DRFEEYMRRhMsBYjc
NrdG3ddncWp6jM5BTuagTVzN7Ssv4k9sPl9tTv13Asir/ykjTo/PjZleS8aEvAU4
r0GFLdNNnlyI5Dl28aVh0lGDQU4nNrWJP6F0pnbp7CieS58ioWORXPWKaoQ8/Eu6
PMP0wE9jylwPyDMnN0oEeA5Ilcf8Po2uvrvo7/w9a9qCD6sVr0cjnCh4vnUV3nwE
Fc0gi7EfaKlMuHTVPSuyPmQtMaYwnbGz3z8C/tnoHRma6ndDb8VyhDFZZzsNo5UZ
aw/Z+iysw2d+LJQYRnx1N/3Zz4+MFeHP6sp5GufdMIyT5w/cWShdSBfaS7ccdJYM
jIYlTcXdqER64IWnRbZ18JpEuT0YUxAcY6+r81s6nPVFlU/CevpnVPWIqZGTbXk9
Kz//mvuxAfmt6fwS8x1oCSSHhj0EiR8gNZg1BziV4lTqIfAzLLnhY1lMUT3djw4U
K2fGkk68hEae2AZ1ERdYOeT2vTwZOYq4CqzpICLfSVDxxNpc+pDwa8xs0VKso6N8
zfMptes2Cl7T9A8sACz8R7Br367WPYQ902knmUW7v1YR5mdL9AN/7pDxtqErNRyp
eTi43QwUve4Aa6WG6LmnAz0rA4NYk1snI06X1p2wLYzuMXTyZSReafHJcbwc4+AZ
y1nXZfFzFL/DjXJZHX+yyngyPpMkLJfE167GudV9S4cFQeY2Jgoqje426OuqYHqE
WVDGUb/a3be7CyWJ9/v2h1yzHJ9U51v/0YIvi6zguBo5IqRDps24L4qryTkBZpTm
xFrQRqktu8IBBmMRuN9heL+5ar7Nt2KS36IjPF0zAR/UUC1OaJJOoat/8ONJzmPr
zP+Lj/5dtQTfBp/7bMTvR2EYSauDVv6uRHQ5d1ndxC6J15iQFAG3nzkC1gP7NdNh
FmBtXL+gve8k9IYB+m1CKkLZxY9Nmlc4Ll9LvYrtiuRhzjVFnwDyGyj9VxSGjbOG
8gwxM9HfICvQGWhYhRTyFxKBbK9JRRUAQIrEnJqcm+xL4ox6o4+6CP92T7jN72NR
bwrJkrQWuKWxZqOjJ3mEnSFLV003ZtIoFGdFqMF8+I9DpYZm7CQ3d6KTh6yO0m04
A6+BE9+9WR5YpCYlAxmNcWXZWN0ncnhg/KZKqno58Xn6TkwCcbDVIKK4HjqiG8Sm
L6vMiR7T7+7Q9+bR0m/jKp5DuMBFV1Z48Brre9MXk8bEPtXwztwiFZgbf0QWHT7X
6dOosT7uunNLY/AXeSeJySqcjuJUIqRxIYN9neFh/zpCiArzJV5qDyiKhGDZjX0B
re3Fd5yQMNDs4NmMCL6c9/8RENTog/KJp7TKD6DVAtWLhxssg6SsUI2LXtD5dT5h
LbRgkZx1eb63q4gfJjiZQeAY9vAArW18/Quly7Lp+VJvqxtZa3EMFFsAZftBO0xB
3SOPC7NszFrk6fiTAn4c7GMa4YqItJC/fIDHMFnikl3Zx6JfjlbAzYcA/+Mb+pTc
XNReP56l2EpuHMgVH2zuHu7GNlaMHViX6Ullri7bZ5TyFg4zgzermKC+ZfhyTn+Q
S0JcXN+LD33vfp4A5KglZWm1ONbwq+9i1qJScxNW66mLmdtUXbvzvA+awcIl/Bfq
naQsshPBPsX7bt/i+RPDi3945jijLxQ4LnqQHMwGztpwTZoy4Qs7c3qil015ZZrC
vup2Ubjwv/9s2TK7skwM1jooqu0Tjp6l6Rt0CPHJEPKEKFHFa9EbNNUF69W3T03U
rl+iZJPo3Dmp6MIILuE7JYJZEsvZeqTb6VUnwNLfOMk65FiyhHfLf3lCwlc6m4N2
kIJoV5aviF0nUOVj3f83BFJ+3Tvb78O/3SVhzeWHlUqTmD5RRVyNt9R4gQSWe7OJ
Ocg1CxZpfF+DILr5AeONliaQ/ISCRerVW/o79UIVj+3/o956nblPQY59pPZ0oNjv
hxn5lvdBVRzn1Yku5CrMCKbxpwrtAZKu9BiUTZtIIKxo635X0vmkP2kGrPJLL2mI
Ook3wfpx3CbMEe6OQk0+Z3Xm2FWq8xAd9JoeTKvRR+fixG1m+x+s7riAw7R6OnZ5
zK/6nrjysBzl4/vs73D1X1wJNLRLOy43O7yJ3hHHaLmYjvzxP2QadBrf5IFGmY1a
24WWTafCkYie20njjzjKlfRg08yDFtDgIilYStJKAed12aC26a6qdk+bDZiCauZ1
kqUCZdHDo+vI63k61P3pEyU4yGmc73KLGmV1k/EsX9rYbIuAS6jS3XANPIbXYXUL
FkcgPtS9GX9CWA2nycoSz53+mj0Ku+diWSkKCmuikzNeTJbRUj7TL9sko75YdvJc
oyIRi3YDsUB0not/k4/DmQEyJBBT7yipIeqjlBo0Uq0sru0aht8aoTO8riSOlUfT
PF3zonsuWxoOm9sE1qn8OC83whmVcv5uHlN4O8Fofal3vV5PfX9FeboRtjs8kVDG
H6uvDlQlt4ijfwu3FlQWabYPOLOgvlotwwpvKnzg55Ci8FF9h34U1lJXoXDkRpbH
lUps/7dJvJoiSDbZ1FdG+OSaE9cOza/mZF50SCEavzxlcliY4CkUfHQxINKVze3o
0tAph9C2p1TRnE9rFL2mUIedxmhh3K0vOI6cJX328PuFNWH4WFmX0msRHt3gjDkt
Ein6KLLg4mWJpRlLOZlJJWbBiimW2RQg6gx5XLVJyE+PvCFtyYPMnnALJeoUL4dG
/uhRtHlsIhvoRcMZO8IdII68bBYB6RCkI4CeSjz0ngpbnkyG5rN5VDHVbzflk8gN
LvSBPiqOqgdB2Kctgc1WF9H+oIctNuqmxjFcIWfaszPVQBnyrax3DQeyQHCKL+fH
XKl60Xk7K/NKQm99CnBG3KMhE/vR87gRNUEZE0YdKSF1TBIEHy6dVMOghpVCJZDS
bN7sUtI5FxsZSzRSZSh8SARufaK2qQB7M6GCYC7ZA7Nkz1bw9Fo3WP3WYg6tfVvt
EqulAXZsy9i/2RT/7wacUn3In2rz98RJrUqp8UIowxeVCZA9d+8CPtAu+IwE5Fqa
hURV3Pzkm/Ifq0JNBQmtdVcqEQPzl66bTK99LG47tbiXVLi+hey8y5esOP9AKRyT
PKyD58HdLXZ0H/hxJLLFZ8GrsJ9pp/7GiSqgINWIfvNEG3Lc4Jzaxad1AeQONpeQ
Aa36APj/TSAd5WhyICPHerkmdr/FcIhikTDnL6aCPxdCy327phXYtZcjKXDoxJLE
ugd8LNd3k6lKn6pAY0pblBTwkVrO5MW+65lkdSaYAwdrIhbtESE5UETj4F8v2azH
wp12ZGBZ/fpZH/iAOquTEibc0M199MSJ4gUEYx1JfZv9sgsdq8S/ZEJyh9xiTuJO
s2M9V3xuxy3oJppkaI8WkB+6hbfyIq3N+dCZzTPBsKNw9TB2h8wM8hiLxoN1erB7
smE1kjEuUbouMkDV0hqmGFMk+XXF6qQ28zBE4F3LwExl0QjeDQ7kbiBFMqd+FnYB
ibDgMNp+sJ/7byVC9Jds0HqI0I13YoQ6Zke+C0a4u/cTXkRGfd8//DzNfuES+ZOM
vMdfT1V80grzT+AtrDkByotHWDY7RqE2FRYn0btME/PEDl4XRZfggDdenZ5ytBPJ
lK99pgs59JFfvPVIzZP9tppPYS+kP6wphNKLC1PJV1EKx+Xry0jx4azy6SyW2KRV
L/qSX244scgBprHKO3HzEmCx9dqNdm/4WOuH9FUnN/VXbQ95lHhNUtx43RKANQhB
d0H44aQpDd0gYwE31XXgLuIWx5pH4B4R4CEu6e4nL+mHSklxnKehkLLD9U4rMLYH
s+IiEzruGFnd926bVwV0541MdLtTo/vxPElvhhAZ+VSAjhopEt3geiJESwe3b11i
v5ZRth5dTSU4r7+lb1b9nb2cUj+FI99JjIySwx+0+SdR1sM+jG/Nljb7dqgDyisp
Mfp/hteExVZWskOYZAJggdwxyN8CmTUJMvCNshhDompvn7q6nJo/EWLGThlC5yDd
4OywO/oHEqwn5qkVNNpLywP+x6L6Wsd8kYQ+Vv7z1qHRJGTx2wAyjnq+7oW3J/EF
TAURtmzoIvu2KFdousDng5WI1HLbeWj6XOOO+oVrzAHcged/nRGwkyOCTEAr0VFm
X+R0JfuHmw4eCLWZvF2AGHxw7Nm+9AkH5quU10TpRasw4en6R9ofF/nI4C/jOFg8
TYVQEALDhC5K/ziTxWnR6Rlu1HKs13l6QpmoYT743Y70kKyFp1s0wrmAXQwlfd1O
B3WJdZyiTiiCPlsE3igElJuEf7lneAaBx9MFwoxAV7rAnAohdR/kxOl4SCRR8tOp
qFpU0kMU92X7XITy0EzvYnDLTSbshbQ+ZXJjNN7RPRY+ay48ep1zPEiOJNtL5sMx
xhsbGQjmibpZDO4oiNv5rCHN5033FxCaKjIHIqlnBQkKBai854YkGVT4l/6nf/Sq
UjfER//eu2eJ+klS54bPgzwtKHsotyn2FHyPs4LG8/zemaQAjzM50azzc8LfOw+L
GXNBdB5UdK7WfVcid4r+cT66ymOZacVnux9ROeHO1+fH/DQleiSp4hJEWpqO8iED
FPXeLSbxl4V/ji5tlLfB2CzfE+R0RZEGRW5vCY/EYrGlshozKTy088SIL8BRLWOp
mCQN27T3GyOCgAczafZjcDvRzXmX34n9me5zvrPd1RbqNNuJU6HMPIFBgqeGsPpz
8gVlJdk0kjpm/FcJS+YQFjWhWHodhmFc2wUFduCK2E9asbBeUe6uNtuE9RvVtGMz
Vuvi+A3czvaTlcj4taIgc1aBk/oI9fqVgP0rJe5pkbUZVApjkDPJJsAErgcdqGd+
TXAf12GBg70S0CfD9kslCtIj5au3CrJeFhZhqCwSgvx5CYSNXV4AD+KW8VGa5d5O
MqAT2MJbRBkmo/wYDF3NmSy23fFSvjQ5HSpEbmyHQPmis2ugwjhP0I7rvV/CnppN
z99L3OO5AK7dYTrKwAXqpEZ2ksrIXN5GN9FRrtxrZM8Tkotlffj2DuuVQv+91jpg
EvGwYybdyzgiQMPWqu45LTn65eRKjzf7No2/LnSwP8ccbEFnOEOf61DRwfgHmfhO
AmzVZIoOJx+i/il1E3THRAz3ymW3bC0+r4p0XUaw/OoJEdb3aAixUsJj4Ohtv9iU
X30A+xHvqOzLiUF0a9XByQhCQEeVxaecJRekGV3OK78ks9/zfhypeaqI6E+0FIpJ
Im9vJ1ky2Dp/GiuETCt7xDGn3sw1MgbsJ2rAkjyyrlCcvr55vhxHAOyYtX5Vfn39
kayv+KwBsm7tDmjKgZUR0W5IsqkpVw4PptpdT5yoJPx5xcK9PWC3fbAlMhhmN24Y
KMA1oHIm8qeAr//fjtvpFzYNSUjlxt9tLny1VZgNbmJaa90phXL0e+NpDq3TGBh8
tYCbseNY0IkuzqMmUM2tJBEMp2Q/wSdI2PBJTl8RheRwBIZ0oXNwQH8IwkAj841b
BOn3tmZy8MKq/ATxrQiDgfpSa9vEXLd+1xRhdU8W7SzwabvoAYGev2ZJKEpnSOj5
vB07d/VZAjPFkvgzuC2FFbIC0svSTdsAH9BBGRfaMcHIVMsLZjQdnywYtuADq3Oi
MiG+l/HYA97jqlkbZ08zxJA7OpXfTW/cli7aLuuwpyYcD40nfYaA+oU8hZkDJg34
ql9CzdqQ9VQP1BnJdLcEpfbWbO3ezaprZLnKMsgDl2VXZbtfFEm4mgKLHclSpu2D
HYQ4toLdwgv/D7BNjXjsG3259YOVgxJAYCabugD7EccO8a2KX+3U/whUpMgTVqmq
arOnB5Y4PtpVWsFd32Abn/PJ+nyCADge6/jLy/597X4YJBkeV9Cel5G4Qm9pCkVb
nojNv3ZlhnTIkl9D/Ox3gvSqcZVTYyyLUtfNovQjA+LSMwg4AOOhPpS4dxU0sDsM
xm5toL13nPerO1U+pzK+J0IhLEvslZF3xa44RQoYGyYzzAsSl4DWRlE/Kk6FJD78
jWoklhkKYA//vFzKsfvTURdfQLnbko+fmcbhOy2NztrYYvwg9nN6p5wOnDmEvsCF
HI3JPRjxttLDitiXNkVLzoCUea8JB8deqds5wGhqfKXpLnsXiVbEeCaCgfnB9t1Q
uLi8EMqExOtyy8r+2XPXgdszE4Pwsj+A+hG+Cp3K1BVe21fcQUjM4//1OaGJo1Mm
oggQ4CWVDLFvbtGUyvdPtMVhIrfLH11ZLFpx6Me3bemNJtOF4T1rjRcRJHunPtF6
iU4k1P9MFzgh6b4vScHyv4HWK+UG5RWRXQp+2ajMQTO/vw1aUPNqeEkN8cL+LoOF
zV6yppzCUusjTvJ4oDcnLbPP9KsGU66KDoI/SQ0FnG603pgHqcpdstb4/rihu6HK
+ACoI1GQ92N/xP5Z37Vx873qNVNkUN51gE3lA9q6YFxFtVZfWH+miKq7AWvKYw4r
tUoHZeF7Ut3rtqs2xyosRsnCPT9ItZ63FNNJG1AFPB+/WLLugTMzJ/eLBa2UF+QT
SfpC7s4ATTfRSzXdbCT9BaWs4vZf2v3ek5uMVfu6kW5g5ibtTsa1PEoWbF0Fp2Wd
gegV9x/Kay0Vn5J2Rq6jfBKQUwdNhTfHYVZKnAjog6YRbF2ql+Y2WEF3FvwzeUuk
YkOIkGMSzk8w52bDe5lhrIoEh0b3Dsgfr7xZZMnOmH1YReqhEMn/2GvlkkLj1IUw
g00OCS3JJlAdKhX0o0CCV6fERs2i9kWv+l+WPte9VMef0IFf0DU5tJ2hKPN1Bxuw
vPB4jT3EvI9xOqg5LENyNYAzIibINl8X/16NIuwKPg1vN3iMsityZrOvUfECWuX4
4sw6bn+G/yxk/quyTD7OB1bZw/g25+EGSWeFOJCiAc7DjBECOPQNhdp4C1D8bcC5
AvKLYK18AZyJbeRcZEDLFAa+toUVF/eG8PR7kdY9Iajx+O5ETYpYRLvbFFxHIr7E
WTedrtxa31NXGGrO1G9uzY3N3YmZTudcNoqTMkNts7jX5840Hi8S70t/nnfQ+w2T
XhuzhKjepzmqrmy9IVnjvqcBmt054jdM72x+iu/e4qC8bhokLT3I6XYH6ga7isn5
p4/Pk53DRkXyvfAOmUoJQwSkJq14eVIpdPRV7Xx0vg5/fZtYS+Z1d67YHOeAeyiL
8b4AiifKFskvil1b2iCJ0n1WFuXFEYZq67ZYrGgVAD6UOq64x1WAeC/WAZ4mQMTk
FwtTlTFjyOyhq+25veQOC0Gc96tEXOi8vasYTr8j54WZRju48jz+PBB56XRLfOW1
41zgRw62LEfqR9TybzYSyyry8GltedaCBwbWhcWCAtSLBw+J+Oz89JZoijkyFEpv
M1AhOQchfNRepq04Y4WdSXge+vWsi3qCnUazOdSUlMRks7y4Kj0LS5oB/KlSIVUQ
w0dBp6f0aIZV0YJoQumuKu7WXELPLacqX929oXl4tAIbwUX7WWtW5h1RvpeUZc8R
1oA6y3yP8cgJw4bxc1DIxZ8kQHcp/AH4yxPllSUM9QIUoc5T1DBeibn1qam4dwt3
bkYRhfNAlMmkE1shX0yVMy4ZeVNC5f2Eci5Pb1eLM9kvGWgnDdFQzrBHQFTl79Xn
kPod7fLN/94HkDCuoolcDhWKM0jFF0XUjn/ULPf74OvVp7PSiG1BPR1X8Xua+qDF
/aSLHVFJMxRfBDZky8z1d2VKEF8BNctjP1YFeGyDWvLjzFh8I2aepsch2AM4WLTF
9hczvq2RH/A8WML4zWRpdVmwfSzH6RaYFamKZD2M2/XVFEhPbvwfG5JcbgM118e2
wE875n8j1KiVmISttpIlla8Q5EUJY6bsoTTb5LA8XtBfUAITlv2Qk4menDbM06jV
MNkjAWNLsBmnSVYTm2N7iTVawlVxxYyFFAxO+L76pV6Ch0lfItyBbyKDxTBa5/0u
nSrBrxA2IkWbYsRH8vWXWo1CjQT3evFlLBeqpGfLTRV5ja4299PCh2rekC0pEvLH
5RQvb3IKkfdahJI6I4FKFfg5Xl+8xdOlnpOrTSuieMvukL1hYmgOAd7pm2Tk/mlp
s1JKxfX/mgrrU9WEmO+/WF1x/yi9/mJswxUMJ7dAWRLuUi9xlKtl+cqq3lB3F5Tc
Y/55D1hLC1GV0iBGyVeTsmcwt/HTBhCE+TDuVQJWvvAPyv5ADkvKRkE0J20XJBCk
xIkWNVKKkbQz2/xvfkDFg97rtfr5dtRiQ29SRUwAhxnhzQd02CR3EqKuJyx3jYQK
yu7ywxM3nCZS1ywl1hXcE4pbrpgxqhdugNO5z5wytF/KvWl/WZrLhmTccnPzwBdn
AZ2HJEwguf3EHQEQZ0nIHy77VFVVWKCmjs/WpuXhuf2CEoFNPfZGRZx92Nu2QN7v
L0UA5Lnm1Vo4Za5E9KrLWoKfRF9AiovsLILktyzi9k0czEClhnTpd6L2SKNlreb2
CfOB2bgmuCtvMKyZzu38qp1rHrrLFSDrGPQ7M2k04izLvpfpIe40XIC4XzkiuRP2
tYWn6NSU2oJ62hbIKftYTSLsEMW2+VAWFk22YQlqGatFOtl7wzXBjjdrxPCHmxpu
DFm75rMyPCpKN2LMu4SoQWj6ICLBXlebj9HTIlxUW9g9E/MOyfz35vneMxBWyCB5
V6XxCddikt3DMX8KoDhgARTl2M3kcSyaIWJlV7Mm+UDLROG2D3+RiYYwd2V3kKKQ
AtXx0sHFO2l2DAEQv8RXLCQgocopzZvZHQ39VDVNaNFXLPvDFCdOPCQ4vzTCfkHU
iLRfjedAMa0RQEZFwBRDYKi/Gn9C1DfL2RGBIeD9OmifWeHTN++5xFVkI6tzRwEr
UiEXdWjwKJhCCpHSVG+paoEG9Zsp38OqSt8G8NjH8ZPxPYTFADLHUr1ZJb2H2HTp
KM3XkmogubGbx7YMOLK+aFOC1bSWI+diwPlYhY9CNNxIsMvynO0Z8Y9iTAcxBrJK
bbF4oDvR8EkgPdN+s0feXov3M+HiJBgAR5pnzDyY5khtaKaEdx4QonkCu8Gn3K5P
YyALIuAkX4hiSMz9BTAhgi1EDyL3grUHwm5ux0ee2pp7ANwTuCWxW9ra5Oc2gV6y
UKgHAmU4xHsKnuOxxTpGZ6EwhTR5gT4C5Ed0jyTXO9PjdV65BgoHrzzc8/2xTlpg
8zDh8Jm3zDH4Ll5zzaPWd18j33Iv7mIKkcuzAdbJ44awAaUxE1540ni+KdUMTUds
fuXZtpxMF9lM48fPRr+K1P0b6HcPr6xV+SgxMPpii7YrW1FTJrT8Ge7/oaSmKcLV
lefEPQkPvjLgcUadeP8I8kqK5sqDcTKZGIXm0IaoM5vD+3kNeaOCh4ghaCoX1VB4
ShkOWKANPfW3i8eXX4udJZmrPPtWvcIP1Els++pyGl9LuUeIjMnd/roq50YssOEE
gI2mwu0f37EZwxo/I9QHJkHevS5XHZ95uiAv052mxGUxs61W0kQpDls6D8d7AcTo
4+KcAJrzFAW63yBAgKnyj/Plj9vij8m7PtCmKLWDI9KXA7nEzRKNQl3FLlq82+Ry
ub/RkXtmwwB6NjHsTUDmJHqTwS/i0v76th7yDKSH/O5Fy6phXO2S+nw6SZ33NGxM
5+m1lDMFynrzwWDf3SGyTTu32ETnyxe+kslJcfNnnpcMj1g/EqyFFZywAi3n2PHV
k4UCdCkghRQtFS/iYdglJOcwWDhTDozH7u4THBErbgKL/0SwHKOhORdOopvl3wjz
JBRNAR/mxhZatw8IlZj4BIZlzdsqsOZrNQEllgcc7AVWdCQCfNatQNHHuTzf1Qvi
F6MmZuf7lJbZiSoTPdIRdQMATZ/CIrQUx8SpXC1w2AP+o2KjDR5YnPY/yPXaEB+W
7TF0YBBh/B2aRq12AYAAdsfKieM83yWB/MIEad7r8CAJEJxJO9K+Vv5JPX9qe8/n
bhOfofOCTDgGExnjVLcuagSELtb/VcmQqH1UxiFMm34POWb4uGud/L9bMQV9Hj8n
RkhAUQHhf6lH0sJB/Twc5P8McA+DTdRiGa8A0UGNh7cXw1zHKs167LAgPHNp9VR5
lNrChwXhScJs4HB0stS4vATKtA8EyFGig6sxzfYxfWi3kVH03q/kMJ+Eot66FRj5
gOEHRK6B290hHWp2a42YHmth+o6nF5y/FHqZOeZUufcx86gpYj12JbXsFej3DNui
5J5+JeMBpdMuUctWTDeWFwEi8A+PWDahVoOpdobqNthKoRIRiKCJDinDVyZyjRBt
RtLqVIUhiewBfmITjHQJt6K7/1HZ+fHhuXpV8W9H0SkOx7rjCB3QJ7K3muJELCvE
q5FXn7or77ZqOfr1Wpdc7jnsodtd4zTyayc5wE3J1lBIKEe8vzGGVvrqSeutbfqh
K/+cwQI+0G640lMwVYVu8UcxURD7hAiDuHUKL9nsjZy0tv63iUPpd5wSbdm00/tK
F8ut9kKt28abRsa4FHfG4z5fSIS79O1ACsmpuvgUWSBddAEByJ2nA9hA3vWjL+Yv
Rr0aTStsUFVcI40X/iIJAYkAm7JgG5btoqM7YAK/KWn1/M6OwgxL4bjztPNlfpnp
45swrMypOebFMEp23GJ4oR5CITVG7WvoBTl+xSE/3O4gihQlS4EX7ff6Ytn5ZKAf
Dg0XqKjcFG/tTTjSk8qUvcIP6jxRkZoGodUcJRX2zepHepdYIotAUoGL7sIRP6eH
n2v9hIzB6Va+Jk+gRALt/Ou50ztQq3pI+tzVyLkbh0RMe5S1G/dUMJ8DFjzj6eSl
dLMmFIO9ugBFjwOI/6LyBFFbAGZEJyOlckjF/oAp9UCdI2jTCLpiew0OowbVq6VI
2rEt7eOnmI+oQ73t8NB6weMObxQzgwsUSPZi0GoYrORrvUUsjS/1qHXLSnJi9NKD
ECKPnAl/0LWOuV12+rY/Z+0/YwI+EfCbu+kBzsN1V4LTp7wwd7t3qWK48M2crTgq
7eejcVLJU/vaYiCM+yLnUFHFrFAeq28YX40W1pCPUxcYVvJ31A5RKI63e1YfLBLe
M8FCUcXKtC9RJirOa7L7sXX+00nOWfrZoPyEAlLAnEDgvx8IPv0rKT7L5yQ3Grn6
oeqVbItJFC+S1L5EHbzYu3uEHXm1tc5muYip8t0RpcbzuCuUuhmR+lFTzriNtShd
Mfy1vP71wfet52AQvZHJqUIthCzUx8t7LwxOilU4KzNiKKZEINq+S2RjEEZX4VMj
voWxA3glj0CI6WOgKHtMVDcwBxooM2jW6XeCaAROABuFeo3b7wF7jRa4AXxd/UK+
XqtaYDEDpT6DfUd97ZTheXDJggMOVbmAhXA+sjV9MqhENC/gYNQcaInTfJM4S7Zp
mToygfwMkflj+nVg1y57QrfD/QAP7MIrLLy4eDf1eMRJFw59uATb2BXBw806Shju
dGBkBFAsNzmQ/s81KAauzXtmTP4IuvDfzTNTyaYhnxv/h+5S8j1pVQkdshS5/oAH
9V0P8X3ZcrKCGVUHVmrmrMwcV3n/6fkFJAEtFCReb1URhsvSVLcjSOJYcApgdt3s
OjfEiITRZZpAqMNzjpChL3iqZgRcvH9pY7168phUVMd/NuG5jv9OQDAe9o34Rfnq
ai2q+Wkxq0KstgYcuYyIIxrc5oi4rHCQWRawqChw1MLipQusemvBUVAPdX3kA0sk
WmeVxDYL4sa83BGqYnWOdhTmmo7GtpQcVmVge6J304O4xuW+vNsFqhVCtIM7ToAP
VMqSD9iYgwqWiLh53ldMFVzwAjcS8KyrU0uUPh96jp3fBR0d670jG0t+LEnxlFay
LqxQkzzinwScBFzP3dzY3K2af0/ivF2En6w1r/LUI3p4/+I/a07XTjfm5pXYnSbF
rERmg5dVuplwzCbkYiGguTuHuwBrQEeoT95Q9P3hsOKsqOorWs4mjrq7i6QrwUoS
x5e9A2e/eBS61ayg8sMTyf7gHexLy7t1BqikIFDtn0HFiwwL/u1ZT5LvWn2ZTX0n
pQIP51ETapY+owoA1vGMVzlLWBp9Ahbi3J1YOoWDaDX863IKT7JZtqnEzq6fcnp4
++8V4hvpyIUeweFhRgZOF+Vr/7iG7uO9FcLUW4jiqwp8OxSj24IvQe/2mztSaZE/
mVvgjrP1a1VgMjajywSlOpOmsEpeiqt4LDSEsXRfOQCW4jz4RIzwhwPUkVUJwlGI
t5eT1KCl4jRJsB5JmVM0H1gY3FRsa+hOBW25N9R4usEOlkPq15CbVz2RRod+GTuc
cUHw53+LX+LpglePDSK5Z4brfC2+5Bp+BjU5v4hILg0JulZxsgwqFuJDKoslT/9f
mTgS0LcmeTEPogbZ2vD5X+lpHDurBUYKksNx/bbF/R5wN2R9J5LkNJsbqMJtPLQz
X0dLzqIEMOm56aVcS7dtuOD8XewuvSLYVeXJZvF0bGpn2i10jGb0DwKbPSFeCX0n
ZIlADdaZLBOC4nx0hjPwdbq0wn2LCeNyOEw155C4DulVCtelsSBr7x+4Z8bs1MTm
Pae8V0YI8H615Y/B+ibluq+wV/YL8QU815DbgKktEYpecwHAY93H0pdWhhLkeJrg
UOKp2JqZGOZXtmY8dwgUch4mHqbLtC/7NZzyzmR2I61P9cCKm5Y1mtu3JCtmb3+p
Y5XCSswC82KdA4Thgmrgk6MRpG1ewBowCHQbCaEOfes38dY2fEMFsRXNSvodhlTT
vzXBGwwt+zKJZCtVprVYV+F7oVibQ3LwFnQXlceVlpnYKk/EGi1ffK/RvqOTRWzt
KmutIwlzbxadCbwwlNG78a4w8LJ2HiW01dR+oA4isBL747u/DvIkOhVE+6GRNsX2
YwBB+OFScelzsz8qqMEvVXCrtm2v7kBYyLA1F25ZzRLa5pd1WUwNYn0fRoQ/l/JC
WpL7XkoXjtD4e1BMzPgwi0u1O33Zl2buPIUNVURIBNYR18Bt56b3SyxxAmWdAEGw
CCpJHm/5bkwTYct+ORZzRy1ty9079c+7Al+BPoVwctfA4Pcaj17wb/EGWnItnaQm
CurXzs2f6AJc7TrdK9Cz3/LjSvD/ul6GSR/7afTVAGoZXwYSE5ZDX6o5obhZlT1h
K1CboLWH1dD598PYnwk2kU6rvTdaiG7C/TZYmXZ6b7GVSnbwkyvFABDj3cp1pA28
s+pD0AMBacLsysRDX6HodC458JeSEKsVXM/VdE0iWK3XJYLa6sRemCvD5gcGht19
RlPkZifRAmLXLPpLmbASDlKcQD5rA2uKHIxYUoxZhmDpO0gL/N+v3ME7LV/rzn3s
zxFHX6aaiffi5LEA5QiUkaB+odMjCwhqGVnLyZ5dsQFCT+1xjavMEiW2+8E+zUzm
IP3v68NkmgE2iJ7Nab26NvxWVSEt9SJftWdg7na0zgXkNEziXOSwgcZLqlzL6lXf
uvOB9zQDAwwoxclIVT2SDWc787yU7wHoV2j7zWZgcui8/YbH4RBsOAwAk4Yg/Y+h
SKNFQbhUyvOeteGqh90eeCFO6trRkLj9n4u8t3uf8asYYIjbs2eQtNFh9j5U5VZe
0P9MyXSk6n2YQjbeYlcmzTW8fQKNmAqBJ5Iym8PEtHJl+KHP5aPWWo3yRhGbC5zX
60OHyldS0ktSYGvEbC8ilqLbdpI+L3LJmc/qOxNVjaemujJCowskb4t8cZAWPNOP
164Gknporz+9mzbY0cuplGn2ak/OluuPR+Dt3f1vEUUqVsHEwC2oRGrtyfMx693H
tM440c+dazV59As5qOWujGrYsYU0Bgpzc77+sKydoxq45l0/5Ot+cEWz4kvX8FI1
D4kezCSp1qXZ7RKP3//sAkZnGV7i5lwMR8rL8SzdpWrCzVARbu3VjGJNc0JgFwkX
A1gY8qYpP+lIZHn+1mjBpf0Yyn8fA9mxXQeNyVFHFHSM98tzHXUZAhE7T8y6+MjL
TAHsX9VYZzWfRpqtGWPUsrtMKOyvH3f+VyR39srHKpTCoDzb/zhq4SjgBQvxBrAR
tSxW9aMAja8VeRm0CLFb8YQSVlZkba7V9QvOL8jYdisBNSjIH8V51KxRM6vO9Qw1
9CqWZuKyIeQqD7eSFxMEwmRYpGs6/0wtlEvz9RQO4B1x9EkQ5gyNKqw6AAgxdTzf
YzwTxAqxMUqgpKYSNz+g8KJeEM1swz726nKXfXa/QFJDkSOZ3RWt45i7fbyf8TMT
d+zruRUf274LngAA2Oz14EQChQ0FNXg3dRpapNWfnVhMWHI0qKsdWgTFyL6Qzrvb
fQxvP9SWiFHJbxwCjUJZ6sxhVcd/iwg+++esx+zFaXiVCLKmRuLJTi+UM2M6xJLr
jLdJbwujz3ks4ROd5d1suu2IUpfApDIxNC1ldKI4bgBa1pJgV/sx8yPrNkuDIAZd
3fFyCAbfay3FMy2SSgNfJd3pGt7J3KRmFpAjBPUXtRmsrd2iV97hlwSFYCQP8h1N
EXdZFc6tbj6lrwEreTh8QWNqv7YeKSPcnqKP8S+gzLHxN+U1gwZUXSr+L1o6i1ss
dFcNxbrxNBBcKhZSGimUdX6i/9L0/L3R04Xz+tF+6t1Z8CSMr2ZFoNxGa5fPW7TG
l+d6ZwSuX21eR/14+sfqWhFFzWT3PwSxQtKHCi6s8NVMCAAV65TlUoGvnjotlxpH
LUDb90Lw4aiQMziJ2jkBx/wVQeyAhA0LCFX5kLgfkku/Z7h9Pd/Ymt5xmeqMJu1P
N2tW7qFpySZ3s/HaiZ2xbFHvQvAenD7kN6Psl0GB0BWyRBHIzw3996i/ymDqwsBN
GyyLkiHbAtK+tYW/JCC/OcRzL44PFf30WJSUCkMaYb37f0u4zYZTXMkruNI4qiCn
LMxwkGtTKohoEou4qcuHBRVfVjTGYt2JfZDMFzo5Yi/5bDqyTT5ENq/zBETxM5zL
opMbfqyKT+muoh5ozg364Tb1vLTLImwHcQWosBUr8HqfUFwwIscSzF7Mx00v0bxu
2e9tRxduoJDG1y3RYrB461z7350imRKp6mgUIN01BO8gB/5buvVipDcdM2xdMsUQ
Emz3bz5ceUjuEqwY1NhQXWPfHAk47vgTvnLXhhTOuOIjLYUNebEz90A1/04EFmLM
uXQ9qxEg+bAct1QFtLTDWBnAiLJReHcRGNL9Iw6sByo0wq7yuEx6jW7kniJHEAFB
Gk1lQvpz8bu7iz/ocioFomR5ADczeHd195edbewMG6nw2raMOx/XjQxSQB8WCeOP
ql17cKz0pJVtLHfvsgcW+FxM9lPEX7TG7MFdqvFKKllZ1uRtzslS1N/yTCgRFla1
0+UnanFkTXYKYRWXv7eZUwOyOVc9ew08echfkywmXUTY4+Ur2Kze3pyv2FkMRXLh
xWeoA5PyMAN2wZan9YA4MHhX1w8NBYRJvZht5q1sJKFCj8adSbvKzM3Go8FAnHDH
5nvayUdmZR+HC/EHif/vfmXeKC6UEJFR88HtAFVrGy3OtQ4r4omLHyehGdrsS+p1
goq6B0XlJcXqXD1F6zds0WtxmIL0Ui2dp0ZeOt6eeoKUwcLxetBs+Cex1HVhTHI0
LyDNOKbog0Dmj+ji5KGcO6yDI6JRYVQ4umcs4KXuvUB6fM/pYHGHD+y2nTLOANmO
7tJgld2cIhyyUY63nR+//WorQHjni+IXQWdBhBCpRCNn/nld4ymjfXxR8SXmkFE2
1ivY1G5qAV9eOB494KIdeDgjHu/fCPw7FQ+7IKxUtK6dJ1xMx7c7xetgEyiVk1ns
/IGnuUKL6Szyx0hLSibRa01cykvYxJe3YFnOKDKrzArWaE3D+U9cCoivqLevXIVO
LxWntvJghxgTYdguCW+rtBTNZIstxTtIx1pgSRM21MBbhI3Ee+DX4XbQDVmZ8Wn7
nMSwYbbJMY9X+hju7jZ1xMFrOT1oKAi6nCr4jxX2Gk7FoPq54/Dy4RBhD73NRYkg
VXb+nmJL4rv+iLTGcx+EBGu9DAQQTORgqmpScFUq4R7d2b5Dr90SnUiAImmNYD+9
za8bp48WncWD36UJcxb2mLZaSrSnEjOaYzE8RKtbs/c9PaNQsTeJJR/o4lopprRs
R0C6lS8iN04sBFlMS4ibDD/yR+RMGtwQ8lBdCu96gvQLqIzBgrJY3C/pXqqW0LjF
4wtB6ZGk9onMxIax7nYnnvKWEY67shgOixeHF5ixqWJ4gMH1nBSHSPr7DseSiAy0
Ie39Gqs0VSz3Pu+Yp9h0YNdwW8tGu0GVRMh1IgHp36UmoCv1u7YFfAdIGpJdYfC/
PW4+uGkzACDtT/6q1MlEHs8r2AcieVozPTottIDnaIPz3cyv1d4V5xQyY8pFU+Fl
y5Uos1BHJAZnLicb6m4oi+q0sLEivvTf+y2PsfV71/9bPLcAnt8ls/P727yrD16n
fJbEjx/ijs0D21tO/jqXmi7Qf9XY4udj30BFLTuLpNXvjDC2wttwtS2WJ+XA33Nx
zAAARPShOzACZ6BFfJmcb0RazF++VM2HM5w02DFOKXY1keH3jj9S3SZ6qFoJdMeR
Jd2a5CpW7Kw7+2MIAlfAAAX40e73KsDyWZ1swQsNESRsJfRCRB0U16c8dVgktiAO
4MrqWSb4yRNhlXcs8rV9NjYj3bOE42GKEY2qzH1hcst2PkVFeJT0HGKoY4o64sWr
dC/y5V96zpyqTmA8rhxH5Mj1U8aqzbQ0gGA7mO7zRnxXKkH4CJCSjwj6HI59DAKI
WfdxbxZaJ69qTZIy56pxerA9/e5xc8XnLIquQpDeFWXIExZ7DNUdvP+UIJb/2t8L
AvAZZLKJVj4HdTwIDOkjI6cUbodMJt4OKkeG5MKy8aRFiE0bq90OJkGvNbPv4oo9
Z2AFzdX6UjhuCPtrloApF6URfspqy3UJG+27POcnxXe1B8AeWR3Cg19A3bPwzTrq
aS6scrADaaCbp43VqS5z4ly6dpIxhWb2ubw4p4Mu/tlCnNDNBjIR5xA60RLGM58C
fCQ3H+d+dEdL4v0+eajKz1vGsIV2pZBmwd73UWq/Un+TURhTpzrY4OnNX0t557aG
TVVp6bOy91zcWvRpyy3hTMOTOX+Vos2Dzl8/pKOlnaPOXXbnGmS+gJ7vXszfX9J8
uyq3Gaxe0OmFSnHvfyMK9OJPUmoNVTsa34QSwoZPZ6kF+DpjTk0QE2shFTH/UPrU
XdBRj1QgspmFKg3jqMuH+is5bWvKGs0QohsZDaxq+DyB+P/p6QeVGpSqsOlWgya2
Nh7Z5eQZyE8NBlmIW2jB9nKPBwMIhX4kwwXdXmSewoTwN6XB5d0PbBu65Yog5Xwv
gho+62vXqPORLtFxDC/i56U0CQASkmDbl5csNY+3wTjY83YQukUeYVIcafJIcWTb
k8ndrGxMRi0AT2w1FNXrLQ4lwIrhS5HORXmA1FX6KAqdqy/X6UdsSxYp7nGZfOh1
W++TyxPpZSIg2GnQXfJtDQ4A23wiLXsewOUEyaoVNSOnMkvfUDMMz/3hrrUV7SgE
XCx1hL0f/7F+KdJTUOIBMkTAO98MngZcFBBcKhpBjMou+nAl5OXc6jm9PjDZDtww
rZqSXh8Lj0S5xWjmkTnU1Il/MyRqI48RlXep3Nd/gibQjtSyMij8u/kvTJ+zot+J
pxDoo+0cVMlJqgp0CupIdETvfHY3Q3jm2nxUcNRwW27y6mhtteM01BVuWEq6DHGT
Uw3QEnseJjV+yfbMotjDJ+0X/s37nZe1sXdeY6GU+0Lho3dIHQZFetgj0b6kWrl8
fvXiHYGa6/Hyy4rRcZtt34gWZaPD5aWEegKNUdSSrOqCYQQBJxIWHruUwZvd5qUF
2yl30CwHBXZn5iW1rUY3BpXHrO0Kz+mklkCDR3t09NhuFm8J+be5ijVbxWOVTUiB
wNsWgZc9vKQz68gnAP6c71/CEAjPd8IMt6bfJDVYKYpCl3Zm4k5zcGwF0T7/C40q
omuwzBxzLluCpaT+15GD0SwoPf6+jcTt4QXUHO0jxszPJ368b49sgcM7grJ1oGcm
4BBdui5I9GE7Ik5uuPkniN+kE+ZztQ9TDuJ+HLirZ7O7Sy7b9DSv+Wpuq7J+7xE0
RdBMUUdTbdFCkYhIa0Jb9gjcSlBdlW8fM7DZl4i9OgMOIUYJ4jeuLNBSwsriK+yh
OE4poCG8HS0rsyv+kXWXlugvmQIpQFS9RkUL3O9Hu8xYC17T2/alDJj6sTMJZjtJ
DTFnnyQE/zCFjUeHGEWIlGdMycKw0XuXje18Jp5l1+louJNWd2ICOv9SMDIkeOgm
6yk8s8yXmyzileUYMIkxhzT54/wYIzAxLZ/IySm0T9v/TWJwr0TGjqhtAQSLD7+S
skT9OrWZtihqxUjRQ1XvuxVQ45GRBKD8abZacT72aNSbknYpcfk0jOKO+nxN0Ryi
jNNFVW3n3gYjqZZ4ZJgOupEuasqXNRjBjSLM8PCs1E45s0CF8MlNVAdhZnxST91j
9fUkb6kTOj8YFrM6YRNRRib1S/+jgUiT6KkohVEyAiZkMGIZMHALgbFYB/+VCnNZ
JCLZGhvgGyazvyvLoLmuYTp8EXrgQtgBVkXuybuKuF2RRot/EvT5oS0ZZXfS5JTi
izhF5NOc1CVeEo8eLK4P/1sRfaC161YHCb/ErKlTROfNwaxl+it5HyN8zJdHUC7s
M4ajT/Pbi1sbomqLiKetmmtQg4eLfYdCnTcISC3EsFy0ehbg1/kCD/3FsU2hxqta
LnAcV34hnUgt8XMvcnmv01TkjHJjcGALUpXagrl8NPZ/9y0lmcPzUFmdIN2E0HJv
iPZV8obdFNwzg8pkwNWaYQWu0yok0F2YCnW7iGODXavIAIV2dWyJ6ufjPaF4zjJY
EWqSd++9+DLpuEXjkmrLhaEEVxn47EylRRKhkMfZPgI3uLCREAK+j5cYWv8PevkG
V9b2q0uGwLksJcPbjrDgMedGTakQygLCBXWCmakjeyvHEWba2qD6hQbCwiRlYsex
+yL2Gx8qrV237Z8GPKAFU3vNGnO1fAO8IxBH8b07fxJGncq3PqtSyAGnGSCgJTDW
sfDYIHrBmoDLeTO0dUKm0uS2+sqqo5IuaBLBysQeCNoNOzTK8r9Kp6uWaFXUdhio
fPbYCfYHMqtu3fgLuuINRzz0e4JeaM2zBLxwaROr387uwNYugTZ0RRrC6BiQWBt4
W12cw5PsKF0aBf0Vueml4ECNFhvDTOoI4yFdGkmAhl7iyVX95w0O7LULoKsqCfkH
9Y1l/Qd7/t5YKkfFcxW9mbF/2ESwQuDSfTTbkuSH0QO4ZUUHcvCzh61Q0Z1yZ6a0
D8Izr04Y9uWqW4wtzTOn8kZ3whCQOtsKj0LSXBmd//KU6e1rtUffIC0y7IP6eCBD
sR3fcaZDbw8C/m5w6Ec/YLOu/uQEavoBCJ4uY3jO3NKVNwr3CmgyOs4jhaMsTY6z
DS6iab04AC3ENb+y5tT0qRwsZywSkHA2uBeLllauyvzIDAVE72OF9mTxaZkuy5x7
tuoVskCfMRbBrL+2kQyMP0+ZX39F4C3qVwgCYpBYVtRIhIx7pUV7RFxu+rXUJYmE
g3FtSZhqJgsL5xMmHrxV1F4T3RJlqCnDmHDaGwK/RVjZTNu0lzaJ/5i4I8UVebIv
ZEdlQ2AvrwgKUpUDhab3dKMP9kQsZTKQb/3blhfqodAm0cHPfLoTfIhORHI+Kx/Y
O/HnVjv0u2NzBVd7ecwboWgiid820UlYvdBZTGnILd4bhisMBoj5TmSNOEmW9Ial
qoLMtGJgza5MK5hufqe37T+kWI+j3iyJuZ65gSlzrXHlGV6+5vgKOn0W0mwM5I0L
/Khd0txKU1XtK6Ifiq3YD4QWOwxkHZBFcpllciHlngcutVG9u1VotysCsGcNn8py
7+hJME7gsBGwVVLjkvLlb0Zv4TsOY5iPOHGLn/Y4IwmvAsZ9R+nPxHt9aJpjGq+D
77puf+Zqxsrg1emtH1xTpUoZSgLHk7m9uBAspUzXKjgPZlq2/fCZw6fs6FDAfZNf
TURiOn1+qDwT5JK3PL9mknCDvqcel0nn6PCcJuvANI+6CPYyQWU3EiRnxCGU1MaH
ny2inX7CX8fSyKs0aNyRMP8MVRkjlkkDO89UphWJNtNC4HjLm39AQHdgoioW36nt
cVpgph94zIYzaLZL2L/PttE/roUB2+XjH4tKRTpzyQwYZNd/820lzvd8lDzNjg/X
+eoS9idw5Ums96FyWl7XZ/gSzQK5nLnj717kVjUNCpEUjn4s4Lifo0i6L5NnVML+
v21ZOzAq7ZLgjirwCm269J7wq1qf2ILUAvBLXsr8aUEc4/w89c62HXCm0KNhe9V2
vDd4QLhEIFAzgyoE2P2BBE+GWZJeDPUgIdowMaT4qMvZkgjo9PlYYVGkmTUzkWQY
5X5mzvjAfh3NQ7vE3f8R5R32u1thKPTXZJSwhYOAVmmpU41ksagh4I9vycll+O8d
4WJhfHro6vrnzTDLvQywstgJ8ohrxINePl4Lrwe2SXTBzgLi5p2xYs2ni/E44/Gm
OL8jmqUsFDw2bCoLp2iqCnl7Mlw46lSQ6KABBbDltO6wKj0R7Wnofd1gV+am/f22
OcFVrbrDDtd0ru61xdpYFBLK3Yv506JI90PoGI5jwmh94tVibdJirvRPC41U9pnp
erOkMYCTeMGEJLXm7Pf97wfxkZU4ZDeZsLKAbGMos5N41GaGeyfhmq5G2U0g/RKo
gldbH3eSFoTi8a+OF8QuSzIwW+9nAJqqHmvTwLHGdIx/Cin67b3XUy0Qvu0FAGk8
KMOD1T4bAUlN9zMVx+bNXDeQJd3vSPGfVPFTIBkqOcjQxz7rvjjAf2/pWbmEQZSb
TiYNeZoWEuphtbuu3m+rui2MFmqkTfKrtOnmro8Tr2MwuYlB617ci5QXJ+WZMYj5
SfO6/HShhmuUoAy3ad8ZOSSRXusnULZ2jTVSMGVWuXwUK4durYKUogq4ZDtTgEuc
4s93M9Jz9SC1dbYLUh0bw7KwscsNpSX0K0kCPV+9xX9QNUcDEHq41Yq15/XN2Zdt
QoZ+fBCPhu7giS+km0r0GtJyZlxbJY66sOwTJEZA4cAXcrpAxIzZEL5A5Hp9QAdv
m9/5MiIcLicEammKUQSbJW585SfR+OFyqt6/jvQrQhiPqbL6XDxMkypIsQbMjYJ2
mUka34dGuVX6DtiPd/ZL1Bxddw6zQA3xgLlUYnvXqVZhBpC75TxYSR9munl2yfPN
80WCAhzQl7+2dh5Dnse3/nHAzNzuRugB0Z3vcFFAm762JzoMJ9zZy3CUxszGDbmy
3TclIXu2T5R/HTbOFevQv9yjIcO8AdhpH0K4keAlxR0CxcD96+6a4VcJc0f+hKKj
q1xZ8rKIH4bM56VzKoUe9QPsWnSs9LasURDsBJugNLTqcCHasXLRVTklgqcjTSh0
Wi1SlVVsProgRzczZ6GnkgWrpcnATZuWa1zClYZb687t73leYPz6wO+NzUnolc7N
LK2swkcu16ULgYrq3detcEGaLUANSV6yrE/Mus3eGhxFHtyVfQF5ns2bwSJIBlGQ
US0SF+RXpoDg30sptwHuAQSCmZmJun6tYsx3BFx1CWcz8LPWRHC3TWQI1PQWD/GE
gDuNNuzKYvBkXeBDQH5T2kuGwBiLJ9EsXZKrXXUNLdVK2uW9vKIrEQ8Oj4sSMVeB
MFECq/upitnhE+LCKQ7wz0+FgwjECr5q2Z2/xnyAKow/KH89A0CeFiUXyKjOwNMU
eUkfgx4ffVlamTkGu4Ys5yuQ8fKN9gfQSLQ0djqmpkTdPIR1swBKYJER3kkxSCd4
BrlgHyITw5w8Jtdp14aacy5mcuIURaT34sGwY0DlEsA5d9vkYgHrCN1JfQBw+aP2
AOH5ZUlhN6L9kcg1bwCDUfWQfu2RhoN1ZW8tdPbyFzCSaxa/SJj59/e3NNGlYmmZ
YORtcPtf/9bKlSaS4+JR3x4lHunKEe0vqcNdZwd4YLwylUPHzq4QtNy8MAir53vS
apdTIiM2dMMd44nGg0i1+XSVqw/WwdXpjsip67ne9fSSjgBNQTkjGfK+vXJRms/F
CwoPTbiJY7PfV7i/7RtZWzDIvMsPspQTgajFAUMc5qKCbhBEWAR0U/1EnrtMaTiI
h/NAK4ASfsxvCPZnF1ZvPNZEGqFU6qH4tEulmqk554mEbGkdual0ELvKFSWt0FAT
6twZEuyG/4tVIUblUkTGNoqQXs90VGv9u7oelXLMFyAsSAPe+rTTBV7dEgGe7Uo4
Z3GNLXy6CbeGRAEmUqtir3IR+591/+aC7eVoK/e2Q3MZPwRdlTSjUdzA6DM/yzBX
tsQUkLEz7bKLXJjDnvwyx4ms+0O36uVowAzvl7EIB4ylOjNowwy4XJSfKOCCjPcw
/sVjjTO/8vnrYhXc6/7JLXsMNTfF5yDGc2DyD3HKwCbsOIXzAwtlV3+jpYeCLfdz
lDusim/mTScT6iZX2Uoapn0pvp3U9eVmZVkWooOJHkekLZrwycFujffevnKiFY+r
APfEWcvZzuUhYAOaP3vyEJw0Wm1Nj/4ZixI0Y0hrdyqbPkYH6nonZ30NdPBmii5j
Jz5QEMtcJtOQofZpTSMDHyvY1nqrqgfoTsteu0MnhQ4H5s5JZKW3vpSz/uxFX2O+
0BHJXUBjpN+9e1UosBcuMExXK65t05eHDl25c97HVQ8VfiY01aIH+0Z5w0PHFFur
btSwz6twPwYLSZWZj0WvnZXYYSZBrPVIFpYhlEsj18Tpl66dw6HoT6RiikvoJBkn
+eIhSbH5TLujLEBz9E3bWj/b6dMcr4k+GZhdjDiiHEwkXxmMAMNLuZCD+7QgbT4O
4oCrSpK6ICNaZvYONW6Bdbts4G0WXyZKTpBn+yxfZMSDAFauBNyKRdDs0kUm6S7z
Tt91lZJTEvfsulItFVDNCPon2kSmsaJAJSnTAmuzRJmKag5qf9K0kUL45f8QIfzI
h4yOMeLnEFkMMGYUlM6mVn0r7fJ7sEank1b+YOcblQqbjLbIIxFDCdjUTay0LaLq
+TqMeGYRNqgwQxP+m2a9Rnmx8yLpJqJUPQaX1zmnzNeKaaJG0aUpFiCWT2Yk8469
RzF4lPToeA+mDZjjx2sL0Xk2nw3WFeVyah8GnDFm4Q6Csf9Uig1uiE+YAjTIJEOB
9Z5V8flUXyn+MZg5ubqx/EX6aY28ndDayouoiGLxJgWy6Axt06p7+5aVxO1a/0sk
Z+mA+iaJioALjfH694DgIEvEz7c7gvBq5P8hojQbQThXObv+FgRoMSI4PaemBGvE
vi7X9XkGbnKcJmvm2LpJ5qzlrcjRe9TsxydogdpS60UFOBBRhye5q6r3a1TMf+ID
HC0B2e51Gdd+ov5OE6U9BbXAr1hp9VLhFRp3z0GN1IBxXwiDLBmQNE1sI5tJgi1U
2nOaWWd2YH9RwOb3pP9kh0dnANGuQUSOO7vTI1uTbRSsbsrY14qAXl7n69+y0w+N
KmUmhJ4rncouICKgeZZD67ROVgntaPm56cyqxIWJS+Bihgu+lDWSbyiL7Kitq6ZJ
MG530HY+KK92bGuhx3h8qzUSUPW/SpOvih7DqktrHGMhyWktIGGlOTajRhAnhowk
CBQJlefuXM77xWliGJbCil1eA/dkFSz3UXmA4YtEximLiye31hMfRP5Nenn+rYxe
NQDtEpGU/rxizwKp8ELpA50e6D5qFRYHvhGTi8nQ47hoOmeMZwh01isdKB0hdp0x
PCrKmVIQ6RILcXRnEGvZurfcqzdzIPGDDKpyLIFf+qVS5FJW7Ct8SKQXjVdfwUpf
bdywbxvkfxL6fUy3FE4gVjm8XXiHXzTTIxmP3MfJSvHod4dtTKNOApQZBLjq1KGo
jpW6R+VoAAUZSekr0Y9L8ohGf0x4NnBgkXorEGotJly3iRaRxAkKKK+b3+wVO8Zy
1h53KWMxU/vaqWokIMTzJnnMHfOPEROu/KUU2Zj5h5k6XnYgGDqQuHLLhH5ATDuK
qQV5dwTabs59ZTP6FCWagqswHQo3LSJffvU47enqq1CoCgwKmSX4y1TqXN0T7VVO
KvnE4K3WlNtbu5e1rBb8/bsbDBAXId1lb+ffJTkVLcX+5kgY9esv7rbxAKzxF+wZ
wm/ZfOD+h7vuSrAe8qt4/NU+C7db8lHaaZ/DJANJDJvlma9dMQCQf0uFvf9qG0jj
crWy3j72DoJcehJDd7H381qDu+AJCKIGYpMUkPhDoRWaDtmo7a8CQBY1E5WNgHCY
TTNz2dWQb47RI/Gqy1nUZc7VJp8PBXsR5pVcqu9ww+XtFYFQvImACYh64Xu3wWbt
BToll9I4yhuMTTd1X77e6+f5lOIqDPVgHmqmDyqD35b5ONVEK8n1iwU1Vh9aiFmp
trj+IZ4408i5u5y+LeHUOycrW4bQxE8JX8+ANvFXHVZ275IIxLKrzy6bJmxWkJnh
h1Chd6sf1Aad6YzBmHt7f+K5GU4zjEmIs0Kd2X+nNfHIM1SbBy8Cvu8Gf44SBUv3
sH3ZmlYZbUnaAGYYciY6nf53XY4APe38FG2uSx0vJcbnOdgzdjrI2G+kaw5dyIhx
2R8rcr6e+AQT5nJ1kBBIjKYyldJ528yl5JyRbH4uo5lAQFwCeeK+b7Ztvp4nADCv
8pUXH+Wo21u/CI9yRQlwjAS6oD/m9nSLErruWZWl0VA/jOx+JX5gF4G8NjfGdqaz
tScqBqlWFGCtvKULaXNUU+R/G6bPLXwHHpy99X6ruVTemv6GRL94lZ6rKVP7a0OI
t3vYmWRs3ybn6YF90HDsNQaDMwGgqn5wwE0SMX109rkr8TznXS5WyLY3G6mIBr7W
TLHD7O6N8usjy8hER+nI16XsDB9GegPMnu2Ofzs5TK1wDXg72hUJrFyGFjPa5ysh
Yu1iu2AYV+KeHy6OeLTI349ScPSHjhzu1RmlB1IhgiU24ufPtxeWz74BHiBS7YIt
ERMJjjwsWmr0TGQ3WJYhGLGkm6HmkLN50MoCEY23aJfQjpr3kiL1bXpK+ynFcPNd
Qr7G7fspnhtmVH9Zy5YbXHCriJm/nMNhz+RrV6T6eYKaMOPflpj7oXwF0qzzIA2N
pbzOHpPvdzNU9Ej2VnLS8Tz0rSwq3LHACtUBBjHgeclLh5pM517CWu7kWpiDztFi
U9XDtR70Tcn3Cy5x8ivOTi8dT0d2Y/G+oCAkrWXtNWJxW78G1NX60HvZ57b4W9XF
QIcNw4juAC/hDvj0liJ/apdXxh1EKzLkvas0Py4UdmHGzB/1OciimKSseKkbNgtB
s8duMpeZ3Hequ1ZdDzR5SZSaU/x5b3htQti1Usvecav0HjEvbekyA4skxvsTNsCY
3uQz0CknkUsdGApXEaUIbScWtofhKg5mPqsNUPz64uh/4gsfnpdqe/DYe44rtnqa
92MUqXaQJ0M6456ds82swRdbGyv2rLOjwchvLaSYmgncGn/ZrBkq8Fw+M27YSLN+
wEgYHsTr0KI1iKjng81p6MeXM0GfmNy3En7QGFuhsdkaZ48JHX9qOQkMGDy1ptIm
wF0C4wm40UwTdR1obcKQSAt+ZiHVw1/KhaHzanm2quj8i0Ddf55hvrCJx6xEliQW
1EiLMw866JuNm5tmyiVm0dI6o94WG7hfeglTmCBmHrFVbzCSZCJ5WRy7Lyppckx+
q/Z82pMaEuJTH4EvrWNrTOXUd9QiDowO8/+cXqEYeBBSsQbfEfpURGlxRo1YvGIB
eZMlnz++4XK2CCuobAQhKmtqbIzo+K9RbkISE11Zl0EVrL/DzEkDaDmE6RQbto+R
Fpr1mE+DYGenoh8aDGEe5vZtantlBsM8TfMxmLxbXLxG5wTmU9xf/ighj4kjan/P
M0Vk2g6WfmQRmOEXTKZFdyhfw4heU6X/rZ8R3lwxfaL6cjlq21WGI9EBAQs9WEPv
xN3VenFmm9eQgktDdd41/usvWrnFPoCJIZ0J5lV3Ssg+hYbyYqz+7vnBkEHti1TG
An/kZGNxilwagsY8l1cUhOg1XRWZE6ZItrAx2aKaRUf0aFbf5Hj42372lJtUSMaS
LPeQbpA+E34QnGq/GWiRjOlzgPiG3OjMl3df7Zlw58XCEL35UGQLr72CxAxSv8K1
IIb2fAcGtYpw8NaOuZAe3qg8vu/sIp9x6luRqEV1kQzoJTlpO6ujsSumfbLckXJW
JMljxMae5O+CXpzCPvogX0WgDyJfJAF2ifhsu3lGyWu1RjrtKsGuX6vDqVQgox3J
/FtJf2CoxJGhx0/McmIdKr+/XSrYwhj+RUXmDXHheD12jC+Jygkrsi7eYGsRb+5I
BUnCTgZLd/QFiBhIJODdWGpTWnw9Yon5AVDch/lDZWY1O/5+fnrKeXspz4m9Wp7Q
umgucEGXHy1SU9eGPVsnsjKpJUpP2AexMJEN+nzJk3G8GSODAN3/OeAHKUpTvjH+
Bf82JyznIgZhJwYe0qlwb5yvKAmIStU4oWBqCEjRqT2ipfd/ydfC/CP5NEevmYba
izxCagPgKLJD8BYiJG6SjSeDKko+MaAQex+xev5yw17FzxRoapWOcpnTjJKjHIRH
+tQH45Ux+11u7X4f6aidAJR3whxfBocRH8MtxjLVT5sCAV68DZaxXC1c+bI2yZjb
24KcFusyW4mw/rzyZQnRzhR51gYQTtuyvnJtfFv+yp8X5gVgFMnjj7SdODYCNe1j
X0qbJG/wm9iX2HzSZnFXR7Jiohzl7LmoYMvhY14VeXdnP1Enm7csV2JF3yVkz5cH
+rPmCGBx935Nh8jDmIYCmDzcpfgG503raUZAJAGToCAMq4gfkgyVMEElJ+NW67Y7
BUvdzRq7NbwZWNd9fqzmZF0C7bs1DoGfJcFVuoLyuHI/6nj76RsPWMSkKg2UmCX5
yMG94/o6Dl5IqLLZdurwbcwE7Qj0MfW+5762KvnEuTAWhm9O6pkUK8aIMviLiA4J
OxdlQdQDHKA0PMDujqDYPWtl3XhEr2ksBcqhbsfyeFFLrlAGr16hdexVeJ35BjBF
7TXJTfjQRtlQOg1QwaBzy6AMIoMOfDfZwJpsWt4vQU61YNZjw6l+kAcraVlCpNaZ
0S3foygyXkbKQQgCvZRbS9Eap4N4KjyZW4idIYkoRmUNWe2feQhyJPJeqG8uaTxr
iohjgme4RlXX8otQ2Dt5wHhm/fQdkS6CfS27SMVgL2D51R9Q1PhsVMVC4ZCZXCxF
hnyZJDUH30TE85sGLk4H9cqjBIDLasNVSLOoyj1lYVN6ldqcgwOMNYtw4b7gbP87
sRN+32T9bpIqdQquUtEYTXZmrD/pMH6QB5jQts8i+bg8MrM2KESOQjQxv+9ZuUZd
syIhVCfVRHiOBi9/RZ312f4fxD2v0xahu5pfTDKZMYUPNVzNgFkv0sHJBjyG/293
ZhFQf4KnQpPABj4qJDlGoxMsOVsJyQeZ+GwXFXcpIuwZ8PyQUSa1XHE5VoDXSYdx
ozvBNb8OrLoauW2iM7/rTW9cDEFfQSRgFHXL3cixcjpnf/QpL8Lc1aGoWnA0UbBR
ZIHMs3MThnMjR+h7M8p8PBNI+eZwNPQ8CeTv+aa+qZ25Q4CatmBwz+XAop9T+/6r
6Md4/6DIDPtPlA0A2A2fnl0qrX65ska7Fm+3jfpC+Par8u1aVbHGZHwHBTqU0GEF
UYVtTykFMNBNpS3fidkMNNMx9LfUPeBmdDTsd91wUIyYaOMYL4RKrpsB9y+e5Zuv
WLIJXfpYibfUoDq11C9LkldRTXG+2QbqOAOiBGQtHBW3fDgPDpX4AhUdAuR5ymcg
jYAhwLvGXyCe+1IOxDFVzQ/hTwmNbciTEWNMCpvtp0Pzgg71pzDkBvGmFlOXjyhS
Nx9LWj56vAAVVSREwEc1BGi6fuJvV2/6wy7PTg+RgwY0qhH/K0oxL1QujZ6J1GW/
CtUF5/CKDMDLa84TMHDyeM3dJRIm2G7sZW6Sf5JZvGdS54uh7md0Z/YHVMrZRBiY
0/OsH26KYhvrEg0FPeDPAmO47XSWkZ4qhJRyOMEwRbdUmzYb5WlgguvtD7R7Mtjx
go8P+sl2q+TK1M4LUXe9RFSqai3Yn0AJQ6Mq7GJn1YzI1aMcPyvDGBuBRejEqvMA
GkA4MnVC41j1v4DUA7p/AHETYqDCNwzMQTiSW3IpjB9lZqOroM/eHp8Ja3ekGd3S
8NzC/6PBpEzV0HkkuA2Ah2XvTKEeI42/QILKYmQ/XdjM/MpeXR7u0sngEZkLuKuX
/C+n7tqPRK6O5NBjcc3Q0BkFLZgGPk80mkIoA4+G4oc/alOLaJgEmX0IG2VhGP+A
S4p2U55TOwJ/47qH5IN74e+2RJSOGn144d2Tkm0CAB1OEOnsfGYxuU5HWirYjq5e
tYgqNZG1nDr2bEmm2zSSwxh3QnMVPx6gBipIIdNYw195hvmNcaq1m/vCZPnfO2r1
rixJmYV5cHdEKvkNUrcdJe+UxGVqx8POLSeMDB81mqAjuktk8wL4yhAzm/W2aeVq
b5/BH1eBglA+82P5INsGDSDm+PpfnwD+VwtToM8gJPs1s1CyC8IFyNslAwgNWxzM
685WW/Tsk7fX1msz4GuJWcTxCgCLXifsl+IVy0PG5Iu94cLLYwz8EFXuis6QfSmf
swFaL2Yeb+6D8Q9ysECm+bjoNtygMQDcIZ1875lv4lUHpbvNWPBgIuRpvQpqAPro
k3Psh2kn1HoOrVx+bxT/stXjKanpjBtkFXhXuCNqX5608UUsvhnXzzxFfSgMDt+z
x5HrfopMI/D4iBWjsyH4uivbLR5nobDkE+PRLTg7wlOATTR0XqxidLIHzE0Lq5KS
Wzk0RsTrpBK1+c9OJE1uBd1SgVleTTbopwFzio8DPa6gETLL9I8Rq4teZfJHEfCh
3d3oC0LiqAyJnw+j3SWku1uLQQJS3gUTTORwg+s4nuKJ64NQgFrTInbyjxzAa1c4
su8J4qiQthpTZTzMHtBqXT70cqiKSEpvJj8uoqCmTrKXBINT/RSVERVdfIcxzT07
CImviXE7mtZ37glpo5dM3qVPcpnRx7sM3CJCXfaxerbxc8BsNuxypkcGvfKgje8x
rNa06YGydso9TwvlfSUnt1KicRXfIy5VIiFe5IANZDDv7iUiBelwQnAvqXA3uCrl
jrlY8eD+7n6MjrokuiRHDcxwUMaF8jRDKcHz4Ws2dDpHlb/Tn5N32PGL1CcQPPHF
lzNyvJynOmyqixrv7ew8dN986Tw3jjwHgdaqRzPeSHwBvVc7A6xtJbVG/TwbOKae
gCxSmuy1/hrkET6nPHSa/hXUOAePgRSV4UyvLeognJUXWiipAdZHDaEe97B/tWAZ
ciSYAm7ZqGwQQc9EN6M4zQaAq9kcS+pQJUA2lq4fqqImNfboKZ9hJ3lBEErzHwY2
7SZ6377c+ArSkk07g/hLeZ2olAAYmVe9lR9OUd20Tkgz12ekXYRVTY11iY1YBwJb
locXAR+yeM00oeERQhlGTtHjL7DJzPHxvMNb/Ug+V37vsVVXVer+mNYbpA8fGZCf
dsf3qaytraDPwLMNbE/yP49+9wH88/rLMM2Pg00YDfJDMiz3VT/PUh1z5MwTiKrB
I8v3JQKVYW6EJL7RICaB81Wpgd8wDeRaVQLSY5MvJmONoUixICjP6eeo40FHLUJl
QA6jxwTW450UvaHyyfJ0Pc76k41wNVvgsDQkHyaij4rVFon0d1OEhc+2FFQ0gabr
GL7Q/aH0TXE0PMht6eVy7DCCsa09Sa+gmcyujRRqk0ohKTSxlNOiz8Z+TLkZj1w3
rQhnT491Ah5oz1145+MZjfSPYFN4iFVn2MS20faQH+Qu3xe2FmLH914IsjcENj3A
eROgrWhDfLKr3ZFWixpaf3eaBrMGswVbQnxKbHZWKItSKCUNWiwmWGtKJTdNDp75
21CpJeiCLwmcWJx5I0EH8Yzd/ibJJN6qFMHmwsa0hufAQbZHQMYxUqXIBffWL0YS
dxRRxzipuy6NkKq7hZCggLORrAVxRBhqnOaWscysirXApkMELVpcdg3CdYpJwS//
n5qr74hOeinEK62gDCzLcX0D6phii5Rg6cgmTTrhBPrLywLtfOmrcRsYRVlLYpmq
cslC8EclKO4uA5qmC2AtjPJ/F+uhn/3GQHjsVqpNBk+LBTwkNaikBasyBjlRC14v
TbyildRBkDqfthe6aez7JG7orAJ8pdtwoVn1MmmsiMJ6oBzk1lBSMM/r5QEc4T1t
eRyIwH3OVBFx9Z5t3242cUQ1ln/o9gqdX7N+OqP6GDJyE0w+7e67YMj+wuXh6T0y
wcz5IO7vrzdxn+tn2Oyr65nRvHwhZf+PhGwM8fId/I6/8g/QPRQhBEkO/8wjR0Vf
nwrOOWPKKRcxha2IeULX9s5LORrMRNR5W53a2p/zdG4MG064ulBfGOKw80fvqyWu
5hUexzikHlllIpkxlubf4RRs+cX22MdxkTkZpzl4w7W6lN/8Mh11wcCBZpY9uvlC
WabEM1NHy+Rv9gd/VUATQ5abQQ0CK/nAi9Q58bINFvgvjgeVSdYOqOWdHypy/Ex7
S5FfNDyEC3xUiJj/gGoIDPIdJIJRtNUfULoPBbFnhSxaOzMOkGUmuanCvHOU47za
hmCFB+0QKflCUuPY9UftTj2bIMGmUcMDfxOy0mfty4i50doE57HN7qklPxwOUTlV
woXAAPVKH+INkoy3crx8hPWKbKZeMICxtVJWx1myPSur8dB6BqhX9k6DxZ5VTiik
2fdiBBtztbeXFah6BOuqP/41McS5N5uGs9boQGGqwWaXPBFuE66a2LNi/wBRbnqT
GxNXDy5ZTBhZkS/qTDBZakoGQILV5DjwT5vJ84ITciYyRn9kZtbTxhOyXUef3SOI
BvnqDrMIWSYcyZNJV1scblU/945BiFN9R07zAnRVRC85BBXVGFTn3R1CzmNci/Oi
pN7shdcpsMYU8OnuVRJcCDrh8GikEMgSt5vy16CwJmOOTtRH6TXGRydYNJapgtDF
dRPwdv0QIS4tDjz1Xw4bD6v997UgkanH2S8KYluW64cmyFzaPZQdbGo0DU7YjHqX
PrrP7CxcxkAtRPcQAu8mAzwzEKkb9V0Gj5G7B23l894kNrwoxGtW0KfPHZcYjxFZ
VpzLtg6qUm/ynF2bNwp7HZ/rgQxz2N+V8otjG3sRmfGnzsEbWT/cEAxBGDZGAA+I
dXtn7bBSEc8Bs9rjHgx2hzDuwBWRDIjkBQSgbMFa/9r6QGzEIGShiy4prbnOrbOf
qU3dlyCqdv1UxKD1QRRiAZ1miig1OHej4uyOobyAz2m/KA4PbQ6WhHXe65cD75pL
sKtIYunTCAJrPI/mqrOnhHDAZhvRVhfZs3QCuo+PBGpi3w6YM4j1g2X95gvwqdjB
4qlNYHCe43eoWG+iKRPopWsMWs9ym+I7/cVvXPPhE5bVgfxfG60LuuH+f4OijykM
ejnNgexUx5S1Eh3+kKboGL9zb/MD06IhlT9l28H31g3sitiPJHBOH9X6+30xgsQG
ssq26vC2XS1qCIQ16JTD5fIm1TRKGaCl0tDxnPSYFeFd6HtiqnvImqB9MG+RYilR
1gs0RO5J5MimWreVaaF994kUzSA/IdKj8kG1tp5+Ux+gLRLVbf1NhQW2zFw5cTV8
zf0KJhsjQ5t5hgnRapKNNfS3zY0nM//qKczvD+5aLLFmE1Sf6uEAQuBfALxhCVKR
upsgRfaL63ckuUHcdQMDIpNtIwymwio3IAL2Xq8+Z4xDlwXPR0gQPJDnhdvwMrOq
Wqfbo8XUHu5XIPrj98S9MtMvAYEzRgkbZkaEGymgxg7Rz+yww+evJooShOpw8PsB
qdFTeskwBs9zbyNpKE+Z3EXeMt9kY8E7JEBF4dgQlxEeuVCuA8R8wNCtR7XLoMZp
vnqg7e/Epx6WtVTKBKNO//epS5AUcFCl6HEzFFvV0GQtk8cYcZOA2rh9W94xWDUr
zJwFsDbbHEL48A4WeBrVrddk1ooOezUXhq3BgotsllbtpAcVSqTLlQNM6EFkQWLA
SWcIVfF7JbKEQ9Ta6L1LhHL4CuWI2QqMvX4H5KeFagt9+NToQKhG6O+hTQUqYpmK
fYr+HIbOwtQpuBemVJhoBcMSPYj4ydDDWOwrETV5EXYGtNwQUst3e+CtjPYZkTID
dzPGCgZBnebRYUSEW2ZMUsUjHVdvs5JevLZZufMMqPLeCJdYKA+YPSTp8RZ97dfz
1FlygNZkJL0njdqHphSe2Qs2DBzIkZWDMgTsMRrGhYYOcsinP2PQuy8ytZ7JgBT4
tZBiSPvvFR0E9Lglz1W1VWhz2aGtTrGpOCIIVXdfvmvRV8kQxtjhhJZXybeo7N7X
jtI+4PyuZOAhyEliVs0LdXJytQH4OaW1UEowgslUI/Hr3VlF2o2TjHkHezfCsw9h
yZdixytwBnLqbG4DfxjPNe5G2B6PHNuYDJbAhB3pZPBsXi2o2VWJ0BClwrHbW2jq
3+xUJGku/eqcrX04GG+RqUcVBcJtPR3m4fMPakQKAEuJJTN1ljjml/MiUMHZjicN
czMuHLv7y/+pEyfJThUIPi6dVouKgH0qfh55lLxstO4iFJyK6xWaYRSRFV0RyvnI
xGGg5nCvEzDFj0wBKoOkVAMjhUGaCSKFxqTgSx9T0loa3xXqPvwhZBq9dJ9OVTBw
P6Z2yoNkXGAWauKIj115PM5y4sjazqi80LRtL03f+R68hM4+0VZmOHPm1efNHAc9
cQ1zGQ6YopOSdmfkim3KTzFw/iapJWtZNZyW8ILmb4LplaXEgCKfjRqz0EzooTuB
fld7/yC0f/YEXDZKvoqFHY0NhCi6U9O25MPqyEzAh13N9ZGJY+Xwb5SinSyqSNbO
wK3SxejVbnnsSf7t150U+5QPo1JBP03voCaC2YCIM33g0xOiKBmMAXYYvJrAQdKF
jDXfS0EKp8GamheGw2cIhnw5518tyrXbElJZTUrEtC0D6NdACr7YshMRekG54ZNi
Rj0Cf5Nh4iCqJM/LB6MQpx8f3qhOUsxXh26nf/9ILu9nDn6q4XqMBcumHtVkpXPI
xOCxfk4x503Y6XaZKWrqTFAWlSEWvll7bDVJ3M3gOoXTzP8uF27gLgPuxlpYOx9A
UFmcvKNMvR3BiQTz23oq69myUn5EO6W8g7+bDCygo8cwf7E9gNQjWmZklUobSCgl
Y9clhBFQGU9mpk2AUgGLeanTzxchqY65G8WwC5xXGJLCnVhfw2DHzahz9gvY93hs
IXfDyoaZE0BzxkITJ2/5V34Q60srkIY59/6aaHMKh184KufOl2jr0n50AxkGBQUu
dsXbHHnGB/dEjOoqrFpvVL1Ylrj5btJvuxoYhsKAJ7tnR/dFmZnDgbYlpjLR3X+e
qRsD6dIU7nzGrqM0EjTOLovdqWkUh0cCiTxDyZua6y2WVBLzlF60Af2QS+6xKjSA
oczZj8NRDrg2cg3MimkI+wWGj+1YwkbVhifpOh/pDbl4efZqIFreaDcnJ3Pqa6Lm
tXVUkyUDQgqhrKU1aJAHmYoTnPpha7ImrQx9ylijyEziKNX0cZnaWYhX1kkGrB4M
TLMqu6fw8bOPwkh/LZ5b4zDM6Mu/XPnuTyggC9td7u+KR5udxPR57C7708n3KcRJ
/wS6bDyV7AdBCRIVz+MGsMyj4TAgAEiTP1cUihKCWnjUyFKsW/nUGQ3Si0giic5+
Gurct6J77M30xDDJIzq0LZUGDiqIYrXxhpCSLL9KcSP4l5c5MK6Q7JlTLrvA5H3u
38O+24e4DPNDIm1J+eGNcnUdHwONAVcGY3ns9T3uuBaN8R1mhRD1odKuz3TnU4uG
oFPL58AQcArlzSdW2Xg7/NHfNwD/dDm8AWc0TwQC97zr/A1Pj7M7FiBcZ2ERb00d
unEuD/D9dByuzsc4DqbRa6udKPuXhwMqwCkjVeqnuxeBK3aUBA/tuda/JG+zKWvN
hu+AysVRUA82Kle2g2jobL/3j2g8lhqyrqmGXIVupNfnSK4px3v5Xr8vnpzmmS1t
a4PrAM7+ttSu2rLTBp5VBgvojMBqFKRjakYotXE/9qhCAxjHUU+JJBR902ebNPVu
lH1g/PhaMm+IkKnaD+kkE+ptBUZM94fg9f8/ouxG2hSnVYIcy+UO3g5/s/x4tnFY
lbaxj/nhv2SBg4CO3fWgbPhwKABzEYbh+AFe8dO3aSApWCPXz1EABtchGyJ5fJD0
8fYSSZyF2K7Lg+ZOSTKHWkbVbeDo/aiRJB1V5yj9ZpJCalkQN7sF7Fvscngm2UZ1
9MG+MzjpwzFgoxAofXtVGK8qDKdMLCbQciI5bx6uhHUVbRAHo2aW8pphzDBoZnnZ
UFFZh9AMwYWU7Nw1zw8pn5bulzHlfHq+JGVNQPRmCxpCu0rIqU2ZO04DjYVcMHds
gc+qrsKWX5+bdXculJX531xyMJ9zmiYZhhNTyTxlLozPMuQTRWLeNMtPqWbBkx8j
qqCKUZE9asgQ9B86E7eV8llW2EB4xOQmSB26KLO0TM8z3ieti5bNr1QS/8ABf56E
jRP6Sd5YasnCGVm4HPj69lSXwEMH2tVWvC0YCL6QcW4F0zsdZkta0i/R18bWsekP
ozNV6xI6ar+rIIPlQLwVA/pfBjMDs01kh8GRPDWPGf7XMeBDJTJ5ocvy6S+Vphz7
qfK0HTpDDlH4VvhjPkklw6yNCYeQX8xGkqqbql/N36HDpyfkhYPktpRDYzA8tXqm
UXiF/SEgDQB60NbcgR9OS9cParohYgud2eny9uzSDP8gsCJZGg7jvyq353wmGLBp
TAuNjwuOAonXWo58Pm7iY0J/t1UXDWMaHEDnWUaTlOdKdhPuUCH4xu4rT8C4regR
vz9tocqwEGvr1dxW/tFZ4NWs5XRax+K89AUewNu1Lxuo9jCapu2C8xWf281VFqY0
b5260V0m7su4r2sWOVwJw0D0+CPodURNnQDYgKPitXudHJl9F9r6Fddn8fbvP0Wm
BnNoe+r5JRM16/3mzEkxTP0wILG+M3FsX27qGSiXsQtZaZM1SBuLs8yEhmO6oXVd
sn59DUlraHfd9MA987KU6YNFKcs0mhXGCYlpHbc0AV/uR0fqaDU/Qrn1l7F5MFBL
1K4qUnMiBlJncWMbn2NCOzyWKon3aryvU+G/LEOTpJfSfyPHZrbyopkBOxeNsWuN
yuOR6G6TO4MKAwD0k4Qsj7TgnpnUHNVON2SV6vwrZTV5dsuH9kSE2CC+nIUbHXDi
BwukwnyOgvBYxUtIEtEvz7dZymTyDWw+Y9bVueFPTfStAifBTh1QN+x6Xiv/YyNX
6btu4BIYnUwMvjDA9pO/lo2bqsBlKXbXz3N9yB8DZ9siK9ielI42q6p+oLvN3f42
En96ne3wmijZ57/C/gUm2wlm2ZGlfs2Ijq/NjltygEeB5lC+FhAFUIcArphHrahz
MGR6mDDHdivJmr/ySNQZl5P2HRnJyHCPcgdi0HraP16rAT4oGpziWThAtGp5yopa
RDGLy+VQC/O9S7LMMIu+hXGF0D8uZe2EHjIa63qNbXMxkuO9QGX/NXd6q1oGtcq6
XH7W++g04dpILc57iD8T41ISMGEnLAkexzo8m77YmOK4WRShkrjp2YAJKpGisxcr
QKc8YHh5wpRftVTCoBRHUUfx33oOM7NGoRdx7ecFFjWqMFARAKFahHMFb5HR7iBL
7Gm1HldlHweDIR5zrk7PvKXY3JwaC6/DSaNT+83znSQyLAtuSNuMdcarBBO1d6wA
RbUJIQkHbhJsVHCiwA+fXh71sOXwEKGBF3LfClRLT7g/OFkHjJxGGosMKYVKKXtC
Hp5eKzjMYwdml3LiMhJ4pMJAFpqccqg85ygaqi6RX5BESkFSm7WHcN1Da+/DcSww
hL05N7QdZreQG6b58udNq4+JuIT52UgX+OZDiEQ07AvuFv9ixIWs6EJqzHEFUvE0
tekzsKLSFAnTTC+xv8uuXpbDffw245LOaNx/ApooYLGPBQQEjpF1ohTz9zkoCH2d
sudUDjcx9KQh24z/48k5kzHaqibV3ZUWKQ6IvAY3ATU9anyowQx8jVII25VH2gAF
VGQyPK4VmuIeSDMcayZI+WsM1+ofPnrS6v+rU86TlSe9OqlMD+emxsfphhlgwT/m
r6E+Tvv8SmjKPxswe+UD889rco/l+M2gwQbVQWxnw0sbd0Bl7nWw1lYNQcuMaO+F
/8C/ANWTkZk4zCW83+Qf0+jF3+shGD4NTgCXx/A2vaVZckKxGz63S8CBkPvwqegw
i6hm1bvRjwStEjR3ROzRC+83LDXmeGV3xln2zs1s1SPY16urE5bgzvt5qZE8KUJR
MoMRXQci52juCnzGQbknFyBk+dNLTbPnXi4uUXF1c9j6xZmPW9jqbt08ZrIlXvCN
OxkP2IQEUhpcZkOd0nWVhA29j8w/qTlrAs4uc3FZSTcN2IP8+mEJIlBXz2gh3vbF
6gqq0deAX9+oRDUaSLoaSav1XT77oHFtzpi+RExAEKOcrIvuEYt0OwhHu/5T8Ncc
INY7rjAWhohaOb5twSoMym5nRcze1uAvwaOkmwejYUz58nEl8Lz9sxddkSyUzTg3
HmNLu0Ydgnu4XzIYKylE+JTcd6N4E01+n5YFjU2XGqJyYvUcV7BV7TRCWTCbAcaA
UM/uSOuVP3XI82mstGEGavhKh0lwOMAK3NjaONgTe7uUSIjiwLFUPiKtXqx62AJ2
PiWuD4nbWI1cD38F1CCVVDommvzvhsz3H4MQjb0W0J5EZ087l8xYJHkX3723yLcP
2xt7U4z55giFtjybxUGOL1F4uqlTzM7wHUOWdVCgHg59ElqLs3WsH4z9xtCV4n7i
k79cWGq1KbjsfcCqUmJFzZdvYdMYmzIoOpHWyq7JS+jT8EJSbRktJiMuTACaH84Y
+udA1XP4inYCJVnxl6ZYLK+O/U7/283FOJuQBoBVOtcCPmIJyotuJ7OvCpG2xOoK
I2vbKDWDPFcTNkZl6FiulBgyUIbT2l2SfWFpGjY0EmsAGK/ioBmEKXk7526A4a7T
JJCLFkZ4nZxrhLWnG/wHwnKz3rJGbK5OUJ5ML6sQlBdtDOssc+ad6d9B3+FWWNgq
75ZBn5YYc85GXEzaUQb2qNGKqCxO42Gp3UujBBVQ1Z+I0qQ+m5oguBpi4pP/I/ZN
2d6nhszCY7I3qFpwJpCfnXg65F+aWj+wW+OZ596+rpOO+LWNwizvanaLSX00WhmC
L0Nwy0MzjyWeR0BDF/mF7Z9yiKny5txP6COjvqZqP/GmuVdu7Pd0JAsvsbEgOpAE
1GFMzCiCg8fXcNfd1chQncx0CJGxDlDicRKKFAUjouk0nvEhuQe+IdUPTz9EpaxX
O8AKYttuJF37XdqoQgxybD4bat+DxHDFy6sn/RQg0Damh2l6SFH5rvq4fAc6JjO4
YEeU6fiyIfpWs+ah+CPXhn5H5HLV9IWaRYVEVIy3KvpqCBvx/REMHefUsRzBQaDv
grbLI1ZEt/4+HZqCgRVSt6O7MjbXVwf7ktN++baFiFj+QMX+xToL0YAb/Na6Syqi
cPNf04RZoFojDQ2IGqDHyrOkRKFLYKVwx7ezJMiXThSWTaBVnkiEi9pJ5xo9HO5l
DJPUgsdhZKzcnHYFWka4ZGBekeow4NMLbO5v/yucpuYZ82XP652K6sl6UI/Ad9Ij
V4CeECu3WixZNg/UQ1lik9v5FFP00IheTdZj6I3Zh96LXQj6L6Cuus1Odj47sOrY
3syc4M1NPKSXF5Cn99j1fRygXfFHsR3HvL5sKnit/N+Uh/XpdmA7WiBM+6r64zjp
7exHe9O93LxfKocJRwtKgIyUfRcFXJTAXAztA9bTl27izn9AyTGqRz8ePxLDoi4O
kCCxRf7J0sdSQJLArO+gDmUPa9TOIuA7walrKumG8/faVNlCVacM4yhjALuJ+blW
n83M6mp99X/4zSlp+vpKfwOmLnhQlcERrrxDe/u/IHKkLTI2c6mBu/8qjD08frGA
ALq/boFgjIXL3fVbcVSDT55QnytYu5ZmZEH4dN0G2rUHlUdAlPFpxoUrIXrKLUxM
C18eezSLczbupeiSa86gJasQmWO7SPaykqzJgTwUF5ztTm9XZoKi0l9STdl4lhKM
glNSk9D8elZhmuoQZzyETlI93rwApWbbYgAcO7gXdIe4B3vWyngt4Dl0NuZeBuNe
I198dIwQ0KNy9GkVlz8GnxoubxjeVvxdAc/DA6Aa2bcqcrKN1gYOz/bWgHYQCLkv
2kw5yfR4LmzbShSKlL+1l1hzmtzJgZ5EE1t5cmHxdbCxVMi7SP3DhUvsD+gpEU8v
RuQstGt87c5l1jmwA+TprM6NNzKNmCn0NPa5TmdZwLd5NnLs0c6LtelqXkvZJxDS
SiFFWKeMf8o+SgkmDthiHc//BVcLi6kH3Lc3X0SGM2UbnGii/auxuD1etaAA75MI
hFNB7o4QyfBWvT1IDzeuwAj3adzDSWg5L21/2zrrMhCMGiV/EXoMv9fXxPuExK9V
YaR+ep9HDvt9WH/gfR+0aFMfZUM6CxiKRSeA1ZDdMMR4NF+jQHPlluGfVVpfboi2
jWN/qCWUVBwGbZQh/HXG4m0fFPzvgpLuoR5qvbtN8gAtonU4e8lwVl488UOZLDdC
iCYi8vB4ieham1+B0j/l2r4rmyNatUjfaw7jqQmITCd28FVewX4ynsfJOCZcFvJD
lddzSWoLOiwsEEgJUmj6zM60varIKrvfLhai4mwJ/c6OrBtcGhpdGQPF8kGpy/bg
YYMrfCjxJWJGkV0lS7WsZxmYSmTbu+L+pjYx3IEuhtr6vwxR/VyRDrsEO4AkzAmq
nL7J2FZwXVuZz3WrUwN83yEHnfMZc+kpgbweI3Hpx2+kHxLWsqq42fR0q/Yd23Fq
cykJ0hCksaFQafCGRslV0Nw+vxoGOMrs498vjNmirLn3jqh501EdijayqYYUMFGS
3JMl+xuEDAtwdS9KjDJpqxsm3oGSyEeBSCsD1Qix8lUtodPQ31x/wIa3GcPalvr3
UhkF2q2cY4QXV3TRVMP2t4uaf193lOQBEXORiPiZvCUCdEDBQdsSP1jVan6OLAd/
9zOjODac6cNjEmGdQk1/zNotgfac/fYSJmWA7MThbVvKhJ8TTK3qC5F1AcEcTbcm
Wjn8Q9x9I51dJXcOctYVzMF3pcNMir3H2f9i5yB/0/ahI52lU40hVi/FVo/mGwvT
ybscokP9afxATPwAKNzo9LFHCTBKqAKtNQ/8H5qdIvyAx0Kp/n3E7UMox7YGGZtI
KeiS0aaSgw3E7YAlRprVp8fNd1Q9TSY2Dt/SLJ6dALRnyKL/RO1y6dKnINdK3qhw
yIaWj5Ht2PIMNCc1+khaCh3OfO004M1od90IIuLLnEb9JL3zhNdBGVgBScGtSiHg
/Y8yMnZckinMXAPqPYoX3ZSIbJjgMC4POJs1q6gz/fgYl12iMJ0g2uQJcNtbN94y
qhLULzXefwUBFxK45Vt0FpjLaaLWboe/ErgxJAYWl2Q6wIGlLZcCYh+itmaTcQlV
tcKr1Z8vGTA3EvmuCuHdIZ68U2ASXTgnMtGnYl8cWpF1nLtFK4CdjRbYnc1BPqvU
8aZN5tEAZcyXKXpIC4nScz+JG7tIyZSiX1yXdnhBX+5d15uM1LNGBx2vp2yoSmUh
tH3FCXhSqtcKm4hFSrCzZycpNATlAgTNLbI9erkvtb3dr0489hMnPo6HEdURYtoK
wcGUs5kO8avDLapFi82IsCQU7xe6x2KNf3hPQ8CHA44QHjvpyhfCgs0eGE9HlxSb
579RkyguotnjV2Nl7vgPACFgiSW3GqVQeG8f4U4XNz9kpIu3b1MkO0u6E7RD/GH0
dePaZTksWFil7pz9z5Upjc3RPNB///59yw5Jy9zyl8Xg3Vd7C8CkE9e0vQdPmybI
j4yFGfAhPefL+doW69ROO8KNefOqpJcrhfZ1o8mc7V+0awB2A1T9XOYZrMsv2za5
5vSoXLkG/DYNA81rvCc1cGfmU/KTT0FDxY+ZJp6gDbirrbuCDskfCxB07nzEug2p
kuFI/ZYqevW01kM96F0y8d1GCRP52hK8sgYLQpT6CxS8uKDoaNVIBAh+UtytDZPc
MDfb++k50YP4S8q3GyBIK1/T7qKqJMjqgFW1hy7mZ+tJIg6B/f+l2A9B69xC4Zzl
Tcp6AGrvGU+kGkZvkxXIfRGh3iOVwrhih1PGpQ1Gpph1NWHeNCcrvYrHNIIYA7Ak
Afo++M+Wm5cPvHdJX7IouZ/hrFrg/YrWreb6XY9yrMMtzWQrS0uPo+/6WI0C/E1J
IcOqHDtLBS0L4j2GZT1IeERKKNZUNyNnTVQNVIPjbRCg45QxLggdOONpDlvccWw0
A7iletlP8dZgLo1UEC+VtTunH5nVjeY0pKu1QmS0tFm2uRVGki32d00AR3RhdzIe
CL0Fmk6iej4R49QbANirGgxwuUzcJqErHeP9NBE6k04UWDChMi+59tnnDvO2EDIE
x/f9+vcpZ7RabnQqc6zqJQhkwLK7/8nQu8PTOGAlK/+F0vuatjuqXJZkyIxl3uDA
zbea6r+5PHftfcQEPBaztIFDP//LbOTy+gIoBb7dVe6jLamx3KMrE2lYEUbSIXsP
mgGTWRZn4V3aYdfBZwBMd4UGZYOedhN/oknrrPVI/O6xK8wSDbtMBse4kUO4tAR8
D65+U93ang8NXm8OupMajNke4RDDmBzF7d2bOs5VeylZfp4ThM1PlPZQpX+Dicq6
V4xf4/jxREv4IXOmVg1A0P07rQxCQ+yZqCASkoa6/DTBgCGm7mGmvBhMCJ+HT144
/2lEIoja44h0j+Dwn2Ixlra0tSzrtTVicA7Ni0PmdPgi6BIJhs2O+RMwpA8pH/O8
+VLp6skViasr0Jh80YjhHn1iWhdVhzFoE4PtBWrSJ5aVt6nLqKjvD+DINZ3TBAZT
TmCDzBZBrwYNmSr2irXAlW6ZOwjMX0mOekdFi+KtUkQx8iTLNinpgyusn03IW/kx
uG2KHYKPWsuEFcr9tgcCF1IoUxNgvKmLICH6sFtim7I5orjfxwXeoO3q1CD5g0uD
DZUkzs6fJ6VaYZqRN+gHlA7clG3g2AAtW0hjUn1EErfQGZDod3u4MQAL50V5MU3k
vATOy+beVDz66fN7HNYGtVmFhm2JgNATua/7Zh3KfwX8DnQSMZZAJMJoznGU+KM5
aswk70MHZEjhAqIoEyCJSsUM0+1cT92qnEmED+a+b/C4tE/iUGZ9vIHvjVVW9iBh
eHPiSPv4Kltpgp9dnLL5Z4o1Deo22xg5CJU7P4FW8XoeEXKY8PyW0bUpFbQHj4ar
AE+cvOMgR3hVEAE1AVwa1Rg13BvMR2+FoL7+H66njPSFOY/KSfN0fJ7CyrBCJUCK
Y++SfnlTno01rXvYY8j7hB1kuMTvJ5npZWYrJ0dhiyvNp12cPHtnUFSnJglJQOpO
OP+syzpGY3Lbon9FFTkFsbbSGZI8ohJUVh01FjQZE/0D0/rIC6ceFViqzON/ElV4
1iRje077mYUAvy2+YyzxakNK200shD3w4Dvk1gFNZFmy2jkZCyRV0+Eur6POcnX8
p46/pC3R5pyC1jYbFUVqpnv0iUf7DLWPrCTrDmLm3snXVp61NC0CDZfWHds8t0uP
Wc7qgmIORgHP/Vd4YC9q3zWjVSQpxn578hvhJYWxH5zkGqR398I16A+Ixy4a9Fbe
FISAzPNguoHvuW0VdwkuZ9KDQurzL0b0IbL0G5EynUWRm174E1fb2HtqR2Vd62BO
9lFzyJ55+DqC9ecfLbXjYQ3rQn31Q5uR69GoLAi66wRQgGEOHHIu+kfsCxhkiWw/
PM/cpDaHSX2DCWzQxRY7WHxZne5sX/eorAFffeHjrDQEZfBRwL1GipFLwTBGAvQb
HKb0RyFDhpFMpru1gp1He4advxoDJSW5MTp5Ehf1YWYuHV/R2cW0op8tJNSQamX5
l99QoIK5oSTq8Rm4bVnt7u7ZyWOut+7Lt48zANgFghCy2oJDgykBXsiKOVnijeYU
eYt1HjGBwosSs1HOPDxIag6dXS4fsXhHP53gkAJthECMDYqVDJq+re6tHOh49juD
Gc/FBuSb791NMX3PykjAKyIzAgySpMjp9LSs14OGLwdBmrFXBHsJS74azeY7BD8J
xDLM7F+qJ3cnHrmbLr+ZvfN6ux8m8C0yVxIM+Iik0PW2r3NC6yrGWefM8e2QUh9Q
KAI6OBbbYVj/41FZhr/E+3FkUVQLxmsRGJcX6AZSxWSbSZHXFyvPGv0sprSns+mJ
tdsttJGmJVmBH/PApMrWxPvCOHRgtNnjYqub0zXw18x4PhKivn5u/iiGN7GP2k+z
Sgtu0vBFMRI8efZ9ECI7qBVMLx1B11vq1ost+tWP3/mZkkMRZhwkubZxrqwpSMgx
FeL6QDus2SJYV5RA46Jw/fznwbvvUbi+bFBaTnHtVQHi1PwJL0wvwV8r9xHh41HW
KbyhrJnzftgDsqhRZnM5ZtiK0bkcz7V55xBmM9h1EC3HTUJwJ4qIQLIBOTOzUrh3
8dOuEKyv+nIHHYyLoiHMKpVKoaP8+/rHbBO5bHbfPZOnrtNNEvVLvuLPJWP4DFp+
KqCP/6Bq899dR2/AmvJOX+tjJTbSKsLge839PqvumhxYbNr/7CWJB/f+KD+RWj9c
7omJfRcooDXVGUt04r8Ujo5+Zig1uKc+PA6rWzr3dBNLI4s6WE4CyKYW5i72pzhJ
vF7VoVG9BsiDkN8LcfNInNz/ykPptoYeuvVUdLBva1UJkkWDUZFyCNMFnGmu1kIC
12ZqCgJLAAhjn4waU0NGIG6iAP3hIUE/j6AS4eYbfJKXZJDF8FC2E5mM4b0x+YpI
xcEJBHmDyyGMkdgHh/K1+Q7idiWxOZPT+Kt4QgpCjR4XafhVfDMaa2WcEhcrk+NN
JlOgbZl3fv8UZ37gOcFdl47sQeRxm3F40FY2jiaOBrrQ0qMSfkSMWHreGYn0r3aV
pe7GLoAnu8wmkWKtwJMfkYg1AXarf/rAtw0oLJSGbMuGLt7BTett4Ognw2Kmv0gV
daaTgdK6v2XuTIRuFMoN0koPzbgXePRKH5j5lVuZeBFqwp2mMYfMR3EJ1InitIO+
zQEfVzNSSQbmIMVwXIcl9PSAl1L+wU5JVhitsbfLIEszelKhP/+/iNY12jR8EanZ
o/hyQsKPxUeqP8Cn2Wd22sySpuYmyWdaiaeJoVAB71FbrZDJjRo8eI1Svt0JxME5
LlJnX7EHN/Ou+IUNLOj+d5LjItJZWakWAy6bz/UEwEM/8lQ5to9j0Inc9OLHSrjQ
DzAJs/jyRfLVX7yJ9p+UyJF55EDy1rJ9/IhmW9syUeh9fzGiLUgdrvfwplodfZHh
aScGg923waV6B9uUzlmilfftqLF/PdFYONBu7EUG/yF3bNeI1JCt/1DPRUgQqeRL
OUe0ys3lTBdZ1zM1tJLwqS9jydvlZ+2yWA85KhbE92jz3ZAYJJiyb2az5ATzf00y
U8H+IXFWQjLf5cD3tiw5f6PTziuDlg0Vua2C4xAHDv2o19ABi5WYf21sHMxw6Zfq
OGj3foEkEbzIvbaOVBB3VW6oYwAns7734v4fY6o1LFEHezY32fsIgo49a460gIa6
iA2Nq1taQC923lPlqajXX30FqKIJ1Zd1mE3zCxykZ0ge4FU8ceLnLYdiLn9Hqept
SfRzKniTAGdD7EUHFwIGaaCi7SBPPR6YU3gD3T5VP33MN92sifjQ8j2cSORPIK8q
UEY+Rtl8ssDI0gYhudY2hErP+tfNn7OZkKLcKsu9doDuSKYaAtToLPG6njnSq7Wj
dmsoG9DUoq7uQQ9yzr9iUiPxxL3+e6s/AGv+KtqMM7W3yTN6biVimihjfypMTllm
FmFbZ6TYuqoSFojpqgEFThMEIFpu045TfdUZbvXT986dbVl/RVLf1gdljAj+ctTp
1NVbMDxQtxuk/8NUUZFkJFhdGNDt5TjS+/rFRSO4Ou/wOPloKtqW1zo6iuCu2IXL
fzhYyyHIrpt4wlNSY6A9IVurbrOt2x7rR3uzqmAno+SMDyTrUIDbRU3tuB01yjPk
T6im+1hU8rZbfhCfC8qDKRBM537hAt4/8fB3SeVs8oRmoJvor4RftYUWHv43WKcy
8x1F65Nnm7q08hlg3W5P+ApWI493xxNnIZWJOTe1cJXuHkGZXnm7zjAfIc8qLaVY
evQREwBa5LYO40VkDQzLXeD/adcjoPpeDa+TTXPqTpotm2+UncIWbHI2IanOZyA9
BhS4+bYRkUYnfjFWaIZ8VgxsBXZy4gYoEfoCr4MbFsZE/jnmCUVLEKDJFll+8vYs
Ur+jZH+vmcN5QOjxfrj9M2IA53ehNb4wTyIk6dkelhwcQAuEhlwoTNrJoXgnyJF2
twv0EVapgJZK+QGLKoVD0HwlVgt3iWEoOH8utOt8SIo2DaaWcrx03HFLoYnwwfii
BQV9R6L3fyZkO3d6UPsCtqVfBiNxBHBfSPgfthNdrRDc4RJIzEJ2umFNFX9nRlKc
9oQcHf4EaVL74BZY3hNYbeVLBORhj1Kp9HP/FJQY6b1+DknFcgejSUlg+d30+etk
4nP82YS8jirRcOK66znUdBpbm2YX57sZ7Nmn3zKPRjKh7NQK5zxUO5n9nPtoedd0
7TBhWuUIpOj7vp4chV50tTOK6p1TI+RSnFCj/JnzIpqcv+27xOK5TQ8iUuKvt27o
KX9FX3rf+SxnClrxhycCoHH9i8KfJnKUAv5hRV2WdTU5two7npFpAKGaSDSO56zC
zjdrh/gYTYsWicq7Lo+JhhH7tFg1BjrB/UXntayS3eveanTP7ugR38s6x8jII5bu
z9lav5117F9vXYwHaKh7z8lIoCatRpsyS34qFRwaGHPXYXrAOuH5KDKRiv4vQmLB
ehZJYdo7QkEPKKYsVpNFy3na9CUVvRt5XmNOtQuqa6IYMn6EWkx5f5xzYsmgNjXw
Tzz5RMjo0MONOZaJfrCeCVCHmssHTETYRR84Wk8pzYqfrgK+kjFxHnW32IVAUEpX
AtTiRXUqsts8C1+7ySrsHNhuBIazntGrQkWJoere5PieyK86sVuI+fG5Ge21VF+H
RR/bqnm28xOfJEU0CGaKdnS4yDg1ikukSbjuPB2j5egXb4UNf5tRGCTbnW8Xb9+x
fr3l1avP8HOEX1AKeoPj/T+v4tRNjvD5+meWsVCfDaFYm8MgQe5imjTg4PRA+bmh
8Cjay34X1w6MpUvK3oinL2BbYK/UwixwQjguvmn+w/P2lblJrgiLRR3a/uQZfy6x
WprjQdQX+ZF0vCeyNOjIe+PYNUJSPjCrrpFdfWIKP7GVB5UxyNAedJS3ceGjGJAF
KNgppL4ikOYda7m8hxm7LH6J1cApdWlpexRuy5jXN2p4VqwaPmTx7rdHMYCFIspB
m6Ej1NVsFn/HCL8xTfPj0jT9Sa6bkY7GG+Y6qeTU3Obmd+w8h7w1liWy0FDn2k76
onOcJXxqS9ZP0G0ei6QNehFp8E4jGQ+Ik/4Gj3mOYd0IEaw9GE6hImWkxn/TPR5G
q4SMqWW/2ark36X9U67PFM3rHRknz/KMBSgIXvnXYJ4Z/sHTDZQ8VOeDjQEAgQLq
a+UwQeG0EUq4Np1SKgxzOFHsZ2nCCqNidi9goG26jc1S2wHl0U2HiJ5ei1PcECeT
zfBp7gsWLVvTXXcxAkNOeEn1lI5f1QTOJeDdH7hVBtPL3QSTvwPxLy69E7kZip7/
UYE6NWC+9x33fBKGMEfT+q3X1VaGD7FBqethZSPPF8XYpOuY44oWR7COzXA5Zsgn
eJZquhl4mVR73OowuIONaQz83zY3OAlHQEKXgpFl8le/vNkQWesTCSK4xNcE0/u6
Ch7l+plrH4xVM4e4oefjjKF/ezeo0GpeIc5ZdXKMDy2iBKPt7g5ksxTxUaclj5zX
oHrQk/rcqI5Q6WpJ1cszD3jjR87maBGKPMfl17zX5ZIS2GK2YdD7rCi1X4zKWaqJ
IWesKbpKb9ShZnsDF+G8H30Zb96dnaVkaWJ3wPnXB5LXwQWmuS7zQjMGAI7XDbSF
3T/0eP5yv8MYE8o8TXkIU1Zdx4R/sNFmzjtE0JuvOBeAnGPvGlS0Q0T5NjbT5iIk
7uZMWbdqYTZYstfV1nBWbbOWZttkhcymegpQ8yTo4LuNeL1xkKGgrWW0zX9r7Ohx
FaKMXKn8r8C/skw3tHGPmHPKY9AMzDowdQdhhkXYjlbgz4PVWqmof3KX8Oqy1Jo8
L9hDHuAqF+YpgcHaICxq8zfGltJRhiECOsh1g8EhK0kEVKUTXFYmVio8nhNyly/V
Rt9KvW40qO4ePOupAVsxQtFPX/DKJ5KkjWLn3UQuWw7sokT4F5aoCcpGnNMt+GMm
GEQcs4TAvsIq2lmqFXb3B78GeEKfROzc9rCLCkLEM9SI1lIaCBtmggOxmeWhgtRj
0j7R54vZTmK7vlprVUrv1hq+7U01aZGCz3mgw8fIBtFso9cJ3asxA/Izcl6kJXML
IH0H1SDvXCVIZEFpP2QrsBNJKPQkulVDN3oiryOhH1qxmnDBwdrwK4RBMHvpHu/R
f1t8onMdPxkbCXiWV1wueo1YGtorQU+Y9YN+0VqUqkQp7P4cfyoi1UBefmDe+KEj
KW1pdDrFWsmew7dGdWAW/6ZeYARNgWGT3spKCOmoPREHw6sb1u0rRHJzQzybrll9
4XfUcm9FIn9CLv+3E6DfbYnAKI2wbtXnqcVBtPKnZ+Z0TDsKUy59Zwza/9t5NTwC
rJc40KFEf5DDK8etaXqAakj/RI6iiuNF9niJsfkpcV62NkrTRDktONnQkzaIQJq+
CqpBp5VW88seR6eZfQ8zx1wQwn28K3Jup5WIrA3K1zowm1k/T5uIoBy4f8nwX1wo
p0FiTCl7nFXXBWOw4RJlyR97nhcpjTHyFpq0fAAbNE4XH6tT0VDWtL8c57E68a/M
QmOL0XgvMGb3/+vAEvGLW3Qb53MWiZmFrklPd4NcV2BeS+t8L577wyCsmfwlOGfn
nxMXJ420V11Tm5EYO91ZF3BzWaUPS61B9TPy9lCzIpm8ATMReLi4qTDv0AkAWuUs
DwxUKImjU5dl4gwv/QMNgDl0RmDkZIEZZdp2cH1g8Odz0Q+sFzl9psMhOkPJCOk4
vNJnBrnexMeBNWdtsjUeDBga8XzkFCyz1/Oqls3xsR3gVg6VkqlyC5XP7VSfKipE
jdgAOJHnLCCbwN6JtQEGEFItvm20Nzys7Fb6lqeR+nKgUA/l+0CcM3uuxLucc/0y
DS76xCA1chRCZtvP4srlmz5401OTVmWhIfNZZ22GsCVHh7Yk1LnV3uuHLvtWEqae
Z//3A5kfCafG6EDDU7kINmJv9LbOtBKbFiUqC2hZwU45XvCu9jS6ytd9mM/BBIk4
kSyLmS+xBPXjO/+E64ymXystVI7m3NoPD61XLuogOo9PKlY3zV/SfkVILqJ9wqby
rLTeNMO5sFIU+RlbJmXSXSowbxirQu+fE6//koEbpSZMFiA6FS+22w6QtsVbZk9I
BP4ct5A/3Q9aC8hs3iQHges8nxEUxX3TIKUkgmRdx7vTt2kzxZwp7iPntdFXMwZt
bQ5K2P1kaxlMdOnFWsWIClqRVZ0TigdTFZjmG/EC9XM+JALWFv7h2J2EKyYEcWIA
1LaC7dZALBe1r0f+9bVR1GXqnxsmUX50YhmHCUaBeEI+qkZw0kDdwuF1pR8f98wL
FtpJ/E+LS3zh88O+XQp2Of5ygsfllli9eB2EmV84ueJ1hGqzwQqkZezvGuL/uYkF
gxLfzs81BgBu0eKn2jmXHebA05xXcxhTNDyk146qgcxPwbQ6buqK4KFOWHrNIK/M
5nFW6SE8mYTdukcBSCLPwG+d9b6ErPa7/MLlV+Weh3/QYQABVPacCzVw+AjQtLoR
V8YXdOcn8IXPFPCppp4YbEfH2Hi6nKVoLMb9XyfmYd7diem38vLLnTpIu6xP9SN9
z+lgrcorqSXJ/OCNx9K3pJ7Y97l4IUiZjpBDKMQszC8f9pj57ckSRH/goeGX95OW
E5Tb3aFlFM/mqvHR5xOlY4MuVs0m9GyOnJTJB6EXDfi1YyaZ+RuIz/RtE1lwcaw4
F0Iu6zq/EWWDgMD8THn+SCClXNrOlQARa8u3WSzfGe/yGbIEhHTkxJQtRRNbxUXx
axsXZ8nAlS1x3RvCq3IOoCb9CCNEYGP4uV3a6pCPcaoZQ2u909MW4JxjFlbu05qB
9Xx6i/kE6B70Ov1DprMJb9v9FAc3z+YFHx0J4sRYX2KrDtvobtMdOA6Ij+znTqKo
SVNWIFTLXI8q+Hh/Td7WSUVVMyyCdfqHJXOHHjzTHgbzZW97LoFXz89dYF4kFhEz
uiZ/VvIlXT/GRasBnqm7VZuMR44KAadQIkZ+KQpkRIX0B+g/c9ldEtYGLI0zV/7T
pB5nu8f2FVkVgUJKjYK+YozAnyvLJwPeto5bjhS17McUIjB4/I9hGPmzb3wPRfDg
nmnHyGJ+JmnFl5XE12mGCEMuZPZp9thXzGsdEwJJZixKRbmv3mK5nUDQgSTj0bX5
DORgtQ1dkgpoeS+OZ3pe+D3d4kl15mheRQyHvb7lozsRqZYVVlJmYlhxmXXI5vhg
gbreU/FpUdG8+qOcBQDBxi+lHeAvcHeau9v19Cak8HiOyzsVdTXUSr+JaogogsrN
aLZ9f86hJKM4UeQUEMdmb7OCngHr+yDUu5MIowxh69ue7o3z/FXrXOExGCMS5nxG
56xhrRZUwpZEqbhYcYjPSKfaOG58kn0SO/ocK44nVDCINi7zyxBXpd5u8iBYfgpf
IrkGKaixP2G503pK5Gr3kqlV93krSswL75WM/Euz8tI0W+JeLiaoGJzq/HLGsJqi
t/db7E4dN1H3K2rpVLoBVT482J+UK+EUDbLa7ERAcgEorvUeXm5N5qatdORqSoyh
IkfHKNdSaTPnjnEA1m8BW4OhT+LoYflIkEdN40bawTeGKMMwdszTK74LOj4IhzKT
4LsMBtO0BnWQpF/1htAHNL4ARfm8H5wfv5EkEnky1BFqptGqS3ZtfhhO77PYiHcZ
rRW1S3KEFWDVaWfBQLt4cU8/KuyHV0w3TpGnynApiLSPKXa6PYdxP88wxYCSV7DP
wFLy2IABeACZRMSqshRAXQendxa1lIzJKmubbpe4VmuRT+ou/eMMIPMYmxli87T+
KQIs84KCs1eiUnGJwuC76ogkiSVAT/jc+gCpwLlj9QRYfBJC85QY5rmAIONkKym2
CTOpOqlsFfFdNrwCqisfCkRCOC759X6A62DYrTMbtqOqFcstFvOf6oVbtqf1vv8Z
UnzTcxuK2594wzbF0ruA0c8qVxvMs8CWSZWBw/Zh5Mo6nLNAxu6jUYniVrFD5cJ1
lafjNtRodZOh2emSIZA19g07tocTou9MbEN+v//BVTfy/L4YIq0x+eck+iX5h/Di
V2MqO9g0CQyrhwkgdS4XczrnYPM3UkbtaHbUUXGcO4dXAt6AbCrg7pPNsCvtHt5G
huB/j5i8qN8XgodSUD77jnwxxBAspqzutWAlBp5IwBPEYAttwcOcgFKa8CKK2ir2
YSy0AS4thZe+TiUwUPNo22P7bcLeybPV1NiV2Kt10WxlO0J7lfgMU19nOxCjxNBT
zKcMMSLMoOfdlLg21MM/6bsfBVAG6tj0IV1hxsJcIrwbm1mPG5B5SGEsU7YUy4oN
AO5Z0IvEDTErys8bc7ynYB7hgw9eRfTZQT2Tkt/K2Lr7IP6sDe8jBOHFFBiGMEtf
I0zZKDI1U36DbKKHcp29+2DHmRO+2H7gaq9KV7F/4RxvVPoLrzJ8ji5N00NHqP+J
yJEZJwzkIRDnzW4SK6gXnpyllEWIYkxRAxqwFJ+oKXxrwiwQMvYEzI0LDOObe5nz
of/ov0O2yiQJjEOb5yiBGbuuQxqWPJwgmJCNqer0AHn+fOulAOOTHiQSZTv+uJUj
F+Eip2h1mvrGDoLuNFKZCJI/LgFwZUwWGhq5qMmn9IxPQizllP2mG6p7s8WxGFvG
zHqyFMQ3urUQnF+NwdiLluvN7KJKHdGMUy2E8lGjuSISmfPiKb16kt63gRyfDvqX
h/WQ4v+SdgYfdMsgfPocvvPb0bkhky1KInhd0xDHsD1lqBY7lmoOT3v9FGo7fJdL
NWucwEuwhlC9EK5Sk2iAAeoL2eFFfmTYGuIjjmOwwMl643xOmwfK1YIZXGizpDfM
lsz8jFjPiQH6iMNdsRaG11dVKrACm9Yuh+1GoipRrQAByg1IuWps4W5lnDjOPHAy
V5JOgp6PgoZN/vphVjlVFJ7DhWllsqVZDSkVKhgLK4WFXpWN1xfTtsw0JqXj+IuQ
M/KEVM9ttZBWEMQEVWXQnmgXfg8uUi0UfzJICDsqxmxAAXPKbhFQsRw2gul28/rJ
rn8VIOTjOYnGnhSZKF0LoGKJSsNJr+6f5nu1bqq/XOtNfbSut5xeUb/S3DygKZ9T
YYXONwDL68J9tR8Rug7ixRFup2rW9D7CacQEXuBme1/Ku26g9De5fZSKy48ZEjDp
D4JEfpyfVHXLzxV4h3OPRkWC2K4OrDUABSacWhlnhPdQrJXKeEp7op9PC8kmqTEs
WuWnRtgnHWPup1P3ZBq5fnHbOTnNMiFE8b3/HVeaB9Egiy7gRIyPfx2lgwq4xwE2
ZJjU6qiD2ca6b6AEoJviUMdkd4d8RNJL9wCo3VbXCX80wKZzJbv2tdkFXdtJjQIE
ulGppgM1HTW9YIWOAsiWq/QO8JxAB//lO6p1bqJh955F1V44Mmd11mjWDvDoFvv/
qVfShm/tD6u328gI3k53hbQgIwYywlVZ0B3IZgASngUilTL34/AKGTI3fuQfVHp2
ntomf2cr64CQBDKvaWxkUG/0WMoqncFPkjUeso6fFkBm7SNRMsa+vio9wORo9U2P
u6mbp3iOk9/wtxVdv059W922st8+xFCEobOia86dERTcYdU0gFPkgYrLoNyRgTAs
tI4LftTq/2slSihzjMY6rC1K+VahxAxCGehm0Fg6SXMrZcaSx/zynQNN1QmhVeOV
LivqNRJ0qUaIBikrtHFp/aM4FlYP1CZcQwqfi1OGjtoSNw7JrSEUnJe2FytigbQV
+HEymfc6IlbrXd91bA8ntFcQ0VKn8qKAQBOyRvhwKo9TXoRVwHtkf17x1mLp5uSr
lQEx2lrwq7Q+wrH2XY3RlvcviO1sxg1tih1yH6xWm1d4lZlozowBU7CpgoKaFL5M
Wn3MrrrAfYHSdMLt+mQ44ab8CudpUHBJ4f7bniviJIza0wavyZOSYS7FjDWJoOoj
PDwLCeLIL+HwlRzA4gTIgosgJqVw9Bu3SsA1PCczK2sZBLw/2XC3UQ//upIgT89D
F5q6xVd3SRiqRV6AJEuazDrkiMN3H9L6BGzcg3zIc0GfgvblRih9a5f45i2ItYxX
Yd59TF7g5wecyfBVtjksA5XKrvHnnHCAT9BmR2WxR4yJRW4gVY/mEEWIqolYVBvu
D72Lf91YYNGitLsIzOQ5cS+6ZpNr9jp74xmFcLY4A4+Q/TRDdLzbf+plOBr86+M7
YVeAMiEBgZTG96JPIeWn7uQuP/7StAwA7AyiLIT0WK+RTg18nc3LCMiQ0TGOf/a3
oMHu3sDi0Vi8ixSy7OwXVPBUwqStdWbAgTVYb21utBvrvJZynwJXXsexwaRaADbB
vtzEpTkqaPL8ZbUMTZtGqOq3dqpDVNb9WVj2GKaN3jH7BiEop7082+QibgsWJiDY
zo9VlUaWIf3rLBdbMu246HITYgYotrnBPNiQFJtkzmLM9pMNXlnXI/vaxalJ+GYM
fVwAWeq3EDqkD8pN6QcmRSaYLfAs8c7TgtxIC4LHjbGPIAdMZuxSluADhHinkdmp
F8kZOKsSOK7OJdBCccb1xsELidd2Da+N2PwQPP1ZsV79EjcuQg6xpdve4oH3FU/m
vlZs1XsUNsDz9o0ennWkpTEySKecdHeX9JQZLmA2k3lVwp/FmYBHLJwKizczdkH6
KbBFgurX+6LxKUOx1DrwKRTSeKeuiTYrNbeAH7MPoEulKaRg29m/tHoPhxpXtfnz
e6hfUi8kf+xApXYKBkoqEyzcLUmkxbA/le4Y9QDVlUUk0xCYqdwaz87u65HczNDs
okN3ZqeuC7s73A0YE7DnijPFWshAF+TVqrWZ3r1CjuNhBGETz4CbYWXVSu1a6Ma9
oDEtgP8mTpY27I56gST1yJU3/3XoRLzR36q2L6sh+/ZWPzq+zEyrpkZZqfoDrpAX
KLf8kp+DS8WBDbUfDBQI7SRh8GRrHcC/FR4cGUNg/TdGWpLtXS5lQc/8tiKZnBAa
GdbU592qz3zHD1RXDHWK0xoDnbLub4QTL8vrLxlH7ZiZQ5x6ytTzQUGdqeiFiks8
fjlDaYCPdwD49tNzqxHI6LGtqfdrbzF3hwtUAkdDZcmrQtVsz0GIjEUUspRjLqx0
0Hnck1vJnbJHVNwzR4d+T4F7TIAC+P1gbnvRplnCeE0+UxXmP/MsYhSrGme/2T3b
DUtIGGdX5X6aoF+zq4LtcJmFvoM79CqWSu9o7aRoNyPB+SCqFL2JnzCWem9MEDsq
zAdvPKhJPD1BW4UpgiCvdueSwb3wia0w78zH4lucE5YvP4ZNwnGLWmsFyqzMbO8p
wNMs35Loz2FaXJR+A8MD3KJjHIEw4UDNQjvcGBR/8JxDh1kKMmQpqySRvYj5WAU2
Sk1AzmmJhL7Jr/pZqfIFEKwzDUiY4rmwzt86lpBT5OE3gsjcgKuEtCubVkWOKoO/
FPxpJ3ERn83/1OEYOTm3vA605tVWt0vnCI2nwJPG924M2kYH1nHmppYmh11YCcFS
Wr5eGwq9UEyCURxn9ofM5N5rq1bYG1j/ZM9I/spZHSV1mkSLRWtTmv37Hx7zyt9R
BcuPcczU/cSgFD2qsngHc1Ds3MH0/qThAhEnv790pjv9Dwoy4zTElf5ir36Q++3J
axxUChHMEwEPF/I3mkEnAnLC4BAwWdwMMswNc7xbpcBl7oSLs6uoSpFj6AgQ3hPo
pbQWNnEr8GMOtEMrpqRnxkdSCuC63X6dz1GSdW0GehIsex51LCufvzQzQty0xm3S
v0IvKSU1CqV731Fo6Rw4n4ai1B6l0uFY8DU120EAxajczg+IBcDJrGLLLdXui83Z
pIvnNYqoyiZusjQQ7jUsBIVKIUe8vOW9GPyO/qYRBYv8a4YprxI6cv86RJK1olrW
XfQx8KBgcKkUbRQiEYMA4/y8XiL/4SrUGMSP/k+mpv1dDOk5wvPrtkb0cg1k37Tx
MSSJ5Kl07Is/HW1i42yS19Ly6oPNesntomzfvWgYl/3nFqFXOXd0Ka9TKxYuEyGa
lxUxaW0i2Gc9TCDQ8GH2FwNMX9pMtWnM8XVAX+W0sERSwGo8YFCDOFBwaXEo/q+Z
WIIikJECdlNi1hoDwXhEBVgV1WANq+FTYkm1yAblaJMuUs9o/9fl3mb5pnUHttQ/
v3R0ZShBm0wZVlnig6Uoo4CSj+a79COk+LMWu6abtQtVSPlDTvaa2L+Tku2wHzeY
Hl49Ta0Tx3uhm2lkt9M6O7oN+/S2Sf250dLAMbnt2wREPFLw5WvhHe19MqCHF0q8
GkDWysqoEjj5ECrVbTPuuqqsRsazUyC/rl38m98T3Y+cmZ3KmmA/oAbAbtM24OqU
4LMsaGZp+qfITYRmGg97ktKY/OAdt8xeT+Ey7mvkR1PfxZY6QR9ix5LRCS4YouVd
aZl4qtz/1t2xAE0f282crFdf9SMxe42i5B1jhH2Yv4H3XzKFkv3/53zIW0ehCpdI
sC6VaUKr1CHQRNunPSxh5Q8sNDoD6f9vT8erKm5h8OcCpXIK8amdxvph640MbnqH
S0FVvf7Qm+a3M0NHkjl+VlR94ipgRL1Iq902V/q9fLanIbqFmDkCPUIQs9IiqOqX
ycl0/vYMzwjQId2OJn0gjsZQZ2Wezs9Y49Gtmp9gtsoajblDhF+ma6TSnvGw+Axo
hhPzTQ1oclo/cYc24SX4v4SGviNZe0+WCFupecE54moBIoTi8xlxxQvD6PioToKP
fGldMxsRjh5t8Y5acr/eyftyWOqhK6LwoXTOn6QYl2h196GTkVP31PxDIs/E787X
DIPJrk4kxLWPcJvrfnlK1dMu27jwXrYL5aAOSFGdlE754jzBNc0hOAVKu1sKEMnr
fjwIJ5ln0cdUS+t1tCwmEHHOF6DaKV8fXFlXVfcLJ8LPu8N7G3lHJe4//ivhOoQ7
JuEbZwKEOlBe1v6loDdxAJLGKxzRstLmeiRecrNMCtQnG1YsvqOnJzOujA24mPws
cS6t9BmdL3TbpJTU9LB23w7eph0eVDRPMBhOm07iE1W+afLkTSEwrl42dz6VR5pk
ov31orjMdnUgVoXvBAZsLcAUm7aMYiBeq7zKh8VA9bY6RCHQ7NgH6qD+ZXYtaowS
qO7O/HSI8e5ILzjc4hP5mGHzSxHKnRepaYlWGi2Gc0roO2gXZWhwuZWUqw7H61Ff
pSGjGL5jCMcCZAE6SxOLRmTWq2iNGucKhSm+cZxvGwBTak/Tk/eV/GvHTU1X4F8v
ld5IqsQmoc1e7smKCxsTXCOaZTUz67aF+k18R8zj9YbCs09oybAo6nvSXTKz9Y4M
Wr1PkZKFEgZCY4ENum5jhuRVKFo3WWc8JPWMEbXJFhGdk8hG5dSeOxH2RSmxKgOM
BawdiMvp2LrcuExf7RSO61T8mhku8m6dybsstvilZnskUhV7mwVD0rOD6CJeT/IM
RG5DX2LcJv2oGF2LIiW21GjUz+bIi/0Jx3r/ed/py2yhBeKwmqHCWrNnbaY18Cb2
YTlnjKMYUeDyTb2LrTF9r+4ocAIhrf4vFnoV/yWNYuwwkIZ5EXjR4nVxutvVIjfh
OtFOawd5/ZOUiCSIW9zKT93n9cOBwE/FZIxKnHNR1z91ohfQuOFxKwgev7xNJlE1
LxCPxu59wKuvTxSxcbEpzqu0vL5ksfp+67ZV/ADEJKAhDKcVPxVMIU3LyBctbIfL
mRAGgS1f8XDPOSIugo0b91sgqqIYa32brN9QVhMgHt3WMsfG4Ov3/V4HprspH8IP
Q0NpOzBLJavYR3RD9jvxwzwXxNQgwDdPqdLMQ28X7EHaqxqt58SW1cpAWmHUQXLH
dYRUoxjrrJVKojfoRm7PeHyAS6RLNUiMKsheNEg36CpbKF/LwdCUjM0mQD7+KVHc
fXm0TzYpAG71vKzFUqNVf5aI3orA3L0025u65EReOz8Nczu2+t7eBLFzZ9+/Stzh
e+f7immFCv+lsOC3hVTSdHIrzk50nyj9hS9+F6yNWiYAc9c+p3H61MnZhSaUZRib
pZzN2FECtDQoGFyv4PFIzcFTpQ1xcTOz7p7rgpQ0GSU5DGqa8pAkZZjW/yO7p+Zm
MoNjbVAUWXwT0ySYPH+8oASEI9M6IHldQlh4yU/ipJ0zJGCHXpcApwzFQV2vgcQR
JFi65puj4t/YLZNDmlH6xclvGEJxYEy44uZUOlCMmRk81XLU5ZaqIREgl6xMKx0/
vGGaeY8BDzDKs5ffRnuhq99oQpCmTdKjFlJ7MMPZPvJjdliVj36aipBMGjUdpaFw
ElF2O4BHuBWx33s+Vqd5hgQ/sljQK1iKr7lsh77xk6gBtdH9uRMkzS8bm/xG9Gxz
jXfUWB1Kf+4StX7Gvs+yWB9squF5Jemur2a7WmPL+QbCFyTL4+L5GUxL6XlqNnIX
cNOROrd8qa4Kt+CM3XVxSAMBk/0YrHHuVevzFF+WnKBQJaKmf8WnZENqhvn9fHBH
oZRW31x2cK5uoC+EPPqkuEWTeqSYyaBjEXUqCWgNH7A1pYKJAhiJpXb/ucfaWnh3
PPhZGSiT7zAwTip01yO323FYhfL7cJjRmXob9I0H0fBxSoiDFjCEU7cbtwx8857H
z+Da0iKcYkbvHgTnSqvcT7kMc9Oj0VjA6GSPuOFMeO6F3C114eunqLnHAHYdNiB4
BQxuvGsvL/tLXHZTmf2E8ziThMD0V1GMH3N2ttUBSrs7wfCxAEdwLKk+VG12eY2U
O/ddfm6yLLsyUcZf7dOSPQ3zcpb/TCaLtOvkYjwlXTo/LoXnnmMVgWZnUhTk2zV0
Z0Jwrti31Nl8ktG4I27uDKFA1TNcvhT+bUd0tBMJ0iD3WOyzWVIdevYqYCxuNLKx
b7SSEK+Qpv42DPevNf6/EY9iX5RHXhSEPAFAvQaslUyuDoRQ3w7/cfYRyQdr+OfO
UHjMkQeSnxEAtm9eNaaO/61RaFNEPxtm0K6Vz74R6GNQvhEogmnMx4ytELoxbESW
BsodZ+ND9hDKX3lQTKZeXnmpivvN34TiwhxK0nAexWVeqVwsicApT4X22xnf/3dT
qiAldGQSAqiK9S1tLzQFQB7tccP/2X4y7cIWDhv14I1GO+/5rmPhWlMNC5SLD6qu
gqX8UgnuAL0y22xpweOEHQqdk6O9EGNWN3CITy7LAX8AHV7J/u0333TWXg/Jv7cs
+DT1XThMyvCOlX0USCDzj2x5WGwfWyZ6IYrxZF+pY3q1BlCcBYSd3w98yMCirP9s
bgMa3pzaAXuV1Lia/wHtIjk1g1oaXsH1pFPxbeOmFhE4Ce6u+2jmsBJVGYAkiOio
Pko8s/NOIYpjS/T9ckAqaw+z8Xttq71aj70B1YoymlEEGBwcVZXZZ5A8OOfaq8XI
rOVL4je0cqDfuZ4o7Gh+DjqcBHetbryFsEgPG/NsE7KkO3n4fAfL501zksXAtMCS
pwq3QNxxNoi1IqAA0SrISrLIzJH3COldCMWdeuhGtCQ4x4JtOZqoq9+KFpuXe2IL
uowA9+TaeX4bxYTsuFPZb4MUMrEFL+OyWEscKs9Rg6qvqIyKc8G7//YVMpuXB2Zn
520pmH1CoseL+QoSdQsQs1r6AkpcOnYE+ro3nol98IBRgqZqyVSYXGuescWboqvN
ep5xie0+RAO9fiJjfVHV6Jvajk0fBy+BW6AXfInXoUSO7zE2eM4ASkR1P9j0G/KT
D1LJ/BKweZ6IEV3OlAXCxIXEmq5jmmgPlxtMwsnliQWCcazP2SnlIDHXUoH+tFgd
J9VQPuole08UJArOh2LYHviYiYkDDYd0iG4+UZeSFaac7RIYtaJuxLoa3zLcicC6
T2qY8aDtrl17AiTT3FyAKV5hzP+eDxNFjzuTvI5RL3/Hvaa/lDMsxTH9wg3OuPBi
mShgUtuk5uN1L3G7Qd13YhQbwFnE6cqlbvmUv9j3wjf80BMf6tB0TNDKtHYctLDy
7e7xU7iPM7qlMXJ5DgFELjDuGoP8YGYq7BagGF/DVRseFYMLIvnQdCgDjXK1Rqq4
NnRB8es/3UlTYTcDU1usmKR0m34HBp5xi9S24vr4qp4cMJONVf5XPcZ4kzzfFM+4
0nBROZLw3yO0DfpClonbpxxrX5r5Cr7O63O87ZZx3rfFudwQLOmTSJJU6vsMWA10
m5P2HbavPr761NEfgjrjd8gwi8QWaKW3mbQ/FbevrvZlF41pDNUTp1Q+Fv+2JKIv
+OQTsMVMzCCMFjfeWbUFbqSy7TQdryN2UZBmliXQjpBcRhpLKyfdxtpIMntbljFo
uioSRQN3UBxvAQrR6nsn4U3B4iAJKaDEPGqs693REt9qIf3oraHJDGRmP2XEWVcY
IEI3avynml9Vk39Uql79x6PeHWrQgG7iqDvPsAFGECzRW4Q7GXrPvXp3RF0A+0dd
v844LUPKT6/2kLgXa4zY81xiZlKva6HmwA53KqWHSHTtl+Yn2QN7mGg3CoQHqZK2
S9m6ACKq3DLfN+latjFcQ5DviMAm3Nsv7zGiAMKqr4lb+UI8LM8gRB0zX6GuMJwS
IEg2fxq1zm8pT5MUSsjbQC2jZHSOASbaVWQt2Xdzd4P9YTXfE6w1dyBIXhOLXKya
u/WgaU/477R6xGBC0HwjDQfbyNNhm5EJjmzWd32h1tkKsENx1VP/pks/4zkEw4C8
tP1UUL1EJmeEm+08PP5ii4TU/m3VkMV1LFKJU5CpKsLgR8PdjYO1hWlm1T2OCGIA
8Cv0jNAyh7pfbNyRaTUUawvXprInjjpLxjR65lZV2sq9SHz6ouDBDEU0kIoRdeVH
/fC1uXJfxyLxnFC1DF+3lotYn46HPtRQ2bASoa58yiIgm40Q1FI+7WeIpoFVisXi
SRsT93H2LoscpI73V7l2MI+pX/xYABhwnWlACG/LiUzvFCDAo717wHBaBVxwLUlX
nC0kIivXlC4v4q9+d7hF3ttxascxUZ0tdaTUs87tH3nMeZrZMNc7KgQHlI3mE+yy
3jbu47Fe7YrAj1yK1VDuAe8L87eJvfLSpd6kApwkCv8fq3tXY8j2ecBcyif9W51W
oGzKwF9/6s81JSnyETltEeqmDG1+bH9L+9Y7iLeShqDE7Qvej5ya32y3ivr6nJAZ
jm8/o6JnxqVgEMDz5XdXdlvTiHJft3hMcNZANDInlgxz8A6NiavrbAOHZmTpOfH9
Kipc7KyKjYllf7Em3xT/heKWRriJmCZRqAMk8jDTDfNn37Oi8IOisdjpcpNyZ1L/
opcixpBhmg3uM/uQr+khw441a/v79btrDixTrG9d+tvYrQVd21HCp7AG1NR7rfSS
nyPG71NbP87Ztn0C6lDL5Z/9WjHHfD6gqNn5q8J5x3psYpA6ZMJJUyZHbpT3fn2y
JKvU9jqUYHz34J0dI1pyUzXQZE0+83AE75T2rYlKxZbBsvPbqlJSVeX5L/qbqPAS
oxYa60snWZRJlNyE5fsURN//CjzRtqZfZZ83Iot9/ZneUkpv5AXubAxV9+VL5LFH
FwebfWckyLS9UQeU+zlpGWnqdcY9dX9538FiwSgf3fVB+PDSQSY116q+L0ladFvb
bP1vVfugMQqKd7hrvwImcuyz+m11uYNku9gW8q3AqVZEk55sRx0ojMvkbYwYwJtS
5Fxik4a9uMVwiD6WIPhK+TOK8WNLxTEjx25LaJSvySokiddYddJQJ8eVab9if3b1
iP2yOXv35kKGPOBR5yayJEYBu4uiU0i8ngb013Ok7xNV69LYkpK2WHvboTRTet4P
/pDCv8fxSAxNc5TBaQkvdVU08j8oDPMrIfpk30LOUcBWmEjXjZ1w+bmhlUZZ4hNA
SQlez7Kq6wLfR1KNvOwkT9q1xpRx2nIyd0BDMVCPV2j217pWzWZmxmSeEUh0jDyw
abFragMGaBdluI1W50HM0uNC3AYePqRT80vST2YXV1FxeEbl3BDPnga3KI7Y0svk
asnndBAuAi/LD7vNxadiKLnXfUix3NL5RBbgRt3tPaqDpN3VBy2m06BgezfZ2MPJ
z2AivZFbjshXNQJU16oAqbOlqFFCmyg3JINpTTbtlsYUkgJalPD1kT0qTaootjt+
d4xBxnzLc9HIMueThUENtGCnk9tHTJlkTDhWgljaYKkTQQBAos9LGtXFjUVDcw+n
hJCq6GX0dEdBbiR0yqSzYMJDvNGoQ4ufpfXjvegJdXIsY/evlSGhQUcBJRiVVD2Q
x4P0K4zyE8aJa/qdndpSJuTyb0DTkAuwOcVIYYURwAVoUvU7NQv/Qg7KO+YGYVoB
AvQeH8kquNaCmsNikg6X+U2weVu3kK0oKhmsO95LPj7B/boMtADrH8czZjH4epLR
Rh5y26IOJak5vkLM54shvbXlJ7cyzJZhbCkAG8826iL3OuZMvMiRozGiNWnpv3SA
DbwgZ/GFBvqovZc8r2CYIc12Y749Bz7dSAYGXF8xdJnKobZw6jUg3HX7hu9px5rO
nFcBSUOPh3lUyh8FNP84TPS/eLisfHnY6XhVKACwOaemcBoUd/SeTqmtt86B+uHa
vSFjFD0z/havebpmQ3P7tuxHiDo0cGaDvLx8wk048krDkGSTJo/fRMgxbmkrI3cU
0+nUgIN0eLDE5Bi4Ch4NlPyFmI8U49bV+25dVWqr4UjImeb70YynaFk8HHtExN/l
08P4nprp4Wxh7U8hQ3F2MlUHXYKUVugchGMVP/LiBZ8HLzLdLs2I3wPZdXZ+V72P
XlumzCCXGiPKUEl2QTSwlb4DmhPGYPg8iempEoESowlKw37WRtKOn8zfyydlKCC/
1oRcO4bDlaEHG1TyRGzei1mI97dw1jm17FSm8+5d3HsPUxowly7zJDcfjfWmCbG6
Oryb1xeGG/bVLmhxtvHQPP87Sk7GbdU0gaENhByXy/6ogqZQqzWhDs44o+U3LyIW
2HPtvJXO4S7/z3Az89oVNIGKcuZgcyKg1gI0m3h0lSQWJOdaJRTyixvPgsyGPXo0
wt8ZOksHbFrbgtPo8WAPuakD+ebkSNvFMdF0MWuzAUFuAq6fbOwVqPOWKIZfNVzx
zv+8cbGNJFRC6hGF/BdXZ1JCyIJrQrXUfRsuk1tqkxb5FcM2dloLStLG3YC2YCln
x1D/u+GJi9imteWJUqkKw/l/sh/8y7UEwl1vsrfJge2n27Xn7uzuHT3TUHGNRnMy
d7zScS4+u3tN1AovHqO6Bc7plBEjPCuGHfv4/2W26K+HtM+j6t0HV8Uns40cs5Jp
ZsVCK11Hnc/4RT3RS3fS62YDxFEJ47i4aH7L8sxk463hpveOU3ZGU6VDPeh7zHh+
lMyYqG4fDBFVItblZKUleX+JNXYF5pQSo6kFk9+AGcEPlxWYIHVAykRyV03Kq+Hw
hjLcQk+EnFt1G74+ShzkprGPrpu5fhx5s3yTOw94O4/l5GU87DwVWYl2stDFaUnL
AQuRvpAoL8V0hZEDLXO9r762IKu6MpHoAURrql3F1EXOTrmtopWl4Sl/s5dWnsCO
joIrHZkiDuRsh2KamHQ1OS8wCaOe8TI3OT1t30ZUEY42CfOvSO4HWZ3e5vSHzuyY
1+tBawihWp4Fhe2K/0ZAt802PhVIaGyMOlAgdZwPwkqIJe6QdtuBQ/z9ccsNDa7H
xTAnmaDPLcoCqYj1JpFGxZT8UDWuRTskiBcgIiiWIz6zKyhyX60+KnDgKfwtn37C
7xisJMF5wqjQSsSIf+eO+/pRdflJCVWcBNEclXg2OX1MOLv0T4Pv6Wvq3QqSjvE5
bRssGCNE+h6VH2w3vgr/KFlpr69E8dEtS0La/ISeRszzB7/+2lRIyG72CkRqxaZd
P9v/4yoa4CFRhLIhbV4iEkvhnz2mdz9R6gbSTTrm1WtdnViuHv4PO8D3bkMIgJHJ
HZGLQ6o1bFBGZLtfZKeh+3r9lXAP2T/tMODA4UF9F0NKgDriude+GV3wIzAX3DTK
WgYeZIXR7QiLK9K4TkmE37g724OfR64nJ/ffBIWDxKC0Xztqd01mxSU9JNzB0kXp
1SDsmG4QCXkMhI61Jdwrq5VhGCixhXrzQsF6e6LoZfsPILF8OKPvAJAmG2XDGVAR
vwS5Dj/YWTDU7T+58VbU1C7Mp2/PThB0O6/CG/IdQO0UKp1mGeVFgc4OK/4vkOiB
U8TFX9LSrVch6VZE9PxZ5JP4p71oRm1q4PbUCa3hLM3hTQR2fb9tfY1vCgdbo6Jg
4q5TB4PCpRU0gWsRNWgkZ0xXl3cWBX90ozGNqVeks+wLvonH6aNXiGnu3EAxCakg
WpbeDAn8x5FYdtXGtHamFogL6EYQnynKetg9+nyJRrQm31gIYTfLHX8lN8r0kLF1
cGreszqWCzH0feUG+cA6+RSIM4QWfvTBewQWSU3gi5H7itRg+PEQQbl1ptf0FajK
kgGUzP4CxmWoz3OCvKRwGv9P8Ux0v2OJ0Voess3u7WOCBaa6F08dBrCh5uLjGgU3
0Ln7yjop8TQAQxXcOYNevpWSQii99lbedw/Lrb3Vj2zkuzyvvUVxhgU0n1k46uqa
8cwb1+1NHS5qLmdUogJqWIOKNvtKPiqK4D/eTY4hRj8cw28bMThDiIk8vcM/gHw8
mYWkSer+M0cufRxRCQjkkgsEz7fpccbIGeeNQdnzqY7VVHC3F2hMn28Re9ZeG6ZD
iviTiGGXu6gJh16pjt9CPG0IUXfLVHMbwUdUPH/qhb+0KUDtX8FnLePtaGUgvNdu
W7/3j+mBVA2j3qe0k//4QnRJJdzc3EeyjQWBQjgpd1cQhwTkJE9MhZxQH/sZ6KSy
eQc4SFVZvdYh2WqBuAAxbfIHgGRv8e20/GJV6vnwWperpmWRdoNCzIS0X7u0/gdi
fqsR/6YSn9vahVwXJVkrtKyrMTp3IiocGUd2xIS47HS9QyLrX822231kfT/FDeoN
iSRoX8US3ZOxFZ3jUp9KRRjp/ZLH15swpc+EzuTcJDlmvJec9C43I+2Jjdl/oAFx
lnNRkBADlnLuWtqlLvWTU9ZJmiSH6J/q3FNxqCf23gKzRvN+RkaB85LCNwhyLo62
fw/wAR7JiubMNht/1xOkhpNADwjO7aBeQKH7/XAa+Med10B71MjLCDg8kBWGC9i/
k4eQuvNNYsa79LE6hQYVi4dUWmfQEM7WTYl/eENLF6zS5iHI7YHbAdezy0Dr+pt8
6UowOnNZJHlS9oiYLKypEUKKWqlXZbnbw9IH3Nlg6n/PLpRkPCFvvxdqi2IzphEp
iOCmVXW6AKKHnv7fxsCZNxbCPXd1/cys/xY/v53btxmGeU7l6ZaWTfFdldbiuulO
nQiDKCcfhkf5Txdwfx9Cls+JkgjIKjDEZ72yWFNNmeyM2Q+moJPmf84tV/nAtoZ4
esFetH/iR5ZxVStUrfAGTrfUfxYCgFi5Ni7Zz1T6TRLkGy/dwNNNzlj88luMKWAA
Hcba5SyQqo/KIBzfAOK0g/83w5YDihWwD4f7EqOiuLdyQNRuHLX/BJwOw4xqpK+q
v9UgfI0otIFJmdghIPxI/Yj12AJ2autC40+bepYcRSZfAeIPx9ysUWD2TO2lgfrz
J+xoOI8Be/zbnruF4qFpfezLJqWN3qHTk/sa6YSwAxC1mJWO3lndOJoA+K9APlrw
kQLsmsFX+CAPqNdXOios0EKK1SAdDn88fk7IcFHs8US059pmGlcH9tkd0xtgWMB/
IbCzO8s2z5rpWX1wdlPEHGxln6It0BU80QpHhbye1EKUj6WGgMoZOV7SCgoHmRAP
Wqq8ZiRDiwSl9cG19FpvWQoYa+bI8n7Ie3/7o1hl4I0RHoSM0rFxtxAmy7QLOe+g
9Qb4ahax5wwfHMLJyn2uIcPXvWuG05AGk/7yHQeVnFHldgDNY+hmcC8QDgkZvqdH
cv3famuB1pJrVnLs4nb6+VPXaGvJmFDA5mu0Hr9Ip7B6NfNmUvP03m6aoQumWaDY
qMB8KT0n8qJqAPdUCSUCZx1ezJyV21tVOBsDiSyaFrAPpaCtwuELYQc9A9faiCTR
xAGEReVv5buNltYPz9tudCi7B2NSsQdIZI8Na0BFnU1rPDF8H33TQqoGMDXNXiVr
EWBqcpIDvr/bhJMV2TtmRsNeEIp06U7MULDKpaeH4R/8ub95OWZdBJr0dC0MGb3v
KptiCeFwjEcxL9N5USO+Qfkfe32uAZwRvs6k+OYXDAyVp4z/9U0a4XaIZbi1L9aS
LweRFWKQU4rWFNA7RQbmmt9+YQA/ILhDP/2IXgID0Y2Sl5cAuTgMeECX9/YB+yYp
j0/645iPovSjsWwpR0gYO9S5xwbd/kZaSpUUQbNVoCm+mEc295w9i/evVTG0BMcW
9tk2XlKFCx7VS3YdKLXg3+Hna2vy+0cQkul+cXO3yuFyFpNVtzgPCtrseeJOBEg/
tQ7kN2sELgdXpxnZHx5BWbOcp5uCCCB1JA/SpOgE1ntS0VDEKw7D1slvLgJauoAV
GtSZZS2QGtILFXwJ3Ghtq3OeFPC+hXKMtHKARmJEbv5t01XCBY5U/VX5rzmk76Fo
z1tb8wJWQhEKE7Pn2/7f6Zt5GCAqz7nc3uhvLsWK3RpkGR4V49U734JOf1ABcoHd
kOVf49eIrbT5jTA0by55WzpkFg5PVJSBbghZrFif4Ey6Kva9UCcXradL9jkgoZmv
sprEoh8Lk57lqIWbigR1zyvFQMBxkSkC3KLmZs7rLKJYcp1Y1iX8Xkp84KnRiwGN
Gazo8D+/q2ge03CNRFb+QV+pBUqU25g+EQ+qnyPcJ9F3BMgIOpf/8KdBbmnZsqRX
CpvEpKbzyYMRTsHimGQecrv4wtE3CzmFedoumZvfFWEmo41N/5Fu5xGiq85LXBY5
riChF7xBl92SBu9pBzGmnV2thJCkf6MAezfKqwEprPIUw0lw8yeWV9zvadVZp3uV
iw78DZEA3qhvvosYw+fvpUZXSSm5Q9F6V5dJgQEns8pW2/UxKLgXEuAfJd1Fuj3y
MdpaW4PmjWmzg9tKpILjpu+94g9d5sl0+L7iJrDOuY1vWH4KmeY1JN3nDUh1RIvT
iB0c2inx6QmFNGg11Z9Y7OT8Kv3EAeFBQBeoEsmUsaLaQlM5TDKqdtkOc9k6tqwH
ZT+keWbnL4bv9BnEk4dcpgx2fzhakXN8iOw1zVk8T+NlI5neCzyDqYB/nDwPa9by
fQBVMh/x3G6k0g15E3dkvUooRzTwuhh2LlXsAzFW8XSFkCtLTUZCFrXlxlDUG5TZ
sBzyFCHHyRd/C0oakuRLLmpwnzsjK3sTZV/b0F1sUvWzy6VTMbp/4Y3Jl6gLwmDc
LDFyGhqPPd1mvd/xw8Vx+k3/0OOfUKURHf+V2y0Il/jhNnHECsbS8hAmnSTz5NQc
dCrHEO6vDo3LPCb3itXn4octZycCBLvUpR1XMUIKK0t1O/x5Dk8IBYZ/5beAtQSl
zC9adYyM9VZ//UH+FriH2mFjWpMuI6ve4/1M4RKKjHCarxXyrN+UVuW42Ild4xnL
B7ksh7ufKQZ+pPpD0POZSyr0lH5HceBGY+gE2Mk6BaQ96P6givyDB0CW0+pruFEX
fVrFTXaXi09wSRE+7HVQ/HdAQem6RT71H5uiDbQY48qE5DknJTuyBmT0sCZq0Dho
N1ZfTn+itkHbRnn6HbTwIV474bM512lh4f5KYi8aOcowkivBEsAWHohNjb60WYge
dPLk27lhrG41gfBbg+pDkGoiruC+LJPddP0kS+4Oa0TTdRUF3kh/8vkSD6C4nYpM
vpgQpL/keh2H0zB7SGiLTgWKKBw2mFQsHxFFbkjyXOoy+yHCQ6fYVWGkYzD74Nxc
JcoScfB0Amfp7BGN3V3KItEdyhpMoOPOCejFryymKV+v0AGerkeEHdWQ/NkFDSD/
p9RYt17sgR0Ib3LgPP0KMVQ4Nwj+IrSEmXkldvpVgCuImrTn7/6BHgh9CumAPNPq
fgaqozYrxNdDoQBOAosfJNElZ6cFqLRWPUGtX5iAF36vU+aOPhlhL8Ol9KfYjxTU
wvvUhZRB6Kq9k95dWLs+BlEV7E4A1T4p4YSUrXVuJf/vwMxR1ibAyMuErRxDckDN
D+HEwzaC+YVGrEyakk4MPVM6QWPS9HgaPnUjKQBcwSPEBlB2vehMcJe+lj+V1nE5
PjrYvmgBrXL0P3RTXsINMe6W5UC89DwxW9QNGqiL6VbmHWtbrMFXzJcldlofjFXA
Hsb4oMYCWLZBFM4/WnAqHHU6VlCoNm8KdsBVX+ss50ONPXpnmPDJx0FJAGhi7UWB
t3bCKtNUZyBJEzIl/4pS17D58xq9KDCPqyr/d7bJCZADUe+gv71mZ5x02P6Bad+y
q0aVFAYwVJS6G8NGsZCyewDKNY9KUEm6j5kxwli4Cli/5egOixSXZmMmJFuzIqyp
ToxEhLGR7bymshtiBKJ4LHZ0YxxmHX0p7shTTzkfGhFIzuW3RUeCRuR57mLGhyRi
749io7jF+76MnCGzE1gg29Cht79JyY+esVj2wcrl8aWpcgRtQbIqyKKSP0cpHHHi
TKkfm+Z/chmmKgT/1w5mw40ch+0DncOqhQBL2/JCw16r0o3g2mRmViixfN1HIlkL
oVZoxyeur9tb9A3OlwWct0nraIsDncnEqUDYlYVM1Ssk/OT+r/A3zPTxWOOcNFTY
uhHXtvovihAw7JMwtPTx+z6JytqCKoVrLSkdoChsNN8aCuXh5+ohckUrxAw+HGed
a43rE1H2KSZJDfE4zZQxIZ2N3MZ0ARBFq1mPYWTGeDORX4MoeqnZDkZUmiJoheRw
/dEZj5Jo+bD+NYQu2JaHLvNIHUNRCnGAMjk4t7FkQPgOQDQKbz7r8xtYY5wTNNoj
Usu2QQ/NOF/OMelFAOFRE6N6EvkQxbk7I/qqfmhTWm40XT40OlhC0VX3YEo7jHrM
IoqqjBU05T7bwD0YLFLa2JxleFxIB6xfJdhkFKxIqwx1F8DmtnsZf1NzrQdFr7m0
Qnwghy5bbOlsir5ynMnXzSQgx0fzJcbtnbnCxBOYYnRg/o/164bjhfNJDjDjkMhA
xDNmUxtjfw3ZQitapdnSaPugLyYuz2B/gKHod7YPRy1J+cAvr6HN+N8jTVGY2Ksn
pxNQEo14sJniqkXGCa+zQ31Kw7GCVnuXXk+pySTvtdejKKrK4HmF0Bw2zrVOjULy
NdPsKfngeAnXvSbnufY8vJ1Brwe8uM+ECkdO+5UQqH+YZ1RvOKFhtMyd3NwyCaJZ
EzuGsFEJ0FtdRQrMS2Ml4bqIG9Gs0SDH97AIMAijeAu9+UYxMVHescOO/n1GwC/b
/wjYeqwXCcJkKMNAC9Z1HvrIIukhqisosuXbZGC4qHkZW1DlGUjGCtf9Nm+kSHBg
PpGBNHmKW9iTWeuidislZeYzzKP7y2NhtTGLVy9Pc+ErfDmaqR0e9/S+NpAFsWI2
Rt+FcU3lbJ75x8/xS+2pms418RM206Ud8DapLqESiwlWinxet/C9PP31t9XnmXoz
hvCNdgF16pFg6AallAIuCSgA7FSLuCuKC2xS8xFVP0OpN8JucGVV1KHTi1JC09O3
uYSwVVQkyXaO/OhfB9CgaNi6lFDww9Uc8nEdpgmtZqx91WAbhja2B0NgRBqWsmD9
SeA+GJ3OaUl+zZKdr7ruGwb9EmiqI6XFE+813dHKUmFbbKEKANOH3mbHzvp0JRLs
59fBzm10r5zZOTzfO//nXn/S5UCr0jSGrxn9sTgpFfOUbs2wMO8+dbxkQ+lfj4sx
vP6QUebAxGIzkI+lS9APgp1WAKAABphOD+p6amd/9D2DRExpt9TX1aAnprr7x+Io
Ul5td3Vfdl5pxpJ+asdIZ10jIYic6WGO3ZWavY1MwasiavKF06uFiGdbd9jgExPo
HFRM0DlreJGlwKgC3Gnz7l8CzceKzLDTZHKDvyIHhaIwxh96Q8gBXhP8YSzCS1+Q
i9TqE4FRQru40+/lTr2U+XzqqCBzxA4v/Ynh2mzKXccnBUS3+jiPNZr5xuzxGipw
q5w255rQDlnJYzQMP3H/eJpSSXhga5NzDCCqccMfDBoUwuKQGPNja8557gF04vxI
3FLBKTju2U2CJsXfNGgppADB+H1Y7sUG6GW9Zc0IR7oD0bT/p9O59nrU5AIhKIPp
RnXpqTUUg3toGehLZY8gxdolpcaCa6LXWLraFxzM6R6YjKv2ne1WFUCk7kxe4YT1
6saiRYP5B1vio+cXLg3yp2GxIiXkQP7IEizy6b2M/F0EyrBKxkwcFG69A1W+r0Bv
DA9AQ6NAnnJOyzAJ7wXjBu9zsobaxoPbMeDTnoQR8cP9nkOduX7tNiwhYFq6xNiF
gTojcdKU4GnVd4KZsRktU7zw2pRy7onSrWv8h8y+D8T4flFteJEqeY+mAs+aaNOU
t1fSOt3GZ/4nj+pdyBr+NZO6jWdg+5FVzHox6WYWkv4XBuw+R3yxPBY91bTLHgNX
wivOeSEHmYSAsT5rrX/GG01pFTZcmqF3vB+xW3H+yFqD4MpKS1gTspJMfDRkS+Ej
N2+GXhNTxLxrf+fasNl5EcKdO7V/TtIuv5ZuvxmrNmv7H/rG4KSrIMR73gkGW+pt
Ef+S1/8lPPesoJZOOQyp5xiDNZScNEKrN1vCDxNkA/xxTPuppvHIVzSxmgap+2c8
fWE6Qih/oQOEw4U4IjAnEIqHS2pHfFLJOPIdZKFtxlaaNg5+uReP/9lwgHclorVb
eY1LDv/rJc1ZSAk0sYDLGouItv416FLeBnpHnENddgPcYHD/7GN+GQ2b7SCJGgWc
6s/wgFXNaP8DZDSDlGPITOVsuuiFnYNWFxxMcZhdS+d5zsWQqWPUaKdYdTE2fVC2
V+KXwdnnkY09DrF65cTdkPWPH3KbCB3hmKlRl47cUlTN0SWuQC3BuIsxQGyaBaIn
39NQ3UBBFPzaFChFviN3hUaUEkZ2GkQ9Yy77n78NS+R56k1AVYAWvGTPNCSQFSJA
MqXmlr+MkGldust2TA6mCYA9miH8i9hzxQjo4kBPJvobMvwfCmAhNh2lRAGuishn
NuJ2s2Jc9AjSkc8KpyYjk6ppd5hltRQhwCLEkdwuRAvQrLJhRF5t1tUA5EEca+wu
i3f+yTck0ZXNtL0v8I1DHBNHh9/gzYic3UxfUh0SQJ7kK1nCPIZQo4xm5RtYbKdf
/eONEOM8EndvDAe2Zy7F+DvSWGgGBv2zEWpc2MVraSDvqMAdlNZkv5PuilpYwLXw
rhgIhRSOvK9yvr+1QzUdlHj73X2myQo6nC7TyKfDgJsoyka1LKi5eGfttybEPLKx
1tKzc4TaBpFJBWVOptqimP6slw3fzRJ3b7gwxyx6bessBGliV4aTmBJXhMTnS2Gf
BGwd7DO2CG/LLxVnqxWMYFbBmsdOh+MCZ3Fie90IWQe1oYD4ZUIG7PUgoX63RuAI
6U8PFNtlSgGPxdiPheRWkaUDZAtFQnvPB72VC0OjPhgPPG3VS3mX4HJzklOrSdyV
7YID0yYZEcIdt/HC5WTpFBi+bEZawGqHofeQPqrJFtckxXHNNUHyAlhrTR96wNTK
QTrjENGMikPmlfYeNAuOEW1jWUzvcUaJo0ao2w6bVJ23LSfFVNH7l57NIUlF0wYL
zBPJfN7kvsFt1EgVZnIC3t8MpZZt/xoTN4i8g1udOEeQJSRpQgRYXLxxskMiSpQA
aaNg2sZxMyLSWxScuR8lQGcrMx0fdtfNcPPmpWxPdoYke+bs3EHvA94rZ+eHqVlH
qu7ZCPd4ykdsLKYv5MDHI0Wk8G+7HLa1MQviUEP14NavjDipZVx01XvquMd3dbYE
PcCQnEy1L1NB3IXMBYzuDczETcbMZsHgenqlxfOSQIYjOyy2955kHT8rp3lfhPW7
9UIsYZvSdTQW6IRukbEKNug6aodNLFSoX0FQJbDi9E2Sw3xhWVmyxHUJ3HTzUcNF
L3GyZbASG8gnDc8yJ77mQRYHtX/pt/kt0rAYMLrDsjvfEh40pOJ4Qmq56KZcaBZs
osWjvpdEH5cl1349OyYfSQqmA+HuDrEaLP+ZdT6q95FMhBDirTVuVES/70MH6rIL
HYVKms4+swYNNV6UZOl2s3m9SXPw5m3BDG+mM7PJsWgyBcHJflTmcWqTTJQf003g
Yd1PtCPFoCK1V7Mj3Jk4LEe031bkY04Cscsnjcc0NKEUW84Y4JehptBuSb3h1lHF
RWP4o56uh1GoTgdFs/mk4B8jnJxz+iR7P+jPh6YzrYcR1cMs2FaUGI8c0d3dT/7p
FgpDJcr0N7v/brj4vnoqTfC927+4Q0E2H4Tz/E2ZeIna2jjP3VhoMHOxpYIfF/lU
XWmKFfc+k2lUepv66Ce27pQ8jUVZSnHU6K75QTE0fTKoDg5q48P8k5Hw2cDDSDt6
NA411a0f4g5QN4BZrOmJ6XIb0knCDF1YJgI7Pt7g2i2MoGq79vddo4+gomk0E2P0
8C1oGqn2d3zwdV2Sh/9pErIs3Zx2VP8Ks9vR1V7xI6gJytzdZjUeMS6kPfy38zdL
bh1cY72bJX+073Phki7Efp6hrSerqEXXH1Y/HiR/z6AJHMJGb7MDfamYpES9qiJv
kD99RHse/BlDOErA/8Ja5POJnXN32pOQsSwrQgA10KeGtJWG148zw5ELaE1NJ8cP
JoEuTYbp0ysEdXIxdsIO8lkx4BA4saS7szsyG8jinCPEia3F9CLIWLw3uNfMVMRk
7yBwNh6QGcqCwDbH8iNbX1GRVBc2zBi/kbp3xBhBAVDhC0c/2hRB3YjttG5OutdP
fvm1eSxVoUe0AxEQm0GZlr0kZXI3kPWrOgwtpKfGUk3CPg+iV6Bd+x9dere6TiMA
WioI0qfnoR0VLed0geI4fMe69yhK8H8h7r3BV9S8Y4ntC4sjbNbpUVlktWKhK6KM
qntP12xuzHW6SNE+Dvn4aSAgDjZ5zbvWEi2LLV42sRqPkgiexX7vpXDVzg9zUYqM
24GoWzXNfgTJnn7aspK5MrhSO7HLsN1VUothr3m8fQmJjb6bktJ6LLIXZ++zJTwB
D7bQOrKCJBO5sUAfdbkWptINOOgHzZhwmGfAXi99xV8hl9tS5uvnSDhNTsqdIGtR
HZT3ScvgylYWKNYMrWAZRW2rTqWuwnHO2zXH+gei/DkdR/ViINSEY/GFZdYsk3y9
lavfwDtHou4ze8+6IV0homqj6f++IvyQ/KbFN/T6cL3IsqL52UoXYkPDZ5osovbS
J926K2xbXewUjGZ7j0diwNCpQ6SfYsXumX+eWbaiO3c1Ukr+lMGnL2yKh8hFsXG3
jKp0WOiuxc9e1Hya+gPI0h2hsmIsD7eN/wDNFT1gZKnJRKUlsqOlEO56tEXS9hPI
FDOgqAJ1J7H20t+OAv/72Zwx71/r1nPqISHo+of0MMVmzo6UDQqbF/FQ561cWMjn
3Mltx/CfwVkzAvE5BkqTK2n3sstd1YBupmMP+kCmgCEu2g7dVJyDa+5SQCKlQyRZ
z90nUqG2OFqXZguT8QQ0/IG7wwz8WXhjHVTC4PvvL2/Vf3VQ53d6EjjFc+MCZ8FV
XXuSLuZoOnKJQnJBdUOyQgB6ezGWSfiRRMKONtnWgl7hkgQVXR+nvBeKOQQ1R4ZM
By3LvmarvXR3oTjjFRgqrzaUMX5RpSczheAzWqNuiePrqYVU4e72GOyei4xoj3LQ
1LVBeJvwCVZAF0+6JPcCTDpHXRsuHcaaszrh/VQ5WMQC5u/uicrFyuRij5xOormC
YLgwaTXhGTYE1nokfjgOOqUE1k+VLRqwiKL/tO2+7zRM49lZPbRXyUj3xlvqO2PD
FUl3oG4gbs5plmYqnKQ/mYtZpdIJ7AqefUE0DpQeuf6P7FDNzQraNJKFF/0mVaDq
LuP0xpYHl0OLemTk0gzeJpf+XVr1QmE8NH1HmbFeAIMAip1TCQDWQTIU5GRQ5j9N
EyP6wiT9smm7/c7Kl4EVINpEG7nHKOriN1O+HyGhgQtgeIdZEnz55laTkTMmSAwA
XzJyf0meBxpjh/EycU/F+HiqEolQqh8RrKCQwZ+fMd8iI+J55qfeXsrpXYAGp5N3
j+anz6IZbs054JnpxM4osRLoNFH3gwxAO725SLAhMs4S9d/IyPhNgWDDNuqWMQZy
qrxfBzoGMc42sB247EU2bB+bfUsOYj9qd91RcmAlW0X4aAIKyFwCB9pnNT0gKWIE
RTJtYs68a5xSy/2MxI6voEcPPwh+PYtPvWLyehWfz2Z0LH2VnjZozz2nBTuGSYGI
pHc6edvZwC0c1OIpJhmz9uJ78sgQvUXG4wvuEE37ooxq2smnv7MQiaYS4nCtlQKj
NaOGbrWwT0mKxlevXDfwViOxOitNq8P72z8EMJ8TnaKlkkglrCF9oZpyHu/kENDp
2XAeYePz7RDNx3ZoSJ6x6uNKGTMHXbyjfU1u5mA+OPrMTxRdmP+bxqY67IoWJzRj
Q2nskWvUrldrS4PfvX3zkSKbKz1iokWnuBcMocUmYCocsnmaJCjri0HdcVqyDswp
qHtwgYggRVIt+RXiD49CY7AUfGuCjLcaZlVGtXn7hVX2U1qBBCHyo5pMvBzDPYrx
xr9CPJtVjsDSTvtl58ISk5pCe/q1xVOMvVGXN7LoptP8X8Urc1iU4CSA3tXFGvkE
XPFDU4jCMoyDw4hV3Sg7FTkCymNKWIFHwZ741y7xshRyzZFkdhN8QtElo0BgdkV4
StXhYff7L6teLXdF4IIGwaU2FUGTmL7PAexCLis63D8Ylx03vJ7pH/dDAwUB7BfP
GYP/TqtV/XDE2nXA17mDiPB/zx18wVUYx0UCLzaAod9QUvoZHyZcRvLsp2XFnqUI
Oe8Xu7KzNh+SYZjEmKbVw7WvGXFz3xZkmJrF1fVWdGHHD11qSMmkeaskIP9Z8X+R
8nAOkmUTdpA/bMFSO9eBcdGN7/pY8h/IKjIG3lk8ppc2ffRlE5ylygPA5EvRimpv
PL6NAfbMAR1ibkSNUXM0VUggaIC8LZrlyo7uDVjeHiopaO+WPeUVGYdYZNHpZcTZ
kSPMRJWeXiyLSgPg6j4U7ZZNdM9WBeOVVRvVYnxuBqlrBHJi8/xYUlpe3uKRKybS
E7XG/neFrzrIsjEJI0kMdqEXVIITaCoSqhIM04Os3sG7pHnMk4gpZ574AHhD/l6p
QJTcyMB83Pj9HDZMRmUY0nwlq89/J7xKaE/nzNt939ffZfpVwN/YyTj6bXa6Nzkh
vjf1Xrma1b34/INiqRlluOK4gm9ZM+nQAZkrMCg5pKcaVa4sVQEjtOCBcUnPrlBw
pjr/k+0IBcca7HDqsIcbQcYLYoivAnVI1xZkoMf0VzrOBYHAiwqqxl/ZmQU1bafx
2ASdXT30Cf49njn1/xhG9CGS5lQcMe+4FMy47rGPnOU8RIonz+tKMBYBo4K2eRm3
c45aZXhfLzuqO1uV/l19oIOtnB8mlY3mjOUl8fPi0AP1Jy9UiKGniBQJ42s2R15w
WHk2IrXOPglweTt00IB9fzwKQjitJpSvgUzrh/2GcLagmWmYRad5JYtY/V0f7zxn
rk+xUfyxgXYcFJPIExGIf4WnSyrNhn3m8TXIthRbuNop4J6gSMt4snF6xj/52gix
WbLjkFHfBsQCBIUJuy+rPKXuhhOqQauqiUN8nDXP6YwtyDTe5WJQYK5YKFjIQdiq
f+VfwfesGnEEjK4bvbwc6jp0ZBNcYtnolCj8Uldrs+S59KyGJvNOUs8WPw22bnEr
IvezKN8Ig4a7M8hCik+a8ZT0XZs24WOHdeMq4VxGX43wVJexnNWdecWo+Amr76IB
/6g1NGsRkv8fkTUk0hga6PjuEGB3TPHErUQnKpTQD7dBlvM4fqMGMwgF2cLBaWRR
6k1j9AZ9qFIByhOtnaFz1xLd2es4wN+LymUl7V6eIKDd9VOZ73gu31TIf1ax6qjG
1akIV9nm9KHHSsx4b3ql7XnCLcqVcW4/xEG8LJm8nygsEFeYOdalVbkXtueK9vQY
DGB2gD7jDvG4kks+N685TUddwR4lP3suGVfBDyOxtY34CqbHREb4Mm7gzyxniDwc
GWobUfQ4EWNrisBI/3/NeQZPguNB/hWl0UyNLWpn9NVdwU3qzJrpRIQ5FEW1GzHS
BVE3Y5J0IftCM8mNKt69jExydCmAnH5UEou6KUYUuNx5DO8RVpitwhu0/VvRK+4t
iANpUqiF90oumFBlgc6S/GvnEg4gpyn0xHujYZUiXGdXvolSJdU9ee//TKXN9XVk
lcG4amfWO3RknNaNhy3nL/+CcNGCOj2ujyuVv1BwJgJTUx/Dn7dZD3GLNaL7NpBe
HEZCDBbO+AZVqRrfbnEI+HEWoojSSEYt2UB/xQliaAYurfCnNoxOJaj7O8LTdA4x
a25LYJvJn/gdfpjFg83Lu6loVxUzwliRTb3jiHTR6g2DRTyhaq1yqsSbg2dND1aS
TVU/ov2/LdAOUko53XHx1pddPPzRvMWCNIG43Gvbvlqu6JBuhMaEFc3nnlmrg2zA
1JgMR24z7o/WcdtUpZWmr9eTGHlNeSuUx85qNC6QksD+W9Fajim44hSFQ1AD/gxD
gv/IC+aCLz4M+fJeeksiN7gYlR7tlhZO7OfRyy2ggIJ+6bad8VMp3o9+YdJCErXd
FjmXrEJRjL7OlVsUx4v0ZYL9SFA3GZ4piy2G2b3+79y3MwdGi6LEB5Wk9RGua4IW
dDXCCrPoLaBbKXrIOQAIs8c6yjxWGbeSuWcFSxiJ0GpbP3sU+oC/YYrxuju2QFtE
QF+MspE6yoKtLWMAqTR4BnBbz4LDpe0ZBI7h5c5kZizajmYvgWIEljF6Rj7QWAl8
G8UKCHl7Cr51IYrjvnfEuSduiRzUkqVJTqTinwrTA4Rhy2YGP+Tr8m9HjOQ318Az
hKcEDzf2Cr5AMEFCwq5qtPFH2ZdnHq8p7EwG5lwMtwMPCn7GdgxCluhJKcZIoC8q
lEcca0hik9vh1BLmeXiyVyisl940Ixg8G3jSILivCPoiYt7ZVwqtLjG63UQhFhcR
fazXhTb5gkR2emDXeVKfv8Mw7n9Cba/49Ojpxr67YxeZxCRx4JQgaQ5mt/WvnX4c
BNrOLCTE8RfgeyRrljNVhN1oUBEs+rxyOQXhVY2jpV8FQvxG/zBr+o1x3JegaDad
W/Rj9ww8iKXhhqJ+qR9rfaBFbh6HOtCPT/lFy7mdNlkjpwfuxJ73rVj3xdVdEdZK
fIg1J8o8r0mjZPp6eNHi3pJbDJo9GlEIP9aX3hKldFJ0AML8XHanYvGQkaJHWY0+
roXFwS3GQOd5CGlT2H7Dw/xV22dRyudYu7LsVzaAoACGNBMDibj5U9u8uNDjsa9z
37/TBdGhwjG6ByUxU41vfrXjX4qrZzW9+t4XqKZrYU3JHRca8+S2VYXa44hnHJoK
UrPM6RPQvuYS0v5r4pYzd7x+9K2nWBrPSP3FVq0iP38scNMGyIlHhtGylgf3TAU9
KLvEwCslOjGxDfSSvENJQ2QHZPmNIxvLuXVdfE7FU226iFwLDNx4euoj2emCRXdH
T8YVf8WRc1yeS6irlElaYzYzp/ogL3i5fAfgPlXzC3bhxEHYJb6xsiwXiRwvzO3X
o6eW7sVFKI8VwPv4rN20FRyQupkFghbLquRE2clDTsFghQOInyjx9bvPM1cDCGS8
uC5Yd0erUDGFjBOXZy5Z5yMX2+nlw3RMxsYF4SDnSqlSaFX8au6m7yv1UzUI8Ijw
ZqOQ62mhTadJu/phu1Lg0YIlRfiSaGC1VZ0KcuzDWCCI0xhGEme1VoeW+iF1zzjx
xvEfVpw6uQcjEYS+gWc8nzA7L4vRQF8poe6wf8tDUqBukZdzU7lDWCuBikp/4f8m
FW2I2PVNvY5KuTWFW0y8QLnCPIA6kUvsZZOdbGVu2o2IkHLHauwtWEJvjuGdWzFI
juTEv1cNqvgTWgwWerOPN0AhkCLZXnRxtKoeivvg5y2ri9Q2Lq/hLfV2MpQRBZm7
2kNgv9/w6lTYYA7TEXbh8lWrNR8jS5Tu3iIFJqten91MKPZ/dEOzmyqwHjk9i8Bu
+6QaL0EjUMfiCJtZEtDw1lILx86VURKElwJp1j+G0DgVlp0cicmuA9L4/uhKq0rF
yUD6+ux3PUXb8IX4LTH2WGmqM9V2HUCFt08Z0oksj+mDHL9yC1ZYagIBCK18zb0o
pUCS/DE4TnndbrxkyFOs6ENtUYiGWxbx5KbOfjkO0pLc3mcCAF0MTd4hMslwQGwY
SxbOWSnqWR7qOWOKdfHln4ty7glC3800AqTnbdL1v9s7A52SyhafPUrXJR89wcnZ
BgUbUKxd3ES7PfRrz1BAxdpaEPUUE5cUNRUNgYRcHltyD3TaGrK6YfEX/86/jA4I
dSeQnQuDqAuNuIQGowzYB91vakMsh/+cfsd0tyWzAtIn1utiuOLiR0fCwfafhH3t
oPRLVpKUV3X8wpcnIvy43KPJPQa/7SDd3e4NTMhWgVso7OMLaEITPWJMhO3IAWi7
p3RQqPEnjq9jnRwPO8+cxXT9vvm5k3rFupveINd28jWv7T87n2MsnAo8tJeYoNIF
hnD5pU0TAv6lXN/hz9z372OU3MNqieV42yFTVfUulSTuthBmnmQ8O3unnrUmJmjG
lo+JRAZFe6513FlrPa/pfUw1gSMMRLGiE1WWRcJsqgvwU/cAOXFcTyRQGI7ycs5p
tkCifwt3L7vBOhNQGZlaUqGCQypjPrVk+oA0lt3jZjF/l42g+AIuyu7rHtbTTRSn
AR5T+uDv/pRf6erGQqDGH5v4WM1fMU9gMlC1LfSsdP6mLEVK9K/R0vkbPm2HdIDM
dS3qPz5b9Mo6Uq9X/qmJdBzbOwzaVkm4vu5LV5C85vp2dtSY8ezpYcKCEFvKrbJZ
17RigiVltuhHHv+OLh36SdsQs1c9NFIDp/0Yiur6SyAD38/f/TgWA4PQWhrJveLk
VtTVncroXXYx29Oh6B125rFlv+QV3R5b1bpWQzt6iNsEprUcYvzHO0WkEZh+uLo7
XwhHUzcabi3T/9GTsONpHx1X+XYWGWu2y3H+PnWClluSUcmSDr0wluuvspXnQNJG
3P594K7yVqquO20wk2AAWKHYC4rZTR478BWkRIIo7jjrYuJx/s24VqCh5taWIQA0
UMHag6tMZ+Fk0CIwBlR/RbAdsIol86ybu2CYi+wTVDhqn0tD2ZrI4/elaK8s1ZZe
tnJelexc3EBvrvDWyg0gZKnDVd0WGfz6p4Wjc0534tRY+Awmnx901fV8PnTE5J8N
pIJJEoJxh9ROxZkZ3CuTvr8DVTNZrsbgltUnIjmSKg2jcH6NMUGZw2gVvOAXIPMx
izJxhU/Hi+PrcO+vebVObZCPCFgNvB2BiBnpCNWhF6LHiP2cU/bL8aCYF9eylR++
KZszgjny0mYxGWjtn18tFgPKnpXKkE7X6jomZbbfUSFwvCrFDFcrg9wmMNyu44Rw
vzfFHtALEij3SzBRePyo9J+PjJtW74CXc9b2uufoilR+AOi6B3sbsa85EvYglxdB
7jN04HcnS3DANIdXgVKOrdpyzKc9CL9xyDjMTQcKSu8Ks/x0pzXgTPtjyVeqKnaQ
Dlg7vS6lLDf9oxrnumoppjGBJqGHmAQ6h5CfT+aPUBG+vQptGbGp/4lja5tXY4wi
+nykTg/IJMmw39zfaQP8l1VK1DhQjreOe4KEHFUF+7QHkeEPC8wvTnERyXvbHVla
9A1ffnQspr07cl/VTGmmsP/+grpdiZD30MdeRqhPXcMJay237npFr0cvRRCKBSQS
lslzgew81/EoyEMFl4zBGs1ukgO1jziL/57ylWLl9LzEj45tDknKcXmRLo0pzJ+F
3u64PcJXiHA8hMeuopuUYBL8r/uHXEpmdMW1BPDo2/TDhq9hAzzhzDa7Jfspvwf2
ex7Us/2cU+JPEdNAOQU9etsIo146DibLlTwBqRNaklv2O2fpgtEO69cY+8UzSAlj
FAYDWVrTm+pbrBQikLEGGqq8KwjManVAWxJNGH74WDbUO3mJ9U001PU//zH4b4aG
0x35r0uroGMcf7211sZ0IX7YEbqAtt599w+8y1RYUK/tgiBicugXu0YlglmvkjlH
yvDwvOUpwlOiXPhxGlG8D8lx48xWsvGjw4/ihdEEL9m87GTjo7x35zH5Vl20dybG
DRghxDzQpVcfQw1MI0PD+Fv3xmK2UzxyB8o9EnjtyIwh2/dnpKHWJUmc+vIeXIGf
StvmWiIRYKmkpf2jwo3e+caTU4119uD0wgDeremlJ0Te9KR/QI3om9UcnmnnH60A
oB5YUZuqNKhIOIqsgVPgZZjiS2LXrcwRud/sZje8ZVzh/VSpUW8GERW+glMgtzA1
k24Bup8ZDQlHV6tWLeYeuj4ViA6c7zbU2h9JcHovj4aDnVCjvN7e1wVYexkhAyGh
higIP+0HiZzKfkPWI5M/t4LHtT1gVOqG+OkCmzp99By1AzPKJ43zzmjOjAACdyyi
ZSmcDkZpjZW+Oi0NgHuo9AWX8M8PO4i9lEJp/vy0D7W3XfmZBZ3xXde16gLZI41Q
st327sroZ4Sg7mKRegqcdIlr6EHBOdhxbz6zBH90rQqLOXLVJo0hsduVS5G8ZE2Z
mNajkNLIfR+Etc7pFrowdKrce1wmInKAn4o7StpdRsOA7AxXSAIAfSek02Q+7PUj
AoEqOijns3Ax9Ew4S5T1dsX951HJS749ALb/PMD+Ll92raUstkkdqM5X7fDTsoOW
xGv6bmybzs2h6kQzDcDC13CIITWWCPlQtKAK87lT0TGCnywpLMW2H5aaGHrw7rGS
MfUbXWKDV4ZQU3E2tRYX6zlHlwfVOf14S55aG5fu3/XGnatmizoWCgURmzvMOmrZ
1XgGPICu5wDcvIfCj0o8DoMrNm8rc9oE5T6eX0BzKTBaEnEvsgy/eugD/DjCyI+h
aORtFw2J4QODXt3t7NqUWEjRvUkzUDUINcIwJ6T+ogMp76HH1c3kgWeov9kMo/pI
K+as0K5SJ8I0vXB3Bm2c/5IPsne/ofhy4k0MFl5JQHmS1/+R2kbfdrR7aGh3veoa
V5MahTq70qkPCAYr2lSO9gIXGCIXLzgU4v0oAbXEVo+hTaGxiPovVmM802/DdOzF
jBeBYqur1pOxfigbESm7VFoHWCAl7McPVQVmdJN85sTaIWJqeuIMBHk1dNd4bkaV
TYu7qP+UhNFMJ8URwt42L7gzNJ41rldmYauU+x2m0KrLqX5LkatRaDBYVPHhuh70
o5ti3AnpYOqugWWO2kgWY9KWoC6O25YRMnrbj8cXMvbDqAWN97mVC4AtS0OVlrcG
GT4TdQpQNk/S4u00BX3cIJt9W54+m/QpmASKgRC6LuLejYh0AJIgNySyGHvvoLho
TDF85fFzTMxZnFngXcteB4gUWMLwPZxqsAX6FiAPTEm7V4izIt6wXuxCp3NFVkTT
0Uz/q+AZuTVcRP9yPsx4jv+0OQZOQUzRuQ/uUamdzJer4B2Y18mhEmI2Hg+M46CA
4xqb1Drrr+MGcaYTi7O8c4gzrPulWjXtm4q0DWzybyJCPurVCakdm5DrsK0ehGqX
4ggSrsjMpUt14TZo6AQkRUw8NfWRymqSq1CWkDZezdOjMabkuDETtFTkP1pIcUD5
Pv8ARuOmpDUjixcjypgPPpPGMDUFS3b/O6gMn+T1O/BcrB/mJJ2Tn25hk26hJKek
Hk1WB3T1AX+MrZ4vvwFCwPiodlJ1FY75HFMyj4aBVcUL6Ld0CyEYDVVEDyUS68fI
K55vo0tjTVUV+5TCsMYjePPRbrIRj9nYZf892bRXu9zefGfKrYq1o+LeFFGWcBXe
W+A/1sDalA4wiTRtqbQ9kdfAa0o57e08X4YRukZHx6vMm106CT6nOJqmcd0m8DQj
XODrXFShvm/VLnXqIWb2Wt+U9isszd4xdWfXfCV0lJAUbWeujMTiNVdTjr73m6ms
sUgDk0zDKbMdOr5ZKriNd30Ip8GkclC2kUPMzi1syveTM3gxpPwHsQJY1cIpOAL3
6kRnZsCJ7KWatIEGGkiNDgidLSNb6LH2uzFDCXI6weTcrW9CwXnz0y/zjNpEa2/M
ijXn9haidmF8DOhuYeC0rjA+eLzDcHHsldZrHeIKbg9CPIeton5k6B2EKmYsgw63
UbWjRP31MzBY1h9Mhukh6P5JAOdsVs4nj7ZNOFDQDqgQVVDArPFUGKnemir2afX8
AySBslonX4DjVpzjqp7G3Aoqm6tXpBFlnvzLMptU7paP0Bb2E1O8dho7udGQSDED
3D2X5qOsW3tVN3+zn35lexwjPpEM/5nWWELdBIoX4dPjjyDVzyBw//iH80SMS5M0
tkUaaF0miSwAesvVBNjGZZ95Dx/1SLPABkeq9vyZDjAvskiawtm1y4AX8DTa6ySh
Xz4+rTJS2jSdF9dnZPHG8Pu4SDVUL6bNXk1Gj3mPpNMyU6LgQ1fWui0m/BwcRCAA
LxQtxyr6K7fS53fGqen3/k5kBRJYx+G77oidGhGj2Hx7tjoR3rf4enjjI5Pm+91U
PvUESL1Px+tfTiZoTmv4d2yY5e7n5E6sqNV8zUDBq7rT9p+chkfluRR1RSgpFLhr
bvLaG4gGBIMnUgEx1wgXzrOQUKexV+ZtgcADnS3QLO+qixVeEEUGiwtDY22exvRV
/2+XlMCdwzTBVT6ASrQsDa+/ppbCPlSSolF6tE/9lhEi/b0+B3H+NNE9hOVZw5C6
7nVldMr9eFb1a9PyH2ItmB5u1dxUYCrGXrsnh80atj7nqxlSwmF5yQ9ucgLIs5v3
bypn07Q9PFlFT1QNCLrJGxcf1F2hM+TdOIc2EH08oIVNv0gsnCjiskJJH+DC30Ka
s+MyJw4FH9vuvZMNQfKbM8aUfJAwrx4XTblDTzsSAbayDDCZDsfcKpdmt2SlG3yf
Af3MUGZm+csCUyDR126hOTJUsDIXwaXdOxOZyf4fxOrEtl7MyYv5L+5YnWAju01S
tlG5Ubt182lyCzpOVq244JICbQVsoISoa9sMidMWcMVm5w28XPFdhcH3IBuvnEkX
XR2ob/NBC2hkDSZGggnguo3qwKwM22tHMAuRkTrIC+DPqWeSXP1btiHtR6DwOLIe
boMq4iaZbceeHnVzB89GRSDSimL44pM2COb6UZyHgBIZ9F+ymYK9qOXQIXsDWNAq
AA/lbhH+1ZPRpfjqJmrOEsWJOyVy6TcPebxBBBnyzCgGEUem9Xvhfd+t02a51QAl
Z398VuCULpgqYYUcnYodeb0uYQSLeEkIhoBaAySfQ4v85DTSHq6r7GqatTxEQnq2
b36oJIbbLt+591gBTgPTIgvVCXOLzMWpBoGN2mXy42VxrHHRXzu0gxOQEw8RW3hr
a1E0wtzEo6Qjqpusq6DNpHlRHy9WQUz4p88Udi0ii8SXTLZDvpHyt81xM9tetXXn
Lwes12Q4CRRzhBpS9OoJebJby6tb9vWooqiP6e01GkLjvh925FGkNQ5J6n5TvjSC
cjFV8PxdlJQmXWA0SSobq/JwLOaNKNmO14o19EOk7xxUNDPiFKoL6cJDrc0MTvhC
8G2m1rod4gkUSQPaaDnLVaONvfhPoN8rQolRU3dnEH33oHaCgkrPq5UdaBn+gflb
+MbB2x1OIiwGQQzNSjFogwIb+sWi/GOJPAD0OJ/QjITqMD4gzXwkLcynzQGH1gh2
NzJFh65wFJxi4XJPEV3zS3kuMm9eg52ugtPkGyD24UrX2RShnMxN2zyPp4RWKSp9
1PAS+ULnqYhu/4ss9JBc6zlX1vCEhEfS8NpptBC1PMYxL7iCu0fuAUbiIE7bPUw5
VkxE2fMdM2bAUP59ZOn4Eb3c4tvxn7pH4L++UpgexD++WjLFH3Hexv8xjARpC5gI
9QsFrEVDV5z0jz0OLoJ6XIVMGvxD+PR/ZkII076HNAj8i8WBPRR/M78fL/kRgrek
Fw+kMKcYgiLtu8mW8kJxc+9kX3QCM3WnIylFkX9mlgO44r/m4w0JKiE4ra/oGTEY
YXCB/eQ6Ud9g/ux0fNJfTo+qahQ0pDQfW0pb+i8arteCPW9Z5KgLKZk6bGyvyhmC
qHa26LbMkC3b7YUxLoL56jm+KV/XYvVUYXYcPZwqAvGXXyYUOpoBJgtmNb5/V94F
VSkohXvh95ixUaPV/h7CLpHCCabue08FMARbYyymiIiemF8ot1dIaYyxHLXdpGNk
q1i4X5byrMXjB6OSG+xgwdMXNtM/YmkemxCAOJO3eUJO8qbnkdu4nYBh7VrbmSn3
jXY+fpPG6RyLVacFJbsg3zeNj+nFM0wHIbTk5zXjHQ0duLGqlsxkUkzcEFkanW9M
LwTq/ETp5stP9j8RdQcxkwFG/6pu9TlqsUU1+NssIteli7wMGCRmu1V03f4MZHGy
Iq/Suhxj2LuiPOwgJFYvqeD+tbd0nuRbu3/hF21YAv3+RorOJTSNmzl01ex4jb9s
y5r0Vt2viEzTk8PvgJjtlqvWE4A8z4buC8223N3H09COLG4xY0Q+BfqnxKV7aL51
W8/QPSEqy9op3g48/mi3bFwm4/lOtLs1B121pArp4/rr+jGiSOFVNJ7HLZEau2vw
rvqoaYDOnp7VKggrg05ya2UtYBauArmvV50FsxECI9e3Z+Id7gcVlb9MEJ+eaXkb
P1bWE9p+SYkUEgJW8KYRnyn8X74Z7cX6TF8wyvPkLxREceKdQWYtVp7aVHVvPgqz
ozBBSJJQLNnh7WpZnvX0nzotqoQQYbHsPvZRyQJmkXm0IvPQ2xkC/+va283e2Kxc
u5Y9qDGxjswSsZ3Ed4iNAODPMIZGbHxHTjfW0PGTCPh9DQ/Fx47gM0SO/UVk+SO0
px26A8l19Uht3dhfDEedATIuDpl1rf02g0DLDn3Ok3xQ1jjtugmrKs+zgEUsy7IZ
uxYSWEwwsCbqK1ldKKQm7LlhAcKPapJnx4djarSUrBwZdlszneOvxG8UDjInK91l
VVOT8Phjcs7jpFClnnZ+BbIjs7lfXGovShH7HYTY+6pUo0rZr98JckF88qAa7lDY
62AQMvc7WHz9yQi15iMdmfwsTKSmyTBz9mSEtExwnFVvkBAjREuncOsSV8A21Pme
4xTbmwq7vzvNZWceL4m9esmB/JnsikOpwGHeag/qXgf18CUpv0G1MBqw/8RXRWh1
4L2YA7xmwt2hcA+Ak/6+km9S0UUbX/RBa/EY0R6Q0DS+GTs+u1U7KQKWLJDbVyb0
zWgQzYwUWiPqDCxU4U+iStMHQSinDX+iKxgxxv/3TDMQXO/h7mUUMHttsrNgRWn5
XjH8JxUDdtzJtBy70QUNyIJzElznP7SD43o9SVvlyDInj1+7Kr0heSps2wZ/+uOR
qOyxnrB0V+fdBtFCe9ELMwyriO+r3slNHt8eE9EvVj++1JvgtuXvkXt86TFhbHF/
oynbd4Or0MxCBfIuARUfXPq9iRnj7p4h6K+qcR2Oi/rsc45wAAckb/xfbkooTJ8L
YjWfsG8wk549oKZxXHYrs3h+K2FZQla4j47BSACSQZFt36Poz2IAtNkzDKgFtHmd
SJRpBmPG2x3qsyFzyhq4HwUarcff/aBizo/14jLqq0NhSwMJIrgQoC5Q2YMUGxXI
5EqY28Z6+hvu/wHMdHJOPRw5RKpccmO09ChXEwjh0UzpIWRmpbzjF1V5yO6tr1LD
jgQ2NtR2P0aSVEXdiSisZJveSSB6ih2NqS9O7BNIOtii46JQYj97LkFnByJnZw4w
4YvutkFGMoeDv6SGCq0TUQ6NSlTEVttGy1GbpGdZsOZDVxy0g01q0RO7yp21BOns
/Fkx2dV/DuT46dRwHJFd2+V0YzOftt3m4Y5TuThQ0IZZggVBmxiPbKoCcZJCwH0I
OijzNUTRtJqvZy5Fes+AzW5xlVkPpm/xq/KzHeeAG4nfjY30SXIMhx6TXS2TWJ8U
Rhld6Lei9/yobsbkGAwn2Ud58cP0SPveycNLCKZs2hHRPgovs7fSCMbIyejxsp/w
8ZeZFH3CK12FAgU/geVEDgRys0arprs6qcgnCpRry8pxI7/DPiS6QRfuVh4F7Lrl
QMxfRl6O/BF9/mczrFO7N3mVRWNg1HBTPVjzU4tK79A0oXasZ4TimVBzkwelvv85
M2MWPCJ056qIVqVGMBiNiD8MrtYrl4WIgP0HX/XWtbtfVhdmyQcBxn8gmASBWI4G
Uoer+f8B7/HG0IORlKbkbfZ7uVyit47rPMN4k4yMVRX0pU86MfNnKzyt0ztC+YHw
IXjRVZ1y4bwHZCFAvjVt0Cip50AKtNcnhh9o1OM9m1/ceiP1uBguPnlXKT1AX7q+
CmgR6eDTP5FkK0vJOO0/FwbHhwnOuWV4LX9gomQNOSExhRFUBOY9QVw+SYONq4fN
Gprq/iTMoecSFb6EewFm/a/sE7i3nZ+TDZgFNcZcNJgfRG6nMu2yTeV/zG1zzAaN
QRR7/LsPaNxE4Nyf2UL5nViDP9A1Pv/G1FRxZIgg3Gi0WKsqV45Mw5H1VCDalzr4
p5H1VbTpZV5PfuI4s4t6KAyiKXC4T0flo2+edkRnJxCP61j7IS7YJLDvXvZFK7JI
8Tv0zgY8Ow+4Nn8lzknlrntMFAdApqH7gKGtbucuAAzhfqqabA625g58kqBQFBHZ
tP9IXspc82zybDpU2dsE06tlO3o3vqd+j7rmWs8sm02NycE7Ph5Hiyp+7W+KdY7j
VVaDVWyH3u0IQXn5wCyC4GisM/5AD5SYrsQTW2G+03JAep61k+HOd/mTJ0YbsXFo
OChWQobMgc5Z7TKWft9Nzcgl1POBWJeuaE7KWA3nFZHb3BFk13KyIng6lNpRky94
Ny4loH8jeRVYbAZLN38y9u2TxhXBieQF7gf7RebX9OZLKvyMFJ3+Sds9PZyTue2d
fnYcdOqmMaQfsH5ofkRrnKOi5fZw/0vUsXzBWnCOqfTHWGuTDvJ8reLS9A7TDMIU
B73VOr/NqxpiMruasxYJ/tSzBQ5XN97oJpS8Nvh/JnHr9rpZuG72VYHp5LZhhZLD
ii5gQCYSA4YUck+MTfvzxdMmyx/oeh0JvBzmNcKhyIMxfUH3+/BzMYN3Vq3rFnoi
BJOi3GXFCebjsPhwgf6QemYMH03e9ipJwVw6j49F5fRCV8HjPZ0L/Rp3Q8WMEHLM
tclAUEaqmV0fhWrvUKyHRNJpuBXnYJYrHq0Lb8I1Id8HIsMKiFLRFtSyiTA3qjbV
OyW7MmkgjhlZ7vmd1YZuAaMv9SO+HjxavX02NzvqK0bG6QU4PP7cm1UwgcyhWBvw
QvwxEM00BVo2FajT/fISnYHzJYIGFCPHlJhkL6o++aMUGKLdkNgbZp0T/gv6fdDV
8X8/RaCgIK9lkcmbj4u64us9XrX+fY8AQe5P74ipvtWdxGhFbac4cdPyhM51ilIe
X3cfR2IzzCn4OxEjcpL7p3x3HQazawthd3YFF5Vz6UCiqydskM4H4GDltkUJMqiH
QVN8zMRfQgxeb5Fv1gGqJh/KmZAxTyfGG5sQtoShEng1kEMlcoBh0TcLlXwF/NFH
CcB8pWPSil9YZ7qNHl5e+LN0UTZOjXVuTs4T/vvvlLIkqfeb2KKirgnpIUoUPACg
KGs2I58luoIunupzcxtI2fe5N9vxbt5tY0RwXpablMB3YRMZ9uhxqbm1dnXrj7dk
2N7aa4rOKaP78E98q+SPbVSL8qHD6vAro0s+p/g3aRzplYioMrzfInlUUQQWq+rg
6IJck/jmSNpX3BsncznscMJm6RWwZ2ZvIH2f8Y2CJgILWizxc/Ye6UpW7DwbgYYO
g7hdIWigHpmUdJDuLqUPfBh2sRQYkSZx2gqOnQt5gk9dRkva8+Fo26pBPFI8WLUo
nlXPckyB6k6Udydl+KJmK7zgEmX2WyRcscc1YfIKaOv1N1ST6X/UnPb64uJ5mfDs
Ck9bBv/hg1/+1G38BeYfd6t91SLWDae4+tf/vEauo40940aULU23858SdimMUSLn
uJz+gBpI5tHkNOtccU1nWrcdRNBqw+SfeaNL8aRVfbzgod9XkFpKJpPYtESLUQOB
bxb8BWTX4B7YZGJAvXGyqTNuGcHMlf90fpcRq9zfXVWplDXvLEwIio/4C3vPpxkZ
d691In22n8r8uSIW+8Lyb9OElA4d07cD2gzBt9JzNb9vPjmMrdjPST7ZQIiqlMvm
ejD4EqZ2Qph862rqTwC4tEKVPyYj8vXV9YPlA3sTiTitDwyUuPkdhrFsC3VwnFMk
Ts8sAVrTgekrZrw9Xv9qPVGPH03LSTdE3T2JDoS5sjfiOzQAkSluIQN4KuBrFi+v
gGnVeYqeRTRKAn43aVHvEGOqco8xeeB3LMlOsbHzw+tpyF4hCnt0vJ6QNRF0OC35
pJ+KQCNBvt5SAZDFuky9jQqblrVyityLZKkLF22K59cNheenAW30RDrBJ1lZhq6U
D3krlCQL4ynmYkPgYqYGCOvXf/QqPQ7wopS/KcvMTMjjdRGHWpNElSEDMmp5pGwh
vxBBS3zvV+yZhqrDnSyOl8dqfshV4iV38VAuPKrqpWbYpaaq8KaTaO1RuS7acGtr
d5zw8Ospdei351aIL4AOlPNFqlEEbQxj0YlCIuGs9x7bnDXkyOMiR9tnppdXerxI
2Mdsc6flXvOnONwodFr4Q20jfFCMQzWp4kWpbNbrrlTETeI913X30paFQ4n7GboJ
O++zxg4kA6f+U//65irIDeAWs4zFXbva/VRDVRDrAcJaZ5MsybcNHdJwaV0cUwTO
bjOmiR1XbylC796OrPTfUHZ5r1joMYAVylovvTAYrRs1Fkb+voMsUcqZTN+B5fu7
rlC4bJD9t3UpQxttQVFOP+NI6Ey/CQ3yY8+hFo+rE+RefElBb2w9/c8gGecUDhCl
1e3vZc7L4A3Fo9p0P2QpJ98AbVKChQwNI79MyGXLDaIQOoUNcV3XnaasOGgArI5Y
bpNxUOU+lX7cveLRlH4Zw7ndyB/kyXJtz5EizxZbCPPBwL3onuYKB2wNnWC0nCMW
MwjfPtQVuQW7nkdCV6zUPwPuJeW5MDz05stBKJtnYOQGGGWc3Umjbt4G+++5Eqyi
fw3I6dM+msmcOztVq49mWJEOboXaQfD86pikRoH0G4Wr7W5DuQDWaP0L9zUHdPJz
ExduCdf/vnStRzmLv4afshtGahnnJIZF0laLA3aK7l9XmieYwltEcU3XUNHRKFiy
6z8W3x73rXIdihAykg9ccuXtKR2JqtkRKjl6D1MjqVD1D8IJgHc96dSVzMwNvR4c
KPPW5MSGtVhryChQnbJZA6HgqZ6SKrh7um/uPPzgXzoA400fn+SYrChW/38VRCac
RubejedX+HTTA7rZcQn3rij2d1YMF0FzoT0lnFf2E9dhgWTYgeUsYEwouXsg3Zf4
v7yChcaWDM0SdCJIVgG4P3WmxJ4wwk8UVRV61jNsJQCOa/aqVMz4C3RO7LDudZhc
KlrLeKY/X45EAJkOyX3/OVqdIcJyQAbkNyg7tQEFSHry9ZFT9tzyPfufvH+tzsqz
T6XD+/mGt1rKhEM8iV4IyvSObXIbO+8sHNm7SF3YboK4EfLkVS6Cgn+oM2WT0ZvK
fEbgefMhSuSnT54MX4JX5vFFqYcstDfSdLyKuTLUg15yhC156mBVpxv726TkTU20
kKHNB4Q6DnvHQe0yvOleFE69ssz0RhLZFitAo10e4xlR25T5+Yrx6MpaRtXJLI/Q
096HEuoG/eXUHr0P2g0uFVRSrwiEXhJRgFvSM9n3192qGGUfRE+zEvQ2ZRzWVtoT
mkPYoQ1VNnJZP5iaYFJV2lHVieuAt0kITVeAUym9ADmWB4aj6sMsIDh/9MIuvX38
BdXZBiZeMnOcC81+A0de4auy1NFaMQHMjDc6V4jskHp52g2wR2RYoicyg6JDh24U
gk9fmmLIjoh+id+5P8znq6VA5qDEUkFV9S9mBJXQQIYzMDxmHmJ8dZBMwBKRHgzO
vDpjb22fzAVC8yZ/je8dG19POZH8Xupdci9vy91Ox5DG9+89wRmVBo5Li8V/0y0P
ocHiVdITH4yJOTfr5rnssFnAiP8OkApZcMUXJrMzjjq372daksuY8XvYXnjmfHSa
ZSgShQ+Qmi7cEKCvbPNWKIFLHX9z8x09hDlwklYySVBvHN6GVsKgoV7xJHo6ZNjX
yKcQrip4Dgk0aQEz6cbqPmVE1Q1P6NzSTUm7gP/tfBWVXqbJfkOze3dZN/zny6FS
2JjMUo79j4mfZ+ZIw3P/1YEqfIba8qZ4mlXIv7HCKG0k1nZsS6n8bbx7HummFaP/
eg9Rez7oRWsBhS3p82JIdvlnY8q+dd4QvLj04AzplPQvmjowpLrnsDFyvq7ngaUU
iJ6Ko28rax6gQ3gNHfer2YSE8Chk27NVqUioEOKqNrf8foDenDV3dTEG/FYyFJbk
C/axxOeyQAKWLzFBru+19wQKoDNA9E2PCz0G+PJ69koY0dDCDylBJVGn47K90bpZ
xv75haJkA51aSlpInfwfIojVw5wQQhw00tzmLAlHEn7moiKLE5C1nIMoysIEdInD
pSEFrtyFM0gQhnf445nphvYkKDnLWP+rcqL7giz9KErXJsm6FTmgnu6UMm4Ucgrt
yRJnriIUIfgESK7pOT0n3j45F8uLf7WnyI/1Ut9X6eObISGIMtpocDnczk5He3Pz
FG5KPEOa1TJublmJAXt8aYcoI8VermFYOPhww5dud9kIZlRIViVcqL6C1dSleSeQ
FqacgnWNLDLWfK5jN5TSOjtLSQE3bjeKIjzoodmth80yXencGEEN6udFnDyaCjYU
ndeaIsb7fdGa5JrhsZvWjw1Bw5M7I23QPO/aDTSSkOMWGDuKL6jnsBN8ZGjUIENT
w6JKLhNjFwDM6PFJIAOyLQT0TRT8Be878i2decu5sv9eQQXiZ655IYSeAFn97dK/
7YvyXpEIWk4XdJHr2hUzFXiuz9sAlH+s7S4OBZSS/Aueuv5wmc1L+/7M3LcfW4HF
81+O3FDjhZ5b0WXcryAEKpgW17DNz8StpdBqr/r+DCTIMqz36sfGEkI/P+4lUIbl
ayjw68WJAiMLGgLnNgD9zRsj8KCvM1iUL5XGSyGGhbZrmo2WUELE3CXgiXgqOqsp
B/h2T+T1QxmCQgJyZWEGdxa+Zb6uUekV0F392OWlqXb6s1r2H77jtyGIUxfUnFAM
NBZxncYkZdsklegUVsOc7OnjmH0PN8hYKPM5B4N5WcgVbmaMr6HMY0blEhkNOMtE
sU4skih2VLe+A+noksf8UTTpgPyKDfI/wHIiPuI4PEC3Z8KU4tUVCemOW4KWvXMX
IejqaNzvHsBTYd2ghm586ZDm3KBGkmilcRppwIShugf6eYKRDuVDVjAb1np/Xns7
2gpgq/BK4aOuGh2sYvbrCwu4Vwq1N7rVthNXG8tTENh3OUQfJQlir7iYE7sDGwXK
XqKNZf2oq7GLw8hHUmXaZbKKlJAun9FPhbYxkY6vFztWmisqhzIqEGVYNf6u0xfS
mh2aIMhB3xWobyfstmgmAn4xt+2sJC3IIKuT8eq7dEIpfSSe9U1yqogx/9F9rDsI
ImMRsjiX/hoF7GL97zrKRCHCYtRW5oNFuncb03LL80xJLn4/mW4g4fLJYgTyAu6d
QiiPWayK/zR2I9sARNj1HMOEcQk520dvU5joKBEUKhu5O8gkzhOxB89pzDEZwvaP
H1ZOU3aYdU1/OrMKXNfFiH8ndIg9WVc1l6/He1KD0UsjXH6FK27gDwBaAVF1uB7m
4z6QdbQuN0iFj93Yf7EUCgsJzauFKReybMOqOi7bVTl/sV5ALE9g6jaEcV4RebUN
tduvmpJYfll+k0SyW4VTA/DJrEnqJHKTB1SfEsXfi72UPo23GGoAJe3+MA+Yej3A
+3LjHGiN3hr7JQ6C6AaaV2DUYyZAGKKNdiEwnO3hTZarkAh6IeBZqHfwdUDpgnzu
RqzS6styvR4zSNFtihA3cih81nO0X0yStpwn1dHPbGhotx5KMdY//9vEs5VZbV5t
51/TbsojXRVBPuLTmgWbA3qgDCD5vcyDp6Kd8kyAqnuoDlDOHt9lYVueELamibV3
2RIEEXq7am1pwFNsEDsAr7jmgt9MefoG0wYkGGma2lfLUSg5GN8n75vna28v331I
p1enLWaHfzD93wodxaHoTNJri97E8rwfA6uojMd/nWqpCmF0iUwTBnaZhRD9xXkc
ZkMO2PYMor9xT+2an7rNnw/wYA/C80P/aQ1G/F0bPXQ/9vVJt+HUxKOMSGfMKGP5
8/al5i5Zq08gp0v3F7DW37rZSRKGYE6JHVSa8nxdT26Zc/eBTTtHXDOciwbjlyoZ
ku5gvFy0Ud6+JPEMO3uBzFjJattpKjZSv947RP9DTPQ+O4tsmMUtf/ehbX+CFPhF
anRXgYVaps3tQkeMCUjJaIcN231MWfw9n3dI4aGNDAaE/BOZTvcj2dvJHgoWDMBL
CDDWmEjBBTT9ClqK/AONxBQ6arBRv11MBYf8DLm4h8ycy9V96YllCc/wHaBOHHwZ
l+Z3t8GJM3vdHPPKttrwD7GIJv5VfYpST4opwK+plEObicgyCB41cwGD/4mvFCFp
zTbLCK8lyi8Lozlw4SM/29ktsZAlhbNPmMh44i1DEtSLQSFVklgDQQ1Wzfug9xNG
J5n+4U+oNvcUHHsjSSamG7rM6LPAOo/Mb81/SnB3uEFdqAyQQ4xrw/g2MoLF8Eoz
wPA5TAEwKyRpG18hC04B/Z9TDZ4eZgZAHT7xaofNMCkHc+1ljt3UQesjGugUqac2
ipFMxydtWdIt3t37SF9N3f4rC99XTVdAmEzut87R9/TbT/Zyuv83rI8FUuPSLXEv
8BAqSFrSkUdT00awPqPF4QtQ3tjA55lRO8Ytk7oQNHJUXZ4LDp3jdfWQElM5Wf38
aiYC9vHeAbglxEg2WvTWjbsleC2TIduz8aT+HJdRR0ahYaRDjT98gR7FoYSukOtI
/9rUyLUVQD89VOvLMB9UF5NCX9wA6hMInBt8e2eqNLWANt+C0iuh/cv/ItsLCyCS
Y9M4/ICxgbBfVEyuyh61t7cy+jDpAHZOSpTLJDXgJDaGIY8on4pTBUtZhk85LVSK
KrEAHd8bGRZvsS98z+aUHJZykC5/v+sUgxT7VzqLs5VtxkcrbiQLW+0d5qaU/lEO
9B8vRZIi84Dz3G2ur59iKDbCmkSiNxz9LYRd3sBK+kD1TNTWorlysN0YXfxHp79r
g0WLVnJew0oeEztoySukj9i4prmnF4SPg5QoR+7vFd/2g7TqnEPiBdgJntzULHro
0vKwTj4HxZe+5IJObZrvIIBxavDSsgAoUwwC+ZyNxUPCXYHJ5g0rfOE8NxrWnKvy
v8OqqDgPWa1MHamZi0/FhjJLXA83Xb2uMNlA+dUlUODUgHSKukFIfzscbsz5Py+C
zRpICxNJwc016NsYsh4+PFfsahgpWZAynXrLUjSZ0sNkGMPWdtPS8xXCvxOoo0bi
OJ9ucr3nzm6ua3wbM/aBF1OIOK6KUwO+70wYoFB/aPF+tDJvTcEy/S5emh7gZEgI
ePfeStK5KSYHq495mjux+KaFsnME/Gp68MIIsMVBk+ArHgwZ7qU3pi5cExZuc2YY
I1RnalcsHoArKy7oalrh3fvKSwNQkSgPRH3nQNf0Uwi77OTP9qqOolz5eX9Rx8I/
fWahsyOlhziC2a+CADLQDWyLVucwcge/wyvtiH+oMa3fi1eMyGe5SowHyjPBWQTn
uo+UVdE3TWMArj5quya0smhsxfeETVbyx2tWxMiMfZAWM75T17CSdINWM281FeFK
RCXi7owkEhpo46A1FzlcWpkifWCCZicohJONySuZRWnMKHSaMeFc84PaFY0+tG0u
/8Po43lu6l6kz4USPpIs+IeZr+iGGpJxt3MBSUaSAJ7AiB3vI38KdWdRbvjHU3dN
pPb6bWr2zLfU1fJMK6+fgapx9U9Cac4PJgRm5esYuW95kUjo9iqd4dNsbKTd8Vuc
XJi79CQuMQIT0le9sc7JRSEDV6JaQ58rvr6QRTQw0SShRwk/fP+dDTj4xxl1v1Jm
q5g1H5bneO5yM7Q2476vwDarVyU1mOFhggfZhzclg5zPojmY5ni5ebDHuW6c13GM
+iP271uwUOp3oe/Hi7b/VwQwbtgRLiuwCGqU/W9pyr4ew+si7lt7l7JEr+gjA7dj
15extxtR4wHzsUr9IeEPPJ3iGE4oEzmyiIwa6dkAmpvNhJTyEmqcthuTVzeH0BY8
+bOYVXHcA+qLpX6nyrNcsOpGJpb0c6LbjmXg64YTFJrxUcuYc/GCSCGork64KamO
Tx6jKm2HkoL6oKBnX2XRDzz/TlK/vnL9q1bdNwb7pG2iUJgx28Ft+Z97xWYX9LEQ
i5kP1wQbBscbiMnB5BOQNFdF2ZYB2C1XV4TqU93oT6QT48Aq7KTSFo3oN+LkYVCN
53hJnDTjEVc/CORPy1ugwFtHZp98cwSKtBt406XqDZe6aHTUF9WOf5WlwaGLecsZ
qI/gUQT8eHs74powYO4VYj3r+Fe61pNSE6mEB/PaOi7h+LsLGcFaLmrEw4H3qzQ7
G1nJIdB9SI/ReBJLU35YUDz3C0iROGVcFxl/Ja+YL0Dhm/2WnfuXwibP/Q/lLbQa
ZfbgutgoDLzPA5pfKTI4jx+oZROphLs49IclC3tO2FlSP7I6hA8h4YWyDS9AWTv6
0i/0UEXm9b6FEQVgy/twOfNMUPGXuA1ABDGN5LmoNoLCk0TE6x74wPMyQty0ikzU
VuDJhqxiO+bmTyZrhUZ9Op/DaJ/bahhOdxyz5MC/2hJzaTXouJSDUSKNF4X86tgL
N4mP9YqAScjBOxkyhFDGfgo5LqaI/EEsvYRq99M2YtAGNgHOALWNRS7fmViivXno
5i4tFTO5W1qmnWsJ1/1mnVN8oZbwu/LWDeVmkonj1NfPdJ7CICuwsZK9cMnHYYt5
2BCX/bk7IlprIJi3ET0RGfSqbkElC6IlgwDBOrIc3lfKgHZBxBj4rU/UwIzz9fRQ
7NC+G6jh97aHlvZO13lt3ILMj98MkzeIpR5qHwUiahhU/qfuG2m9iR9BSbJmDvN1
+oCnAgs3uZD1aT8yNADfaZQUen2IaiKOj8Tv4GrNzfCpf3LRIB3ujXySCQ/ngRWu
5upPIoEOD6lnALGScrvwK0tVnwbZ7LVEDFI35q5X6q1mmO/yqbr2lEyw+xt97rqr
q8haqCvQetdVd8JXDHVTvNaqNAEDptNoGN20EWMVCmGj1ZNpP8z5QPpdUeYYm62M
4aTjAp7XWYN7AVh1wl+c1Q4GwloKs0iYsYMXkrEipyg5PpVUMqFt6843WdFnpF6S
tP/eEVaHYAFmLnnoLz0U/QmcLHlidAmZr46IflAPIRwF7spIorPnkRf4czlZbhxY
QnXSriuj7Fqv0JTztTM+Xm7PURaylJXxY56VfbU4MkvslWGtACxDWfq6Kh2Cuyqi
sPNCIV6DxDy0cMuHX98ypx7qMO+rMiSRHa3rlWoAfx33oWtZ+lGSkbaEWpD0Afkb
EsoLQjFEWJCzaOBqELe9cKjKXjOGQhkID4Lf8UPqpmQQav6ho4BWLtrPQMmrEVZ9
aDwLJT2eaSo9ofjLhTozjXyQ0ZSeqIw7BTL5M7sH3QgIZIYhsOAnoGfGX94YMJGH
M5b2uxza2MSInidhNW/BdMMTAgcS6s1SFRJlf8ZFaogMtvZF8SOvoj5+d0bLRBSe
qsVEBGpxvJJanWs/HE82Uw6ZwIWFoLADcAq1qyoU2/WdO4qfIf7bN3mDPKgxS15S
wFkTY9+5ChKPL6ouxHYfc6qsC6xsba2JDaOeBKMYOFeLi3rtZjOX31LXX9eJPCd6
1QTBXGKGSJ6mL+V8AG35xfLN476C4y3OVm/4F+TCgkYXJOfFaRs+gLuvK3ThSKPG
yrK7VihfpWhL2yrTrvAFeHdDK59c/3s5aUAEoD9LNVWFWPT7V1twyY9hQo5FVWwl
pk59AMgZjFD75s7IySxOxEgG2HbBdpPbTMun2UQW8T8q7ZLdTih6YvhI9WPcaUZV
g07Ullhf/Uc65U7StF8aC44cAMsaH+g9yHNPhCHfUgZdQdf5slPSE9B7YlpDjIXC
RFiAjleJv8yL1gMwVVGfne5Wu//mqcSvuXq8yizFLfxHTR6NrW/PfVvYiPvLrS2D
f2Zkco/p9zdNtveq7gjnJeZQUt9WkwRcGzf7LxWT/oAXaSpO1Od8t4LlYYYZB2Oo
wvq0pY01G7gCemOktj4cTPkZEduyPxFfAb3zAtZs2XCbK5qJs9qHQY7MiKcz38Rg
Dd0Fkn6t/vJ2LDUQpknNL1S64o+FyRhEQnJxp60DJPE/ErdE3pqKek6a56GnL6BN
0WYJxPqNoeAwU+GIB2WlbJuJUA5HJxBsMOMvnTUknfdhaMaUVIXfCsNFrz+W2I1B
taefpbFNw58wVzHhcMj6LoMkVJYrsP344FHk5qUl03MwKhxkf5dc2vBehr2zK1EC
hQhvUKQYlVLnMMX8aSpbEYiG6nEe1kDqd6ThGbTh7VRvhLwAnz7yjgqxp+edKV4W
lr0Rql4qhKKrMspYotnsnpDHak5lMp95GTDQBBRhHgeN/StZz9CdxK1s5cQOvg2u
wTfjnbOi+Qd5NOW2rLXhm3v6V8Oh3Ck409q5MGqTO7FnmWfS+MX9wRYoOuiHJLR9
t/CYh/YjvAdhztXtW21dr1pL2cgbKkjnZFTj7aHs9Xu+GmOAaNqu7kH97Y9IonEG
qZ63pCslPYJltKcO3R4uw12Zo/izir5p0p0OQfynBwEZXBkviJVkOTjdR0hiWFEv
k8G1aF5m21IEWmoMhFEpLnTLxQRn6G4qFDfqWRm82Hg6/IVFvTMwnQtumYEem9J+
tNT2Wj4aJR+5GG6fSjHJHsOKt21m4iEEAxLVXNUlFoez243jLdH+3YB+Wl4aoo73
N0tqWCy3tWyMw5trcK/47yA++poo7/faQx18EsyYcogHyLR++uwhDGQc/EYH54We
gHudM9RXqkN7Mv9zcDXiQljodooH2DDsfN2J7L7C/kBpX/QMnnQoAfgltZdNi9xE
kNMINrbON5VGYeB5L9eE/SbJRxzS6KPVGmDEcxn1j2eiRvnPhiHjx1rGTUYriKYB
BA5zB2ultV6oRx5KprFJx4c+QoL0+Kba32BcYdP/xitDWS2NUZlC7qS7eD62gbuF
6IL00WtjS+gLV9XN6sHpXZ2anvaqtJ6COJxYdV6WXVWrF6AtdpWbYtjD2k4Q8zFX
jqTP/HO82ipiz1dg3/2NQI7lmwcaBvQxZaeTjn4X5iBZZlJQ2AXRA8nkin7r5iji
vF/snkBOj3d45hWbeckLU45ragrjj2pLFLxWJr6vic9Wkkg7FedZDy8qTRWcls1L
biQIgVP26ri/RvhCJwnkLhkEVCIdS64Op0+QZyF2gK0LFQe2Kw+cPrNqYrFDM1o5
eR/Sos+0TfiHk6fuFZs1VfmKLrd0jlYB86Bt81tgmF1whGxz4I1eXcG78Xc0vDvg
fK0DpbjpBKb5MQqQHm7zmEshGnAUHwMEWBnNZLr8Gp56XullZbxpFgNhNgsZf96W
ytv7rCVSooEWT69iqRQeqLMY8o3fJphTL5cbBzMqy29v2E6Phm3wLICKrFh6FzIf
s2H79DPakjpHWYfzhP6Y27bl7lV6WL6IL6Te7t4CXYm9ArwtXI8GxmcyFyb9WOL2
h7SCOU4gAQNYxCltOMYIRgaJR8ZFLfXGDMAZfodYzoOtlyZuMbLQep1A4HwvSJhc
oYqRCrW08vrCmjU3+yq52qHFbQeIbk3ZY4fTf2qjYVSz2qaVkLJyIKXlqYzoSeLa
ZDhMpXH0VpOZrYjsImGUBznRxOPDKlXDGPJ36WGcUlx8XMa4PnJpJdYeozAyNCoK
2HWlSOK4rDL0IQK+g8IX64HXBWt+0gqZZH5BDGDwvgk/5JjZuDPZwzDQVvMsHPE3
6QG2CzAwtCdAtDjlcisjpp4OHW7Ej85AQBu7Lu6wee9hB3cVuFDTdOIegMtoZwcv
T+Pmggcaf68K1W9myzGx73GYeNskE/Dy7G1bqzXwzFNpl0IsjLNOZiLiA2MifvwB
OVOxTR/KokyTEtcNhFajz6BHqXLoXnzO+ONuKsLKFv1zFG3Jg0Hu9mjFBualp6Q2
EuSrkaFFjXtxk9n3uamS/zwuZtwwd6ljDMy3qH3kT+1JuXDUUQL329VMCYHXUVQz
D4bkIwBnTYFWfdjuLqpuAAGhCLkEFA36nz3qmfhXasVkmbBKktLDFLs7frAk6cWK
MkvPGqkJ5FG/5EqMrt1wmQ6THjiMCX6r1s89rvxVQ3jX3Nv7mT08UzYPdmwKXHTh
VoV25U45trahzAgmTvLwL7h6Wa6zg6G6WpQ+mG57zJxq0X0LCFlJLzwu0bgtEeIc
jU18/g0UaoC/HsrKTlvlvsSBvNUNmqC3ZaXLj9aBxncsLKnJ2XpgfikObrfrh9Fk
tAA8zNUQ2WsKupKTrSTt6x419OFtsrcMXTKxUtm4lJIbZ5jUORB23yRtEUK+GCDN
ND6tM+FAoR9FuX0+QVlyrSoue5gv3se1Amn3t8V1UlAQmv8A0qF7ukXRpSqwNdT+
xoZv0sWmzBxcG2fUUbQqGxRimrNKg49YhOSy/bACZoSLTIUhcb9oDpAwqSRcv+cF
VTDjbV7BnuWqiq79uMvHrQTnng+fG5BqF+fym5ulXINl4SlnzXb98sV59easefJq
KBrJMR3Yl2I4LT0V2plSbyRUYkaHnGghuGG8lKosGEhEIFfUWKdaUlZNFLJBgb7C
vAAhOJEiEvIIB7zbLre/rSCynqqSJgm1vpQmRfZg2S54iTTQ7PYdE7klBXw+wWNN
FjCYfSaSOMOs/kNKWNBC2w4Tb2B0VDRfOyaZmmAXn0g06H2sPfpjkExUMdD/NLFG
hZw6iByoJZXBBYr/Keiivn5lx9V6H8kQohIUaamcKDaGdYC2Ghue8cH2DcEAvYc/
wU8yIP9QCm9dJKKxIUI2MhnJVTImQKPaJgr/t9jPzbiH+RwBAbQ1gpx0qXoXVdaU
hzhFf8vq4N3SgAmbNKMfKD9THrUBfaI/ZB9Cj8xOeHjird9zMgh/fbZJKcyh8mnp
xtLMishOcvtcRwQpmNcjAiuzdFDoa5nDJKgl81U5spJKK9fEzu00TywdAHT5cDLk
PHwcI5aQImhj7U4nmO4S/7+xZf3KFkRnl9/fajPMC6i8mOtWJepPKTWlf1o6ype3
MWS2mXcjaGLn9o0HXnywg2bgqBmyNnflH4qD79k5uN0+Nhj8IdTKoSwE/YDES9Hy
/mvvejDXah/qR6FhvNzjOsgbejew+fG5YCQdoUD0wkBzN5PXcm8VmMMDkcbtPsW+
WyVvnrX4mBNoY/g+6PvChIw0QV0erie+N/XtsM07OXITDFYqrs83Iz3iK2so2QQa
Axmuah/g70lO4WpaCQhKGimBjfRBZSLuED12hqUeXPF/yUutsrq6ZoVKgcVJrfu0
e4yAneuBRC5SP8o6ZujUpsuVPDqN/nJcM2E84AdXSTsrqeHcYAtl1QVI3X3fBGwq
9QUFaK11VAjwrArtuC+SsJX3ovfA2f4fBhIC829V3/z774bA2+OGHi1LcCQetWvY
XBi7ACdNorfAYmlnMxPJxtb16bqk7GHqvG7qXs1zSKh1t6lPst7pxkhZIFydkcoy
LcHxJPxPfNy002NqJ7kqyFhbMqvKXPcmqOGzM6HgUdL7se+gWre38sFPyw4YiGo3
pnUMV8XCwOZtQhDpKa0qnKiPtytDLZ6QxSAmsaK/gbwZPn1o+/lhdT17apUfYUXl
07X/GPADvln6Vksciq6hkvDWOLZTGRAvaG37K347d1i9FgLRwIBnFulsqiz4sF1D
WozMzenZFQR32RtigJJHGu/+XAIiRI7yAM/W9F5aFa8khdxL/prRZh8/ZYbo/AT5
aRxafV42a7TKXZFBPndsfTAJVNTZrVS9BlbM/NkIpRG/LW9yEkzUxSI+agerLjNV
ZV50I9j4w3+XHQfNpKpiL5OqA2AHudneLMMcvAKnRLntJdUWkyTl5gq/z7cwhh+G
Uk3IuvnAlDLvHZ9I7fpqqZ7eoUAnExVIZtB+05i08MsOKTvCdZDARhsxrruT/kJa
l6dxFdSSiOc8djf0OQfBrGZjjnBBYzDitD6rHSps7J10LSYd7ysoQbYT+yAT5Ktp
PBplU2WEvJLuWx479190OwXAkTyu97zQ50pQAPWUj519Epuzxv69wvlHdBGkE5hQ
1bL7Mx+vPs2ipodsR0J+DNHHL/hePbBnGjlPfM6UUmpbOOGbz09Su+AuMRIm2Icf
U1cqFKQEcfEYiHYQQ83TnyozfRxDhgNx0KZEmMSJ5YETVnRxNi0pKleLGISI6r1s
hV1U16wharf3QJGxUCaPlf971aaN4mvZt0TdmLFl1+Lsq1MXjMvI3kxvlbgV5x0C
H/aMfg52Cu75HHI7zlHjYLwE+xYwS2arlSDoc48jNeHuKUH6WM62OHfk86oW8KVL
3K/3xYPGThO8lpuCQ5DBsqkUWFPY1PAM5Hc3d/LlnfPT8uZvOO1FCabUDJvWHsjH
+xBTWqqHgvgGGeMfhcT7iUV1Vb+HagNXBIl9TAXBZSAfSacO+kifL7P9WPiAhX2q
EvE30RTjVEQlaqinpcj4NoitiM3vkyvtZGyr3fPvyoqXn9SgOM7qpDuW/3cv7tvR
oN7KBEwBFxIXDumRAanm80kwMF1tZnvlxbtEp+RFfu2WIUxBFIs92PnIt+hsrQSF
ogFKrBoNdRGhwm+UQIpKAC8+lUorBxGqmtOZL8jLUSZxfmhScBhaaM7yJHwUFY9k
qJdrdSZ62VmClr73Pfup/AOb4J953E2TqLdCr70BHT2tWCUeyAphptC/nRwqgKrD
A4Y3WrhiLugyZLyITXjbgUR8OYNpeE5huI0/BOf/T4p/T7UoXoZhHTMKBh7wE5YM
VjDbYjksa6CeTYS4L/KZbN5qfzXP+3yol6CRahPWq+CFI2aUrXriaILWuiEBkos6
DEv/ZzDngrhHloxh1tsdGpqd8YdMIG2KMXPg1Fbi5lS6FO48cuJ4azCwFcaWOKtM
aXLyvtzBON7/6qejdIzeZOWiQVj40PgW9cVGH9M5GjFOgp+nUrM7vCYfWt76ezRH
PpnVMpWtlNNWFzK6hfwPEhEE2oVaGqnlVNcaT99U1hVdUfClkVxDw1tDYBliYdjU
TBws0Skv+Cty+pgOc2jFX+3z9un/M7GeDBM+BhCM/bj4uJqMGBMnk1csTrmu93ct
jlqmQUsnHgETWv88eQvS2yX38MJ3ook6MRr6h4YE4EnTOGj0p7R3tB6X95ii86sx
GtmjYtl/YdBMaWRN4P/bNgqEyJWqmVOYmMeyfDmmry1/NAC9eOoK8FEsnDT6vbda
YiqftoeHrZhrksoj28VXdk1+bQ7XuyYlwnASE1hkqimMQHUJkokmhnvNaLKBFB5L
0yPAmL5CV3OY95TT8sRVu8l9FgPHbCzRXSrAgjz1rnG3NNC82t4gYHvyBtUrtqxn
mRtYjNYvgPo6tyYhWnlr2ghBES3rdClUAIs3elajX20ZL3CAG/fcjjmJYCEukGAV
EsTSdwvLfTmS0xLOZkCekabFieNeO6K6tnQYuZtBUbBwILfHNlEhrF/K6XsP1EQO
n6+f9wuC5B3+81bXkIlyfpMFY9LnL1/vXQhHi5xLgUlM5134jRRfQTOEARLzxyXU
Gye0ySpvZjVfgUROzhZlI9gxoOEibIcIsUv7+vC7ZkQZ1XZUr9x2xjSLS3UhqTKM
cDlZ0+PigLFDD2qU+qz74LU3A4fwBLTAxLmdjRIkcEkk2AT17PvU6Xtj1Y3zTAz/
FoCfvAm4VNHUOQ/Ew2LcA2+dZJbBCUIhcKnJABbMw2Yq1WO+26QaxhJZC4dFM2Fj
Qqw9qZmKot8PPvqfs5pGZqKxDYyUqMImhjkOLGIFQt3XDFwXl/oDtC2SG9BlhuM8
MP5Lg2L1xpsmsKGtsMuZRh1NNT7zyebIk1q+7BkB5DVFnBRD1OES4iQhbgOUQYrd
TzT1pmTcHIB5yfJHKEzmgrWajYILILgKzS2brywwqKz46ld8ixxK1sVhWn87G8/V
PatIudA6bbr1QYdaj82GxtYnsVwNp31wQxcRJ7tsipJrNIJwx0cNCe0C37+z9/kH
kBQf1nh09noQRS66JK8xJEpimGGBMeuc+ytLvn6H8YKMbSdzwBDOj5PjJdbkyas8
mwRASJl5LB5Jm0zcyC4D+6QMnU+/zg6Z20JJWaApddij4s7aiFNoiPvg1B2Tu/lA
YoXKZx5hhrw1qAX4NutqhGUk1l/LsPyplIL9/38hzXqMo6Hz6Wq6sVKYuy3Dyx7q
+NdOPuTUY5FeJkQQp6cN3WQV4ZOX8kcH6si0W1q72LUCeH3eyqpnP88w/uWP1pUI
eDTSru5dL3Ww5p9Zg/wgs7dvjtx+EYUH9FFWe966xVsyDUXf8b17bcVDIRwJYWIj
o4eYpRs1Fh91iH1QKJRs9LN7I2zN/RP4RA6P40OpGG08il4UP32G6xQj87PHGVBB
jBXyP1UJfi2kWvxnxxFyJnPfrY3tM6H8qp4HjFyrEH48zCN9PTormfJtCy6RKOXn
X8Jd0OovQndsE6cOzfrJNYBwaS8l+rXvcyhPIEg1stGItOO+PGfVaahGZwL8Q+49
OfVVzzymVQ7WpG1tXbRBzJf3GlrBBSoeAslvSEOHbbKZ/HqhV7iM8lfv3rIYYWGP
8pHTY2Lz2PhKlrp4n5Y5TJ6d1WYabsnTkeUiP/z2Ui/G9Ck7rhr5ojgpR0bowMox
5wAvH/sbXMDeeQRc0kGKJ+Nw3akYaMOfmAHs7wAJBE6OULlfvb3Qf6a/wqdwE2jj
sfE6woQxqkl/o883hp9DsgTWEsEA/MtS9aaJIY2UxzN3ORvD0f6qnHN7OXYDoQMG
I6F02rR6zxRbST85ooLtdA93+i7C1tkz3uGBbTkqDPvdQ7bNBJQ44rNB3RbcIgRC
ebsk3SMpmUWUU/7Suin69e62BzH3afoSJwwzn3/MHShwH/vux4Ro11iZWLOECAkD
48e8bLpOnjyw8eBrgQ04rhaqf6UQHvt9eJwMUgqhMMh0Q6Ny0kC8+WjUc4D1ATRD
Tt3fzL10FC/M5jWQ4JdW+70dYrqFY2eUycYVCTvor0QzluHLVrIL9yPudnx75qDg
7ktDxEJegCC4bFf0J9BYcAIMQutB0gxN+4q+u7LoQwIPO3GUt3EQ222gTcDUi0CH
sP8xEpEvEqiRpGraky2QIrpuoWujNW+mjk/EwRs71bPeILM1NhRclR+jOfrKfPN8
bYovnq3X6KTHWzZgfSgjyDY8f/tKKhuemi/M7PLJ3QYaetB/1lR5Inb4/xtGcNYb
v6/fJqo+NVjCv0Gq4Br+G8RuYbIvfPCCntY1DuLD9N8MtGYqiyycT1Y6kHVKlOvr
KNbFB60jDggDoC/7SNVzKY027GRAJS+4yD9KYe0PuD/j4H6lpF7qfn1KRqmchU+b
6eqbFneiMuSF+Ub25RTOT7CR6aZS+JOW5OJODto7aG4sQ1CaCmljbnJqhVDhqT/U
FIKkSJ1SMMMVS/QkFKTERkJayQsTWSSM9C0z/9Gm4d1YCPXDyfzSkCBk496UJoL7
gp9ZIjXzKeVuAc6kKUuxRCmS1QSuOOwABObJhKsrm8H9lnVf883MRjk61g33iHLU
U7Cmv3BqbGDmfpPDmsgmlrQy6/61J+eEzPTDazEknZDMBuX/nbdFRAoo95341FSQ
WJ9OvnFpjQpJDjGFUni9Ah7qCSom8RzqHd4jAANgFX8Uc2KamleLnNUH4Fi8YwNC
sqmHzHwOjJdbTvr1cLAVLHNi068puMATKQd+MKGu+Wn384M2qHs6252RN/G5jtV3
bYAr6Sd8hfqvcsj26wa+0guoyADa7ojh8svJm861sNa7j+U+oI0vJUfOq9Q4Zjvr
lXBUkOvo6gPbj9jVrlVQPiqk1ECO9qzFgCLRNyuC1EsFXvDinO8NNEYCLFr5oZMN
ZUf9ydqZ7817pCLiEmp5uIy5YajIDPE5/CS0kzll2hAHPqtzQqW8LzjDI9y0EwOA
XqmP3kxiqCQZQ1HXRrCM1uSSKafJPWOS9uUUqxzJ497pmcuE3UcvLmMHuRaXfgZg
t9ZL6zNshUbPTFpO8R6esO9VMg7uL0txo3P9FQDHrIxac8BFv6Zhz+318IhA4FVI
kAOzNNBMM7J3w9IkVx4JuyZQZnjJvO/oM0tXJJX/ZuLK/iW+CN38VLSAnk8mtGFU
C7gjMs1lXRMns3WffH3v48VhqwlMaMO6RGuOJ1FJhmwgYxcBtfNK/Hj8NU7ooiU4
wjugRBLwhXoiWqNZssf0fox7cuKNEyvZlGmExMfwMiLXpCovx8o4VvCf60TUlAux
QWwuJrN23BSf2FLf4txgCJGUyJxvfVx23VgEHGpDK3/r/0TXMfX2Xi10GhtWSJ2B
SLNJsUSv54ymx8LpZfBRDZNv6XNTwLRNTvOi7Kip6ExKmv8JMzbiYX0cN2tHYhUa
CUvIDvwlvBhkhqiq3y6CmuWJ126Q/pEYlclB0qWHUrhRpXzp/d+Yf/2Upnj1EH8F
KzeTZkQmzjXEHIK1phTjHrNppFGAV4lTSLf6FLsDcXxQZkwK26Zdy02j2vxwT8Z3
ND+XCYWCXA0HkekRUSKh1GOtBODfHw1sAg+Z+rY71a88u4OEUGLXHuxPRdq0nOr7
TV+uYGPn/r/EsH5oXMj3grnhxf7cY5H6YkCzfqHpjuVJ8NtYMpwtg37lnUo1XF82
ZtqdKyryPVoAh5z9y4KT0PY6E1d+NUvQsOYIGdfA2eExyV6ZoP1JqN1pH2oryVBA
sfd2Ma001jRJ268kk2F12ImQqxXmwnfg+UXmJoSKEFti4idE5u0pToD5/dcAAx8Y
FLEGBPsf9CsYr4+BkqR+wW5dk+aVyYVmupQigflXq0l8Ir8bOkqWuqpeu/j2gf4C
UP/MKRJAZyAe5mkal/hviAKFbNoxfULFBIpRvlrRmFzSYwh36w0gCHTuB0aUFFri
e2hDQpYO1QydPU0aG0hV1pQH/9U8UWtX2XiHtg8AKEhrSLnztCgEfQfzenCxiNI8
SJE7HAY4SpNR3taCfmwLTBR5ofP6CRk7D4rWuIXqZP5BjrD5T+EOU0ODH+wmPto9
2hqmM4I4WT0sspZp5dngjZ4WHkz6Y0czT97/5xPISzNav+2CPkMmplgShmEqDmEE
nKr4IHu7/aPzoN7dc7vS08d9480lH34VRBygo7z6HpFvuX4wG/ndfmgl2QBqer2r
HpCOHtsFQaHUHaho2u1trlYRtWeP9Tk4ZGq4lUdKEAZFvYM/S/QnBd9y6nrL2yDZ
WnDelYME8JvlGve/L3viGxmMI0YKovjHk98IrFBmjRlsQKwD1r/lggktdTOmP+Fs
zzRsR/ev0uQJRO/zaQwaqbl+704eyyd5pZq0q8mfgKGNIo4Rxx9gJAHkUxsg7gp/
g/xBeoSLsnsvqvhROcsDkp1v0mCBBQU+aDIGJIoc/7pgfW1krq1YlkYXzAwF1Riv
PGr5nwqYUXjENmqTdINLgmevpePtXdUz/wJ3Bn9Db8/c1XDI3ORcXneaBfRhH4zV
7lUqPtPMh89X9MB5FnXdjvhwnz2KFYoZWcPOOvvlU5EtGbKPzGr0sY18Z89RI5CQ
pPnEgQhUW5FM+RYxCQSZDLSbqwIEo1BTPwMWNAl6H0jm1lHG8CdVcbsp+r1u7nU+
UlMn9dxMQwb3ScyLGawDZAPn+VzH3Gs1ltL/2pQoE9yPb8facsWHbsMkaqkgXnL3
JDeBqya+arqyk+hJtFrm+w4BqzVDJZZcL67GbI0B3tYTQnikiU0Tq/zuPNFxB81x
anheKyuUJI2b+RL7V8D4U3ufRpt3hzuL17O8gQiYqwlfjsgBJ5Z3RFisQomrN8w+
rX6er1weqPSwkrdSkRIVrKqJsWdLl9Px+2uaB2tseZ1+gsgnBCNdRadd7XdML/z1
fQnm60VQzE8oh2LzSfDzm7ojzCgLpfLTd9FplxmD2q9R4xjbSIndgJDs3Wt8ld99
IuehOymOnTFzmFVjSpibU37PcXT1iASbNee8DVbgkQJnw+ugpPWdfarDTPGhJ0t4
u+2gPC8MVKHpaQ7yG29KMyDu2aZ8EkS1IVc2t/Hid+9cOOxMV8fuMybcLKO7zcdn
idLc3RRqfcdppiW2yOADDPGKaJflxc/PnL+X6n/GgD2+iufrqjCK9CE269i50mfE
vVSm5INMtWq0H5h6qcBRlrfY8Fn9dQDDIPB+WdEEvVAIMvPEMzErQKfxC8zN7OYb
0UcCzAmUBi5+tGy3Xm5bpMLf1Y2Eun+P1ddzpn5JjjqhDwjnR9/1qK92oEARZ0cr
Tm54m29Vhon2oYSyvzJ2ney8dbABSCnvYDfod54Xjqmh6HAMpLj7iJ93726iVp5z
DnhzIqtneMyI3IYcOnw9QeH6J91jRQ6f8j3gQ/Sc6G0RQ1Po/To1Bx6gA31ajJmg
VMtJYVQpw9N5jRf8C7JW/jaYjATvdhTZCxPuZP16cxjZMsiGCCMOsId5JQYC0oMT
FQq1rUfSvE/HV+n7mBjwbStyvRaOKJQlZ5wqU0LPr4RNcX8x9CxpozkgGv0FxTBU
GEVtCd8jsCHfWW1TN035sN55c67S/xuBXf6gepBaH3upeLcrcd/f62wthJLA1O9N
h5qDH4bhOz/ws6jU+nW6EYBZFLQlCnMof0FZaa2+YyN+iAzWcqbpq2OYBnV4so1o
qSbnYUg9nJ7/8RxqqKE1r1zTvDNqZXu12G6hXkObv4yefKtxv3hXx7TaDCVDi38w
ZDlCZyEJnLZFZtMXgITJ69w/YWSUjCokjfFprBfYU7aSs4lpmd+6cmdd6Q6MPMWX
aOivSrVuGQ5UPHTPeYhn1sPqRciwXqO62sFpPwwPh7XbTFydHiuPEgqPLzisnIbL
RNtHFd7Ojq4q2+vLeFVfFdyHyxfGeI8TuEPqStCul5+r9/qt/l+e0UkNlDybLWs3
ExyTuXew22CzfXdal3ZmGV3Xc8Dh3m6TTpSz70dFKwt0KvmjNgGhVU8ZrsIXkC4i
NvNL+Wnki0fqPiNq0ARPj2pDC9BWGpIXUX1e8x+z4yU+r6vhgNmwNgmUWtzITYui
84RqDhSqoCTwsmDTkPCzJgj5Z/iXLICzJqHcZeC7AqjhsZ31Zz20pXpn//gseRCi
u+j6mFIMs2VMz+1PZGVVTsm6Ch47GilJYRRW2dHMT2jaZgPLU1J58EsCukvQvcnX
ieD91XQTC19uVnaHsKRVVP74a58roJMlDpyf4WJTskvewXNOEP68lMdZ1mRO9cl8
VzWuiVh/jDZHd4DBUOCwqzSwIRNQOeFvPXZ+CZVMMLMu6oIVZHq7YLxI3/WFNtwB
VF3ZumPjk1J5P9mldj3NNOXk7efD0L00fzs7iUaO249At/znhSB0+LYC2XmSWqNx
NJ06tnbObeF4ImoatZ35OEtLg77wQfxqI/cz4kY5Ew8LUHHi2qGgVure8JCGPAe5
xDSpzfd1zYMOXfU72nhRQxKyxbkIG4zpYLmwr5XvzLDc0oazBjsqKmDViTnIbqqM
Wy4nH/8wLFWtV5l4PrDu5c3zuo1qts9lLCjr3F5NEdmtv7VbYI0iY3WoAYETXA18
FzbSYlm8vXQF6iw/KZJDOZUvu1ULvjvPU1uRt5Us9hMerjxwIwoTzuekAJ3ZE+zQ
6crVjhqnY4uFeoc7ofKKF+ioLY+FzpaVOe28zpDdCLZnJ/2bFYG6MqLzdzFSPbTz
6qvShzN7468HoeACoj4VnTEEJrFijhMc3PZNSE2m25J2lxl/jD0B2fGYM2vAlSJf
mDTQ+47WA0e3oBiVeQkgAK6Ktp56zDEOTcGRsPTVknKpwctplBknRJuEx824dGno
e6RvYxh5uE/3tW8X+3jkycHRgI3YGII2cZtH+TTBLbVpRq8v/JwCPSTVQxXv04g/
U4oDFTpINx/UfB7qOY20sDsALRMoPgppA86T47S1p5D6N5tl3PdJeidjFd+4GDzB
K/03J1FLFF2taF1SEMkDO+iyf5ZT4Hih5ePNl/UHVsLPWNS5knlkcm0iXy1ZVcof
5L5MZWNLrn9He2tBrZy1mnUiA71oa8cVDXCq0O31IZg9T0Qs4h5HmEToNSo2nj2N
YVOFJ79uQsV40qcPjzfwLZEd5qIbyaw6EaTAY0SNGuP4hlqV9GgS63eIdtXQL+oE
jvihnJ3Zv2KeDQbosxod/0wrRsMicU1rsRMV3UoCONB4wGfPFrBfop9S4zzUA0NN
54z9CEq5vv2VxKxALxHSHQjR4AoOYn/2xivtg2HXOQhM1Z++ZM8p6Z6P2XrRCDWY
RjL0JD2PJnXzeDAgJlH7ldZv5REpASyhjg96W52w9x029I3Ve8+mLdYfGSpqHGuX
B2QBugkra+9pHHfRpUxX7c94HOnCGzhRikMeLFF1O5f1NItClqgGqDZpOgEWz75w
F7XYz5BibBvmAs2Pjl6wo2J8zUtoXbY+FO9NVni8OHZywCYyncNHAyQJyACnPT/Y
Gct5+YfWB4F1TYvYA07RqTwyHHj78nKg5rLDEymjxxl3ZopP+P8bM5Z7FmVYiV1O
dTmMDCJAL2N44C23iOqbWSS+uiAuPKOnC0qzyKEmgmU5VQneztjGIzstsn1hNubE
D+ZWFpD4nq3jT2kF4krgz6cUea3zNjyoHb7TuJ4pI4fWnuiNjqLV11WbjYOD6cH3
cXG48oHw+b5HvpPNY8Yf8SHEKCB3j4gD/MhG7Q0H6YUAQINYsXpfjp0/0yW05t9m
XdzWaFV0VgRAN6S//o/Rv2PcMdvK9C5xcwdlqmZI03g2F5dX1hyQuDLr1LfYWdWg
H/G33j+/8tmh7y3Z+zOfhOZzW9JLXtgaIvW2ck7zvCw7ehOhhMWpIFp7qV0wX4jH
VxxKvZCE9Oi/d2iZT4l0IsYbfn5X9Sa8MBJGY6FdAno75q8bStKksNuKYUQDwBxx
X31U6d6d6OiwVjhqv1NbnEKx71HEXfShJcdxD1VaSOtOdVLX3XqgD8mfenLr86Xy
t7EUEZXMT2ZpkgjWCQTlobiV0D6Wvew9xXfR1+4iEXdb5nQy/+sym1NbixvxjNkM
cY0agWa+lFg5DCsucbniISRQ+YXuwjYWHzeHY32Fgp1wciA35+SNAH4kOC7rETal
I2thPmWpntHSMBavUoeimyim4IHhp/YooDCLnUr9xibOSulqyG0hqU6eAUcvj2Z/
cgFiVaRUOk9Uxg2blOH2J3eeo0fNnS0G48rnfKjOeXxEU/2czIhStT8HgYwxUZOc
jYboZ+y+lNp5ZDPe7rwcPrgL1Y2j/M6wxFfPJPE0xIyE2V20VLBDXAmFXo2CGRwt
wQYMPkViNSpMf6nOW7px894XOOwkJ3aeu2L1wNtwEAhj5ZXTpWwPgNdHibRrig4I
QFG/5IEDUF1BjRmuHElENceaoww+puRtqytDZv6h+Hk7Xx8gjyeL8W4LfAm0JMs+
srM20/oJxmJySzo7ee7DIDQGb5TglrXzrbr8XqxlkWSYFjMGAWOMqKIaSBOlBQWs
Bp9Vt2xUGLbgwjAixP0qaxSxPrlIcTNVW8bVlQ2DyCExRBnXNdvGqNis9IUkqPD/
p/HfGP7eK2SQM6EcnqWUJDG0P7utxM/ESEjBf81dtawL9no6b4K8IXEaBYRJGApl
IYxUNxPM2ga0BlFlnDZ3rpVRkuClGToDGW9f3CBN8UDePBq0Th12wj7YwEwlCD+Z
Qc/g3sMjLUmDFklCfrZrl+HdHnbZP+byzm+jxWvJN1M4ws6NIGMF+BZh9/HaGItS
0BOL30cV/JAZQDQI+lEdWIhYiW9r21qK+a7CCtcMnNVCSI4bfjRzic5hlEMYOhud
xr8A53O1OMiDtqjInFq197LbWrm8vs/N3OgLmrx316zMQOyupimufFLvpHGVza3b
XnS+t4/g3SJEKwbIr+9GXT1xB3S6vrJok4AiYXmmp7EnHSxYaBCJcckFQt1OB0Jp
cL8ZeV84UIv0OkEqWNNDzW7YaYoui/4FTrfibmy24/zSCLWmGmfhTAzSjHSPTpTP
5ZnrIFZgb+ONV/KXlxWTtHxnM3WgEaTmNPH9KAK0RyJPG8TgiCMnrgN+UtU1jA9/
yZsIWHgq2TUx1isjOPgPR1HFYrABsxc8FVvkgVREdTLdFTWEHFpQmOY1GAIEBnOV
iTzmhDEhQEruLdF9ZEDzGbCdvDjDWtISX2kiaaZAIUTDiSVfdP8JWMAkJ4i+TxXK
RxMFSwI4UH6/BRODSpjoePwDA9nc8Q+hzKvduy1z0zUdxyAZjbKQQ7UhGLI41rtp
FadEuZg+0lNScHdIn0UD391xojJ867jNXMfwGFMHrLj0C7Kid0bVSRyXRIuo8hvy
fb2YRzNADsEudo2c5vyGPC71Ure9PIGzbSdfZ88mRGfhD/KybG6ZTC7/tKVIFFgz
+AfyK9ibkgzC0haqvmYW30OVRbRs7eoemA/m4XhLxLRxXEG/rSKlMUFiVSfyPpat
XkGdiYWaxbi2xJkO5h5VkidoDX0K41di0nP9Dxt9bhvV2CccgrafwCbjMA3NZoVp
vnLIhTPm2AXEHAGDjgrUsAktkC+LCis3FmqklfLm6ML2XpB2506fC3qvDPD9F8l4
gJ2PJvuBq7rLn7bByjR1txMGf5AfsVD4oPcYufHI/LHMsJHvVSEp/RGMMeXNEWX3
oHNe0IvjhE6KIH+FqaMaVvnEMh3VYR2JKywfs/cTe3be2Xplwx/Wgkf/GBIapOhj
CNDmLIf2s3EMuZBrI1uBrVeluZzJv3Nc0uehb/wVvJugGB9VePZn8J0YGN//d0Qp
ZmoogB4Tggyo0XKM2H8RH5As1IBePScpWzRN6JFRlcNPzvAyxpltVVljLIYhkCBs
djtTOfx7hCyMvvoN3nDJs+PQ5vFVZq7YzXhtBtlVIKDHWPm3luohJweMjcltJjqm
ud/e4L4d9MKVRoCfLFo12kP7ImjaefXv22bLGDhtoQekonz3+wcAK4sMGxTikNaj
Ecikzq1rq80DLiNabocrE/J/y8gwYLVurKVwwKlT6UOUk8JkXmY4CMneJUsk3UPk
Dw9k7Hka4MdKWz8LojtheT1YyJQldt2/WLJnhvW9nrrfeS/alIGxwvX85v/1LqX9
bps8ssd8DaanA7GgiJk71g/D2GGDvxTXa3o6OPlsfM8ix4B0yHGOtcoGwEp8qxhq
hEnkKrUbecR38wY/62jhQQhhBveLXhkzVip2wx23AW1T5px4ifbKTxO1oHkUvLKj
HSypj42SuR4lWS8OCvlttkBnCQxujNIMF3thiyVDRQksDT80tifP/l//IDVi8Z54
QxJIhV/Gy02Gqvh2tH0EM1DaSgA5fIKq+LAb+DBaKaLhf/JIRr2Ealv7f1oUlWEq
38gG5JTnnnf0NECAlFhX6vv+MwEM6trnoJI1obGVqqT7+R+3Vq2lEFd7or1x01av
L6L/MQl5oaZSBOM8j59yfv3ItSmHr7FnFQYPwWU+e6VfEY31ZgzC1DBGtjzpPxHN
svoV3x5jsG0sLO8z5FH95QV6w11LP6J9FdgaQM7KhZ29Dr2nsyIgACAc2QuJ/97s
fcqL8ab2HGAfRKYuEADut9Pc2wIF+ZW6ld0dIVu2rMetETRZ5Nh8u9fYIs0Xwd5e
HwqZ6rCcad3OkAWPXZOy0F16cQxRYiAnfn2cTTplZnV5O/m0Zlr4LeaNZZ6o7Vot
1I9aEjwJ8cBUDI7aBO3vjFvfu/rOj17uPcyVIvlz1P/nkTy9jNCjmHTbydDnvVG3
nXvwiQDEGtuMv8y//GPFdF+bnpfA0+bTi4XEtuwIstgrfdzbwiiyQJVP2KgWuDf6
8f+DqJVavMLanLe0182PPcqgm3fO4QhmmRYlIp0hk7EjTm80rgfUT0r2eCXGV9h8
KxbLI2RyqE+OEEeN5+sk/ve/wfqHV4LHimYvi00Dys1RlGBsRfYS8YHG+fj0G9GS
BTXb0IygWOXONmUngWm6NH1W1P9giLfWM+34KmvYOjaanHHvyhSSHkwHh2WnJgNP
D7LoU1KoPmsY68Q5oeJCUFWxIxcJHi1nj3j+7jcnVadfGVWkVQ8BzxR8H33u2vrl
bHcKn0EmE5WaiwEMuXJnxdy+TgLECnXUhMwiKlE0Tfrj9fNdwqtdJFkPgQJMHtt6
nkL62a0BcdTGNd45J6zAReBvCUNbKetUzDICHYVe8bGm3hb7ixIGj4dxRIdfmz0A
63FNZkrhNF8NYLTkNeESXMakxgQEzQBgMgwrkfRa7ka8IIVWcNl58s6SlJ3cqbAy
TIqHjMZJaCwZqF3ixmAfn6pDipEVAs72FKvJ+n4Ozhycmsu6rRT90kzvW+HDBzT+
W+DwqwCQ0/vheMe5swELsENkkfX1P3oxTGRmdGDDQrQBFQTpA346ByrkAP+S2yKr
qChJpUE4NGeS8s5rXRvofYoZh/lkTOx0R9BN8xZMFTITGQBVHl/Pe5GIg4WHOigR
fkRzxP3s+0L8fLaU/k9BlBncVUFi+f+H2ajDu73KG2OhSHxyaXPT8Jm1yicEzF58
oDYzsPxLqjCL1GuIQK02a/+JOhnwqbYEfALYHsCu6WXQotF7wq5x0avoAkCobB7c
c7ObaGp9MeUo6/dkbnsXUwL8RhNEQVEZeliI8J62xzc5qNg/ajpfJujekjBxdgid
DNrhbWi5wqqSXJ/jqnTwx291Y/uhWwZhL03pKNd9ZbG9YIL8CKe18eVnHn/a23Ya
FgVlYB5Ft2KotvByzbaeScEqR3QBn9wWd9e4DM5D5YY9u9A/Lpa5aIC0cBTfVuxn
2gaU26atA/CL8bHq8Uz+PRpjwi0I/UTsU60C0jhEKcI/P9fn4OQZspzCKbTVmr9h
4itnZhK/QvMMBYUB+YXjJcO4d4cpIYGOi4DRIUa69VdJhOtEDVWYCLx6KwtBGxuV
Qn050kECxqRjHRaHz5sec3YMWql1Z3upkKpPywUhzeEn5B+mwJq44FCn7eRghSEE
PXduORmYgXx5B8WBwoMerKo+sw2SD5t6ezdxaQPrgoMXzLFNvRdGLTH4om7kUcO7
8EMq6YbdeTCV3Pf/YPJtrzZ9omvH6z4xCW0WXKo2dr7qXx+AZNTjAaGucoD31K0W
FqYv7wgG7o0/D6LjzysWjUMgtl8qFooZyVwL7ZNOKLaolIkWoJDEglL0wQQTAASO
oK5KbB0Upwrp6EVN/YpT/dxeZE8smMseNdKIKPZKoxq9/W1kevTijuVzRKgTQZmB
Td3popXV8kjWpr5Yw7YOeEoPt3YWp+34iubA0lxY0rLWO9XWBgtcPxtdZLqeH7bJ
+SdekfvMHKyKNhNsytgYXaBSgAubw1hMxxhpJLxe2VHIJSVsB9qI33umud5MH7O9
iA5L0qdf5HiUCpc6x5MPaCMsGs9x7a6vvvXh2aIjZ3qEHpXoaX7IXEGqjqorlnN6
yx4tpiFI3XcZXvMEKLPY7Q8emm9zBQaXI/etU6e8SNM6afHB6Vcath9ONKZ4XLas
VjnKBxzV/3gN1HqXs0lYqTJXWJjqfYnqoHqam39vPlMowk1VxgLHHM0bGRlqXK/S
af3s/WiY3RXQX8iLJc1oVMumNREZmSgGe/t3RAGUgD228UnWoWfbOwr6peYjTe7A
RW7OsB6z9q405StFGMRg2XySzpOonOfIcWpBcG9F19ERwkWP0mvV+qDN8wLUTsFM
sI8CG42MF7AdEJhcV+BDbvPErk9Mqz4wtmqyyYCkfyfRZ91DMdPHBnbm/TcMz/K8
jnVw70Ybm/OzCFxNI3sGUzxl5/mWTimoH7FcjK1MfGP5qV07J9C6t3joFyUwjVI8
lziznl+T5RChFa+Tx8ku/Jaxv9irl/NEn4W5vrdnXRXtD7GXNbPbPhb4IyVeI9MV
WrEZUXk8yV7+jQfNpwMqmw5/7uTTI+ikCdxanxDSVg0BUV2nqdmMltvZ3DOpPi8n
Thz6gfkTqO+A7lYvAeiZ6PsPxYp47I1d0XQR4RHo7nLz6g42dBczFhAw2Oy9u46j
dl/tDYq/wtarn5hYQ5WyIUW/w3b0NL9+0FCykZZQYH/UGvR9kx2VaiRsMpXcK4Rc
uiCpq1cmIE6ZoZhO7kc2uwYZrDK/G+bfcmoZeJCUdSWzC43DH1UZpuKkdM6Rjx4n
/P0+7jw8cjrFa/GdmVvSpJBIempObgJG6LOcXpP3H7Rd8csx92KOG4hS4Cl+x+Oi
bG8spHYzUoJgL2ri8TfbkZR5DCzSqf0NV2T+8sEH3V4ec7K4iU7gSnO2w8QeY8vG
UWHrR6LJJbbKMs2ymYmMx4j4DpldtgMZ8NxApZ1lsOpZ5oB36oXnoiGpnnng+CuH
QXpW+7BUIm5BCXRjJKU7/Q5c/uNA9xNuBh23wlDOyEaF1F4qriZLdIMrjmdfkawu
iJKancE608O+uw6soiHE/9aYL4ZbMIPBrAYOXFi1dckhNpUkRoBr6w3gqKHneNRm
KXnpfitUiGJGkUy/W7wqmjKHv9aFPQgfqj3dz6kxvdJK2RhrejWCAzCykfroZscR
jD4HMhyB6Q/JhuYta9K/GDanl7z52z4fyzVQHkehp4VrjCsNzPUBsnCHAaTY04Yu
odPaP31Q3ocR35I9Zu9kOjgATsF+IdfebJWERecCCaKoeW7vPKfVfkT8ioNtF3zv
YGrKUgW9RGtq34rblrQ702xX7k/x74903anjtz2MWYAw0psue3or+oi/kXhNrEvE
PzxUHQSw33pBziRpZ4trp9z3IuY1fkUMD/P2xmnGGH1fuTLLQN39mXDGoSCyvwNm
eMCg2E1eni/AESV1pi3bbOhhQSW7PbrQqiWV6/Sw2ICE3IeIQYWopPSomkBxbOby
fxSifLi5ZqrQGu0qB2OZvmLePDpYSOcCvytZeJGytEoiBvt/vpJsv5LV9ES77BcT
+WQhq0G8MEDxitIujl5Mr7wXyyicZWU2FhTwKqjvJaCasOlbyuWJrcNRN7cbyJfl
T2rvanIFaKtlCZy2tNWScJiH5vmWlvdZwUsjWFqjD0O50i6VHCBPSfpyU2mV00S2
OWvIF+giF4wLPSmnmTw0aEtFmqxirE6iWGI//83ng/EhX3pfhV4LFvwyqIwHamLJ
RxZihxdIS2zTR2WX7i5gAMeCIT0cIn1jp4cMrS6wnc3utZpK0gGlpDeDKXPl/aot
GiqGomUTjQedBUqv2d3svgc2PhyRPeeOUzGf16bw0VDoZkMzTyMANBSKVgvIHTkp
Rvr9LUwJH7BzCApCErA+g63Ir8bTOlEqIIGktnqBF5t7sp76ZtEIuAQHp/MwpIxD
h3daY/j+tqIR0BI/7/HliVpUcfQNAZQUKBBaRFNSfKIUm4+RM9eBFxDpvdkOY4ux
MVSrsHabLBZc9MFlaTSCbrhPw0NyBXSmKblMLirFox5g2KGrauCRJ7U6bgWz0/iz
h06dW0phD9Julsp+A5HlFcANWElFOnQ4skt1c3v9bc1003rjd5u20FtNpOdXrdj7
Ub7xbFRARCqc1CPTqB83DizF/sVR3CuOXrNZruWZ0hflVIU4Ru56TWTpwg/EEhd+
uZfvxPzg8XdleyDF7niD+zvy0725SPIP0rIcyHIkBeDVAwgIzybMUfeI9yW1FXGG
bDTsa06vn+kXH3pEAbu455aqm1aCoZSOscLrQr2rZar026HLTbv+TOmM5yvi4gJW
AExtM6uLrYEalywV4pc9fe6pKYxIWYRp90uLY6MLlCWVIp8uR0/51Ts+BTKN8O1t
VXmMhESYFc+qM5O+YUQJD+XYvRqaU9EhWp68+bhnwxEzG9BSXTioVndaRl0fiALq
P+kg+dYDo9bLaYmi3LZbGRKYImY3EkfKTN58GRQpKmNOaSwt0uNZI+JJbnlGTnmO
6SFSBiU0DWT34nbFO2RqfKzjR4HfKm+e/wJA+c6sFE+sqwUedq4nJhYSN402700a
/mrZx17HEulKBert0vfNAO8Krn/RUgvuLwllSaSAzDEQcemtJiiHfLuqAfeU8r8W
l1deeWBWnl8gK00Ad7nZXx/0Bpl2rkA+cmx+PCfGZtUQsD5bMH8dFx2RRhqSh8/k
Y1ENP9cTZkSLqtM0et2ugBR/AEombSVHNgX8MPWM9Ku8Kg9yrpwCkumTfkY6VJtK
z5Gw5cqX8X3tQd9cgdEHzZbFs/tMQ7ZnFDTIGef4qJf4z9DrM7tEScBpcYCz4T33
HtxpdTCO2DDq2iC/4WHQIcNNz8u5wzWGL5mKY8g0mhhRyfMl7Ybhu+8KzjhQQV2z
CiaYMYXZpwuOIOEFmmtmATvKdYq2UwTQ+vacN/HN9vAlO0kdQSs3qHhTWWDV0+cP
OlVQjCSyNSUcz2kT5vTzor5ap4CpNg7T+qgfGftTq7kvlWhLrXGExKv4NDAWMYUF
m22n2BbkMX3rEzpFmJgEzptpYDhg8MIgHutklQG/FbRrup8+Urzw52to82EfoSiz
ElHEzS5G4JHXdw0W0Urei4SFaH+Nkl3va+2I1V0MuKAaS00TRb+3KfcG00i19bJB
weUGFox82/uXak1Vs7s2CQoTYE24PMbpw899Jm6oL+1NIYLX32jyysIALia+j5em
1MasQo2nNujKlAMUUmTTtcTWRPD/yhwjTHC481SicL93rAPv8LzJOQVyq82r5aQc
//8uMVIIKqMRsIQ949ZnR5Os1bOGPRu2z9lcwDpwl4OXuB1j+AlmXJMBnYfB4+WN
TU9U1uwhfzXcaDRZBe9wC9caFRPmN4E1qenbnIhkJE3vaOS3RqHQRqORC4Rw9eCS
xIzyUBRAXdqkEoQ8bo/oITH8bBLpNOB3x9QcuxSWB0Ew/KWhwX2Q4x6nwIMoZOy0
IAnj/XZ4XkZRw5DSUHjp6MzQboKVShfWYWqwKvB4I2YPefGUbdTbewTBnjxlegwx
dswDEcM0MHycW4W/8DSsMUJV/6yK2+iMkjpCZuIOvBsUXc4152iBSun4L3JcUDbA
IoJzPfLvafipHkiPxJfCDU6EsUriBmkzW2IVT+w0o3zXiXLDDVpX/tUdPYCJkwfB
vtiLfkaslmzm41trImVglUqDS4sQi4iUki182SeE8KrRWoSjoZ2DVTo2p3ENDNSR
WZ8cJma57lmRJsVMqEUhcevPMaxcLooVYY/M9ZaSrhSkvutcyWuybJc06l9VKk4k
vGp2SC6m4Ky+fMSauuhjPAEa324tqEcg2A79jam+fV/YrWUctmEbGWJNsd0836R3
R58uVXXF3iakeWNXiyC0dDR1eROs0mQtHTu00HicebSAhiHIYu/4lNK8GoHwkh8U
ssQKqOmJNXQBq58v1bRAcmRg3crtOvNtYUOTf/x31gUtXkmh1cFLE/Hsh2LVFHZq
+eHXqMvLXfFhvpoYbIK2gEo60uuoHK7DlhY0G3ePfFHHmhauuFkjsWUSbPzv0WMg
/ZYz/LkUI+FBKApO66sr3rKjr3UFwEwsf6mb5RXUbt+jE6TCpkSQFbLNEQ5Bxcnv
3FaGvM4+ZZ5wXYqWgdAqEcCUO/y/vkJPs6caA4lhSnIRjBd44k/20FKy04pW5vYe
2adEakRND3ar+l68Nko8v4Omf13LyEkZAtGS+zIYV61xtKDW0IwZPbjwSRidaAPm
Q5i1enn5hB8UtbJnKJlugP/vPkvfUqK85tTmxoUAQRnHOOw21c/9Knb+eGkaEEkc
q1oqeBcHy2+IRk1Xk6bFILLmISnvb6bjt+tXTVdaoFMpe9KPT9pv5j3O0vM0cRKW
N/vPqQpQggKhnat5/PEJh1/u88Lq5mk05KHD1Gon5zQykaJL0hzhKcLgYDq+WHFT
7pMJJwY4U3u610oBMkbXK2W+PIQW4dtIVZ1UQtl82VzpdFSTKQ9CcR9KscqiRXRp
TR0YYRHG/mV9Gy1SHi/cbQMk91NmPoFDHVJ0OqVa1nHyUwdO4Ghy98/7MOU4xAvl
4y3iRvJeV2dEjaOIaqr07YCfc+1EoF4q7voZQqraFB7b78iyohXRxeJ0J/d80ACC
Ib+8TRVDpGTWX/jQRHacpYte8RvWiyaAFk0n8cNSiuCngChHhMiGeWqC8NX4XKh/
LhisUCR2DuC1+9x8SzDzPSbQlEMAVeQjUOh467qJHx+FxKL+ujKd2jKDVExtLDo2
GMeTYkp+IohBDDwAghxZ08adrn25V018OFOUkenGrp/nMgi814LBmO61GBvewqmY
e+1Yz8WaSZJ1g+lyrp1oKlj2mbVdZm4qB8qwCAD9fgy4zqM5qvS9/0m+4mDNj8k/
PdR3sy+gswRRU0ByXhoEn9UVN5qcHNKtwY/AKY25OI2SJqC0kTLOPINPB502HCVm
tu2p5qM8V2jzU0e/wO9UKT4+V9Exti62XVNWmG9LrBjpAK5U8+iiXPa1WsvXtMrv
LB/4aUV39ybhv0mKOXwAZicHKIhq6B65aOCXHyZFKH5RXKO2Ib66uA/CigMkFJMz
9A7O9fvDpbpBbBSwWXs2dB4e16aysQiY6Mht2eqhP1B1Z02j64IohDeROGqwD0KX
5quYAXS4cVK+I4j2edtu80D2TaHZEcxHTAV598wPJRokXfDEQrZ3kn+2uKpi3zwR
ExN8pLhugwptiF5pv7D9PMpEK9srzSIa/C0IsHyldxRoF1vJSEFgolG9TGgfcStv
qIOR2apjoP2u6PLeW6Ssivh4uZ1lyWUCCE1vMbhjKk4adK6abdxurkuk9BUPcE3z
c2LnbflFt3eeSiDKarfH/8OplLEikpUfiusJXtVzVzA160pnu5842WuNmQEfOWoq
eBIiw9AEs8xcjIwZ/Zfuy4f+jL6klcZKkrWL1h0cHmJgo3uOEKS+BqAucK1wbLCu
AP0VM7TacxqyRFq0K1GVy5yjNjEEKYZ27/IaDMDEpjzxBm/GeZI6LjoPIDy7AlGa
ylHCG6mZkumvXS0CYKRhfuvgexaJL9KDVeg6lSnb4rBeMATbvv3Y3+c+QhpaEcc1
LZeHvD4+kWrtz6OnhYKmOkj01JcuDvZNRtvTPUMdn2zmbhIs4mbtz/iEak/cB2eq
laHcTIcX3Sr9CCy+zKUioS9B+0sqRz1YodAFvXiPiK38uIyI52afGjXXAsSoiTLU
l+KIC/TxJ93hpfvrsZ1jO0w+VW4KuLY8S4EWat623cQFM2//keEjCqP7fi66F0aY
vYHnuMK1Dsu/rhD3mxlWKmb6KnishaztpY8+dOmkdXnNb5x3tBiK7C4foYix4ldK
xkwQe3zYEe/LyFJU9AdP1AouTL/XJed9AnfL/W6NNnj2p7mLbUwUcyBLRiywUQ18
T0mPSw4eZM+C6IMAo9Fn9C3O0mCKmI7TC0E4PMr+WkpbE6gnElUA/Wh3/jkyEn64
feRPERnnYBTJGOnLRUtMdHTuIoCAjpygY0XKSYS4a9IGhxGKzfCZIHiCXhNTj+A+
tIc2q/A/IysEnpamelR1iJroEkvODuX2wj4ntW4LLsSD34b+af6y0zS8Uixu2rVs
QGOwzb4E+II3+z+B0CG8IAJK7SmllAJv6HtgQ6pkqGKzy076AxP/mEsgmdSoAvxg
+0JDTcevx7HApBmG6jq/ooOkt7Rvw4n/uUghlVoKzHo2dmv62+gERAOlCbQWIJzf
c4hjYBdiZVXQ5SHfEin3ZpgwFiQKHAjs3K9l7/mmaRsMYxqmT4uGbkSP978c84us
OCupOoaObX39UcAgebvwyKRRFcGRb//X2hvyWiiC77Os3VP4gf2iuwEpr0cOLFKm
zIlBhhRxF/G/zpbrAqVCTDROXzM3VamB/zWR8yvaADAgcVtn7gnIQ0T1M8tTM5At
U/Rgs8J+NDjMyghHCMz0JUFMk5bQ+S7ZHBQhQX6PCRUP6HcqGOgxDbdYgLwHixjK
VEAXqbPY+yq9jjMxTBmVe4GFMWd70LNaomMbqcpOxUi5EB4xA+xXBlrZHHs5bYVt
PNpsSu97Dy2i48BNurRelybFNsls17VFeScdNnEj1O6nzZA5HSGsy/fy45Gp5S98
L1+71f72DWSMaRjxklBlkMUwTp/txf+eTgK5qYwxkLp7M1WesVSSimmgub0LocZ3
q4UKTW+DkWDt/TcStuvgHX4Pj6YQ0oDJd86rbOB85nrvW7Clo5q+3xLRDVlzfUND
rpibLp48y5+tHsTpedB7xh64fzjO5To5hUjvYwD5d2Zao2rqNCT2zWwX9WqoZ3OD
yqgv8ko5EKIWQaaPzxOkIS1UYc7xOOiAcXIP1tl6r3Y6Bhr9bCW/KTQu1s0CthS4
tnwhtmvoo5fLpZ63WGA6b8uU6LR1ToQMV376AKNEuDT/hcuUQ1G/O6EJQ/kNu0mi
hDpfdhWJAQ/g9nxUFtpuH0jaROlnbt57AuG1ssb3eobgGxcrbPCJa4gu5YCSr3bb
1xqIcWoOU7+seyeB1tRd9gDFl96nueesSPgQTSFg3u4p/jFX2LoO7LAblpyseYo8
uhd9yrTo90i+ujNk5yMFoxRp1Lq4aAtgQ39rHnYzuDncJF22FoTCgjnpsOgxAO1g
m6fYPDoaxD87nZCZLD4Ot049a0hZUzrQ+GA/cjthv8rRQA2NkS88o5sxc0mvY14l
LLRyjq89U+Qm36SIwcDXerYX+o5prnpWqB5cItYP5ydAWmkZwYo0NS/g8heYNp9q
T1ubqf911nShxDIl90rHGTpicHGBIOrXK7FnWeknkjFU/v5ULJ0R3uT14wDbK0iz
LlMeAKKjfQxyazWFXW+UnhIuk2JGnhPkXJHv5ifL+KCR9RcKZ5LlCluRUPv2qK0O
G9f59cK5K0AjtwbQjKppaiAjdKReOayiZD35q583kaofZ+OECvTP/QmcKYkaPBUJ
LsyxPxeSPXHvqDV35zO6lYAruVcVQbuwYd7jT6hVqbHVnWR3/SgpjI7YJlmsbJu/
rOv+o3s4Ddx5xFgrjC7Tp1TFf6UNdbwHGKs+WNUKI3CSBQ+Meegxynkkay/tuPnA
oPkpZwQaneSVe6XyOX+sK5UStFLNd39a42ieditBcRUpY/jlT84l4hRM5zsEhgdw
3S5mfXJ5aKIabiCPBoCFnw/+qqsW6XGAgs7w6AylAf5AGWNvi7hrEExR7xNbclZw
/7yh71zuRDvxJ4Rh8v7InlqJjmOHVR9evwatxZCchLd4rb0KdxewLpMfO0L02UJi
v3BQQukZhC4V+Uthtzg9mtRg1Y8tNYMt5og6vnBZlrnB5H7f+4mydMKYnoY7mkmB
5Fyv7aVhq17gKm5qPBjQ/ats0ggHFHhVnOgQVUcFvwZ6HIMInMUI6tFscV7ubFvV
rHlEPGBHDBo4jhwHGhk5ek3T2PgVfu+v3dU3JCeHYefED3t/Od2ociHyvAnZuv7N
ZeidTlY3TtIKLJeG2za4HdFrIjyl5XOEae9pXBv81+UQgpDFQdtKjyZRiTJ+a2DM
VuQzYUC0RfYbYqMf5V4WMrnW4NF7G/9ET2RpBESaG+it+wWNwe65tngZzprQtFMP
m2cy3pEVHCQ37rAFTZApfTih3IRvxhNDUJQbP67sRajceDvJgbWUKU1eWyIv5VfN
TO1+UDSXvFtnedNgx0EFETDzmgvIay/u2MTlsP/XBkUPAW0VYpIQPN0iaawFwxkA
/X2SQ7br6FYYC/pqbiPy7fzVI9H7D/0/vPhtNmRM3ejEuzrZmicHAqScQ+nMzqZS
MuH4wXM++GD/VYfqq5XnRpNztYAmiCNJLzK9Kk/lgBi9PravYxulYTAyOBcq6RBU
r8cYvqHnib1Dst13UObpppzcMzwoYLf8mXsmhvy2KuQhpEP+YxTzSjsvCtwAXh6n
HhnFKcixyAh8XuvdSbrogZS/eDSOetKjskq+xnLnU+fUZKo3Ir580gc3JN+avC8H
N/HLCFc43uCcm3C5030BC75GPMOe5iWlNspQ8uZrWRjjkeIFYo5MYSjNCVZn0ZIX
0wq2nPu3TbTqN5ev1b7igP4xP+DiDjj0AP7hNbdkie17BLJIKGdlSsnNBIeMuzmV
esR9pfnaNC/IfO516Smc+zUYxeOFdV7uOpA1VqIhVaym94i1sgQwG+KgllscP8x4
4TbJmCm1snH7FM1GEC76R8BVwumOcrGiMbwc7wSp8FjN+vtHWyaFxnnrX96E/pg8
iO13hP92DEE9z6ykz0rYydMQuMxZaeadCuIFiaPsPlZNLdqViE/ynyJZQyovs2dR
c75rCHzzhHgbBCBLlxoI5OOZhT3N/U+2z/t7A0OdHSXFJQvmj4/jB1AMwPCvN1rg
AdLUfSqKtQsUKs+/Q22LLFbRQJdDcKQSuRjNXLfpfrI/2LIL6MtS84a0QWJKhQmS
38RSTcTRgygTGUSXsanDWxQ817Dm5DPHcQCBd8PBlOMDyq2FTMireATCbldoQaSz
kgAxHJ2bF2qakw4NscVMecmySSbqFWenwlVVCaWkC3ThE3cLZwXKE2Kz+eOSB1h9
gkI3tukOigdi4d5Nb81sY4GLYHLuvxyjb7uirsGsZWmBlo4gGuQBplEDr64Ev44N
9UZ5jazxzy8gbksqsqJ7bDYetsZuaCfgpf8puYk3QqXz/xx10YBrlQ2JhewHvrfD
oRr/YHSkyhQf6PCdD2gkZ4s0AQYrVZsKf46K9S+EfC+idPUl+UN9vkMUyWtOJvlW
fL8qcoBLEVZ0ay1PTY0P18Pe0BGV2tWB9NMqBrK1DG2N23jekUL2+vv+2mckSoCR
YeMQTbeCz+FgNge1QfdTYFQcD9SLcz41yQh4Im3EuU4AfgtG41aPR1zxEx16Sgcg
JTK9pNApxIpAFBHuJKKW8P1WDxCrCyNYQdfTjN4sjv8l4XFNOM/hyol1Oa9dsQ+1
JKV1w+WQXLecigyuq0KjjdaXDhuT9o5VuDGnOKf7wPpW3lxxRMp81N9VhuOfD7Jm
vF7gNhtD9nQJw2giUHCYwuw8I4UuzyXYUCktz2etxrSkAe5hwHUrlyR138j2U+g0
dFj5F75cf8jBLI208vGNvlrFRur8Q4E14oClyFQxCxiygVtrDLV/nYu0KR5l18y2
wkDzdqomUKrLtAz0yx+agNHbd4W8zw6i6UfqVXEbgRiwF0TwtS8ogCr61UjymHwZ
L73TNZU2HCatAdd/7+Rh4GpZWwhmEdSoKmRp8dwPKID1HR959pNTlpdICda9eXi7
jSZouMGulQT7FYhZzgH3+DDg0hcAZ7NgnARCwPTF4+JoaaKp8Ci0TnUooRztHygS
+r1j+KF3Rkb+CeMq87LNRfusg3IpEqhzZeNFxrpI0YWX2puk6FNy6r6sG9uu2TPm
OxNgkeMYgdY2IUAY8+3+Ih5b4Uc0NrVSwZM1x9+LaIP31fKlLjz24w39tJAAQWn+
V4ShS8u6QeJHzAHpOpMm3duR1vYDZ7G3Ff5GRaIEJklQU0gKuVVCQ4hTW+TpTfmk
J5jZ30Hq8h05wiiLqThY8hysT/UJcLN9oo85JIgE7ojuB3LEgVBxyGMwL5GYUiY5
WRXqiqCi1BGE2JIDNjXYZTk5VF47iow/3kMuACSHi6P2oozK1rLUH5ce3DcHZHDP
uHLu9yxoNjB/x1JKIUMNbMNekcXyxybyf8cfCkBv62/jgUj8SV9sXBHZo+V5pKUo
6YSVJH6NBBFsRSpva6ii0cE7OhtaF4ySl4XsKQ7MEFoZo/PO2xkhkSi6EVSJu5du
Qhmz2fBmR/3LNKeff+uN+IIh1sAlQKwq8f+x+shbk/ESNmv9+/jUlsx8D4kS0+nM
XOwZCb+qJvID/fS6RvzY5zGPEYeC5AYgeMG+1dAKtL+eyQY879ryaudFWNAcvpzG
KVcciGi59lfLxa7YeAJRESZ7yV8wVJVZWolTKzrsL53dJrE4UA+r+6vl4bpWW7PG
yo55Yw9wQAZ+gduvIk5IuGUhpupeytKKrf7nC2bQT7YS2rF2K+D1O36ikwJHQTs0
8/OFCTxImUZAmnsEdn+hlFZtMN4bX9Z9lVMK0FaFmFMQgMXqVmNGfNLS/2csJl9w
cRZ3BBgyZAewWzMEtWuhxVjYLkmzb5n4cJXdO/d8phurf8REwbrNuBIrkuQWyGLc
IqRI8mXc1Zs5Kyvw2w5iACD+ZXpFIN6VlVi0+SWiEnoOIOnGpRSJhIk/ocGXZ902
UH0i2P7dtuM9u+0y0aSGctpTXqvmG0eTtZP3CsqGy+6BGPk6/kwGLSqXF1Jn6QlL
xoLxCe4KMfjYuMyXk5ik0/yGYKDfGD+WE3g9suX+frz1f4+dgoAWCoTmwU2be9bC
EKab+dCajNofKspfsV0/3tB//IG2pxhQxkgWQ4OehoVQqX3KWFmRP6nhyRLgVYk6
gY+ya9ibhZYHTIuLDAQY0vgKeHevQFC1t+ihumSXqpW7+Zi6JFmwhKnEranh68DA
iraZ7Pj5bu0DemgKgxJ/cRPX3VRuQLnODJoYMvFseeihGn8OHSS+miRJ8I6e09Ii
SrQdRX6o0EYTorzWcqIsxUWEJuNQosTADXo1kiB3TE9pstlPMiowpd4EorJGAm2Q
10DNSKLCboX44yHJREn6Ya3QSfRNaKeOHvcwImsIUw7PGqZe67nXtvaScsgy5dLF
27TTgSiZLlEUUXGbdyyFDajS3nuQ5W5y9y+lJpomX56JyHwulH7tr5IGULpTASBR
C4bS0eaCH5FjbqS3p7PATDldv05qJBf5TaY/5cHA0p/Kv45uCx/207vF1ln+6g9Q
z90VJCJG3M/RMNGZfIKP/QxVfZ2MJpcXZLUYSiUF0aWV3a+eY3ehvAemge0QrM5/
E7jeqZ/cl9QJlQeW1A5PTnSjmgEEANxWAp/w1d3y5VSEgw4Jw8zfw4+sOAG4HGWd
m7vOPue3rpmZeV4Bs7zU8+O520Iwq4+05mPNzp7RSrRbxzmlm9lGZk/zYb7QXpAq
zpsRna56+ChuGQR2fAuhA6vw8R5J1Uw0awSVvHCs0jKoZKe+9vx9PQN4Ju1Fy06g
gAQAVi5LKzpVkWn6rYzUFW24HpSNsqc6Aeiwuhsue58gd8qCtUaZfxsZzAp8KoUI
X4D7rJH8uhJg+RTQ4+RLQjndigb7i0JfDO6fqm9Xd3QzmgT396a8bX6trMzHhht6
nxYIU93nFX8br5u7GX3oT7y09b0zSCt4XaHoUi+pAcQ2Q9tDt6JZH2TSAwk6Yp7Q
NL51bXfuLBkUbXonU3VnxcMv5o6076F+Rtu+AXkgJpYitf1HGS8cFFtMyYdg5hZL
IsRe2Ml7DPA5xo+nwKZgBrMRXMzQ0M6l6lkbFIXaXrccH0+kTis0/6lPgKQoMPRM
+GhEiTnahm8EvwwRwsbCKE6kuMMk1CAg8ajEQYns+7i9E4sqz+ZzLVrbO5HzxSi6
+bKgrqdDpigjHZNXbvt/gAQLdTR3xAwlqdBua+Od0c40tdk+kvCHhTPA7377deCv
1ARCxh2th4GnrKHY87tTgre6azv5o8+xA+Syb+8ZV7aAcl78brDm+64yfjW9kFf+
balsco3WbYiE84G8v68yd4N5/wcdPHqD6xhETyo0VZ2x9X8FGozZT5lD9qAfMRcU
GICG3hGnaw3C9S+ot2Sri++5DYBwPpigh8JnemNuRirnG+Q9cD5rEBRv79s80IUD
ooKH4ZB8slUGc+kxe+tyVoWDkelfIYbMcvTotABrmxSj0oeUeGCY0d2Y/YYtELsz
If7sjTx/4Pe4rNqOCLrNCpaUyv+k2DGEMqAxI/ZcOSctyklZ4DsaPVLvucertQjK
Oiva+wFZ9oEp7bFbX9sxAVWF/EoVVeamJjCSjF+y7EOsWXnAYM4dWWFedz++I2Oo
rXxSqMlQJBPShYIabJZt9FDR0T9nKht+Mo81G1KJxN7Wj1q7uRmlV8ORHlWfpLbQ
MAqVmEth8UP8zApfxQWQmbqjOLo4Wx+R7oDgRbC70hfcNC42CKrmrcxubFlVnoka
+sSYys6XKfo69LYV1lWjrJS98JjfE+S2CCZryBzEB46BVJeMJFqylLnLLDj+sFEI
6er9aZ+17kMtEMqmoERGnYkqfP35YzcO6HLhFIP941VWsBzWjYvmpMyFyAbRMEwH
VnYs4V9Z9d59BiyTao3YCyXvmqs+/KU21oKMWwscQ4Cg4xJdy/vy6vpOef+5JvLr
ALQyOBjeTiCu8neKxiyGwxSOtEe9vjrLBXrTXvJX6tRA5mXLmfCl1/CKy8n0RDk6
1dtIYRWv/P9XJy2ShegWzxoVRrVcSlUFBoa5MnwokdgklzsALwLshAdmGY5xs8sS
tdGbMR7dFXFQ9tzira8o9piB4+ciZeaqWIPLWtqJcQ1gMkVvCkFRnsGqT3LbC7kl
Jas0I3a9+H36aGiGRt0xrCWT/gj2AnzSTnCB19634O2hTHHiKOHI7UtLBcq6Noeh
iT9F/j7nBm3Jz41xlThg3wZZD+UwLqjtT3OiA+jl91BGmQMEao95MCH7yU4x9YWO
na26NQh6sIBAGJH8DFKXQZZaZSk9iCz0HN2qq4qpuPJMvDuUZ9FrJYxqPytBgldk
igfvbu2W263nTuD7gvl/YwJJZqy0iKkOR7UPhQT/jDiWTKQrmR/haal/l+sMw+11
bHwsuKTHrWlbe2YVALUoFrurPuoqC2UvwdpM9QTj9MIkaWPuCwJB0LhE0anpJ4Sm
ZQ81ROFlBgN+X3WsLXS55HUo9LFEFIPnPfGxRzO3LUg5Itnf2ak96awNxbgXm0Vj
U6pf7MEjKVhA7JWLKFeUK65ftoblN+OaqH30ddllSCtIsj3RyHbfWVmHGcbYN9rq
3Ufy3/FBMNRALcwKYdySiRQgXj+N7zwTMV79mQWVLWUfEfGV+StbaJMdfxz8CvZG
gAjVjbGAt32f5DA9x/tpj1OkbBO4AFJPrc6qKus8WWXlQ98eenl0hGm/2eWgyURI
RR2PY80oPzeiZxNRCp42Trtklz6oyknHPfzC0U1sMQ902ekxkMF2Y43XxwmEeXMl
1iwhNl//WIBVScVel6rNP8Q6YEvHhzaKi22Z+6yYAOzVuaakoMD+mJHzw4h2ND3r
j2twi2BxBMLwbVhSvVX/muj2n+PqgD9Ygk8R3YRBGYFPtY99UOkZou7jXTWG+KJD
Jychb1cfa8H+ktLbTDyr/qB6PYXPo9n4aRJBLFvYgpemf07AXdEHyP75dFKu05Ac
7mp3PxZOO322HzidvJ9n4fQgO1JIKCpk+EZ8QQesItLGFZJ/U/tQGqimdg025YFy
7fuY0bxZ8MIW/htbldqkx7TvM4IWic1XPpwg9onJAQ5+bfpseRlsR/Vdl0haIigt
5gsCxf35QT3xtPQujdNbRzIBuBAgWymriGd9CYXsKdzVOMvVDWFAcLtv2OHd8v2g
k+cDov+kIgen7r7UlI++TIMjoOupHK4vbaKPhXI2951XE6QQJ+qWtboGHE487a+b
CjV93UpQF3w3YZ8zwnn/VtEj2p7olTheDCA2blU7Mbi6YNZ83v8HqtVSpSpQWVn6
nDGXJMRS8fVm6NVp3DUKj3BWteBt8a4/n1Ke4Tki2I8mtHShEpFrcX7JQ9fMUGCq
9GTCXAcAfAGkVyi+LcCLDkK8Pi+klmiyDlUd5LN2xHBfCb86LzoGCRSIch2vjPFE
YJtiqXLIzFM+PhJ927Y59wINe+b8saOxKeiOMs62CFdcmdbrJCFFIvsdyKUYCkIH
J70fkagyPlCrSDvyfr1ibgxEGF3htcdrOnyzc8vhj13RiLvLNJpEF//oflFvM8J1
MbSNdKq2B1UOzsYzj/jgmvFsB10jS9VN8/IISscf4j5E8k/FYvxIiXdgSpMOfomq
1++Bs3dRm3rHXMh/KCZvjJayCKlw06igPTbATY21AUEAW0jSQLkrBk8CuFu8BpZ3
JjFZCZokDYjEVIjOG9Cp2E3cziRuogbiFsjNpWAyfAuFWLu1PZUIUZGv0f2E85lk
y6Yy5YTl2gMjY8ml2fEZOI1+GkcI7VkKefFISqxC4K7W5r4PsGc0azUOIoll5Myt
ou29ssbwEm+A5RA948x6dUC04Vn/RLQu0iqHKgKKAhsko8wninKjfK+52/Y1BPZN
kiXu9sXZ0Zg8dJky1AT5lLQw9+fscEPt69+KM6kpLMwUwbCSkGn6Qb8vsIOCEcYr
oQ6ajzn4bL2KicKe5ZDlGL+Z3YKQssWAlpWZ8lhhM+qIKG1+erz3Ws0FR7xinD3j
teyjPVuDKeDAWmqNTHV5h6Oit/355FdqfAJ5f3EOswgRuaG9fVulqq8QbFfJTrJH
vDmwasQSbJ+hMQ9RFgBg5spWlwoAfmoMqTHT7trFau10FB1mx8uPY1x0YJHR8c32
qc4cSQOxEyLXSnS9v3KEnq6h5SjlHcCz+eROab6jVxlDckD5kjn/sXu7wg+dBnGz
AZJVrYrExMGsZCdeXUVimG2fuTfivsODbwWq+cAZyN+MYVm3UoDkXSGLvZ3m0deo
tikgdvf2sjm8/5qkzG+TAdDQnYOdGDupZ9vzK63KfqshH7BM25lpIvn2sswmEYnt
ZIp1o8l5RLc2nHeipJJ2v6lYl+GAJERGWRzleKgi5BTd4MI+w++dQ6yfmhSDCu5T
ga+dGC2jfLb5bACeIomuFwR20xHB4vsX7BbK3kKZGaaJVWkhoz2x6cmastaGsLnR
M7LIZuS7ExbQP+1gKJ0UZlXp4OiYdioEnKAPSlook8lLbzTKVDLTfE1mSuFp6FvU
laxv/KWCFG11voz6zGml8E19mvCPr3HVC5YLiCfyzX34MsES2HtU0jRN8xbw47YB
UzGTWgr1Am/88fTgVy+kqMaY2IjivmRXCEpxWpHENEvp/WL6qDAt4bG5sqJXqPoL
yUUMlhl8bw43Jz9UCnl4cvWgomlKP/0bDxQruugWWDAXtH0ns+oTgiV++3hdvO4w
QNJclKtHdaavDdCwf/JxOpY/EstgMeIWFoRNBlG20ZCdQoezz0t9PSiVirmsOZeI
CuustIoNeDf7gIROMcCb+CG4xKa9oL+rlaH8YFkCI/8ZBU8/2OjuOQ5NXqzWHpod
Ofae+ZEuCpI2sXbntrDecfiwW+pqswCtSyTl6AbiMD+1hDh5GXJPerpKcgeT/0D2
iVkRZvsU66ixGXdq5qsGmV7gqHZlVpSBp/2ofaxS4VSKcUmNsYCxMYSc9rXJtG1r
evt1MLxgencqZ2Gb6I78MazxsLmCdYVKtzLkT+cXx5BUNeHoNsQ8z46H3QfiFZg1
dE2Az22okk8gxP8xKPuZVHipPN8Lj1STezK/CsitxR1Hkj7mfxgL3TEjZvq93N6R
UroKw3C53oKEAraSOkxALfohBt+1AHeHcBA2FWA4v28KWmh0Ib+GLyoxhJB6ilOE
SACW/n8l0TJmAx75O2+sopOcJV7RdpVdnlkx5UkMKZ07NLGOh9dy0WQLLY9zADFl
0FPu5gXAT0NQ0LIH/HGGEXtwVOUCP6numhAGHag91FWxUgzUcHxzl4NPGEqpsxuM
1A01wSUFPLLCOH4kfV77u9T+Y+xHEgi26E5wZKfOxl36W4O7MAFqZjMsYJpZk4Or
mmQ/CETLWhTtHg8yKY1U3mFoAf7CHcBqOvZQEgmHB1P8HRi2T+ZimG5yWW4wcfYX
iLD7cdF8psl+K4X1OU57RvN7nDiBe774fDNix8bdxJly/YrQ3FXOS1qTVf4ToBLL
s0heEWmenvWgT4gV7nsbGMZ6kuM6JUaMn06SQe0R4U9SfXQTDptl/zDwjzUora3C
6Sc/VdjlRCp8/bkjdBm3RtrIyeovGpJagA6CH3E2eq5/8V73Gj1L40Dk4PwIUr1X
ZC9wzBMVrHCAfSjUMKOo6rka/QJ+mRc66csycyGDCklwfWXNzLZIAt4fEDebp6MO
WsvgiwyzOLu/+k8mfUBsdVmLNxAIZuNBOaJXjRCgeNTJhlTplN2pCLsqNsOcxis/
qWx+c3vLYPlRrs54KDW5ACUETxMOqspgU89CtRhhC8/ITHq5bvBDKHUib4vlA5v4
tbDMzQeKCRSilEfWRrs/0tixk+mUOyev+fb0DfGDKa0Q59+zY+tnU0XtO6ZYyQH+
GdgRpHPkxJLS2HxItmvtyPyr/d9nZAZ8fHdIgnPTVRPmZhZqxaVAnroyljHr33Da
RnnaCajmw5oJ+Qm09n/tBqKFQuZMVRn6FBBeWNV2tju9DTeT3HUhASm1kxyb2PoL
3klbSj8lUokJuqRn94W6d93P2MyxoIi7CWNdvpUjJyy9Fw+4kzCsBivQjqGsmnR+
DxAGtHWDHkR7loMcVKsPYwcF8WgyJRvL+C2J9jx6nO/RqIGm72dGOvE6eLJ/5f0r
mHbH8f7YVdY+yCMKq2vT9cPXyidTYrfmHbs00IiF+4CCbIXMTtNAp86IAUI1hLAT
GAdkCNY3KNaFhpPzpvzChep3UE6fsFGj1dz/IGPt9KsR8RSwUvRephdrkMwYjLPm
N4ulOPoP+womb8oARiDxD1KbJ9MaTXgBsCE5Uxb90QvlCkNIOJLHOmWv47yjpHpq
1HHJETXn8tPGHu9PhvaipdyTfY4MefqHPop8Fio7LtEqWY6N/ko687cw6NAswh7T
Bov8JPIyiI4Wgr7LegcH9zOX+p4vC7g9BMv9HFycSRzphlNVhxZXDA2QE67IAkG9
nyNU+dqXF+hupnA53FRZJyZl74box2ERq2lpsV9oLtDiIpj4KlWEJr7VrdZhusIe
bC+Uiih1BZchKvCqxX+/c6bDQrX7lqs5pv3AvRTkkE5p9qNkOGbhTpu1PCv0tEGO
icbcAJr/58w1fe+se730/6ZXqX6WLS1q+kwhQO83Pj4beTmo8D/y0V5yCkTv1gXy
HbEdG3bN43onAecTVj2F7nHhK56iBF6RVCsJddkV1yULy9KPyy2iRKLap0lPDfzI
70tzuW6ZvDNlPbD/GljZl3aqLa1IAOAraFt+jbYidcR68LxWg1R0Ob6XEfTAqSdJ
dz+IIFsDzmAVVRP0tbqzcQ7GPjlSSBeW8aekcU6KnvJ2zxA/dX006dJNKEmf9F9H
srTpNZK1oe6Ni9d7rC8yfva2GFQYmWxhADOh8CqVp9VErKTjbm1o3Nz5dkZ19V4w
rRYV9cFcNd0ff/wkaJ3YmL1iRqDI2IlJ+JtVzuAEOCckKHi2PtVbz3xs0ojNGW+G
PEAb29yUifTYrVxUvDD//CPLpDXDifvCcYZrIJXwUtrkWY7r2TP8nNhvKowOBc1a
Vb6pHuAjLjYsMBii6jvBYX2InjLWT1gsJlyOcoSnqLGX3R9Id+E59iCFdTBrU26/
BTwiyCRN1bVlqTl33gEgH0VlJ7nfp903TGINb3VUY/tEuZOs5Pi2H63BArYtJ2Ek
iwbx0AZvcbBCqZwhjkuyieRyyBkfsGjjgxNjKZ7OdgzsNXcXQp17XwaI4X+rdvZj
9RY1whTV0fr1JbVkOt5Cq3W3slgajnG87r3NCsBgRrR3HqvKp79zuWlYIMpw3mw8
1YD64JO59DMB0HuuH+EU1YKJf69fNUkazUouPH2JkV1a3oeC9LMVmioXQnofBIlY
+RsgRYaGUoxKyTVROe+3al0g38DXYo0cZnByLxzp/Te/RbyirceQDNy1Tt0sHjWP
3+gIyIzqbE35H6gJRzTTz3/yTJVBN+RJ4H4JEsvoqm3S9RgNfWCMY4i0FB+AjOK2
/6NpB2GNsC+KRIQUFQctcHznVvG5UsSlmQ8nUcnccE1STOY8dpO0At0Jxzy/+L/a
EgvxCMgmfo8DlAmtkVgj9Up0bupfdvwyd33GNxC5FDHSICIJMrRIaWDIy8/i7k1H
FBAyYx3HRwOMEVBdQX5Kpsn4f/cSQt6h3scuoPPkLIXzApnI2z5KU1W9bNn7uxjp
IDLCyM4CKyBUiM+tKbOAxr1LVfN9KHVmDhDhdEWCm3DmAMMed5Z800zRlt36kz9Y
9adKw1gW+DanQuMuYljyXXV/cuAIh1hWtst67nvbk1jBbG+tPiWvViqnkuYfgmAr
5HoYFl8+lrihSbqWGlxHgml2ZCiKHmcCnIPjvTRqytE2UeOruBOIiVS4z/cABGML
yuz3Aai6EzFIfJezJrk2kiq8NVnZYZxAwbTHJKBw2koF87vvGtpLMs1SXrzWZbzb
oNSs8rTsfMheO7R0K/xrvVJb3a1tTR6VQrq7Er1rbJzBjmTJ6deI9T9eDd7MAfJN
KQwETK5HXe2Q+FjzauuqXxu8YY7aveeAc1KggTmKohfvJVCq32+0Myv69jMp2EdS
rkAEiE2F/Jy0Xcr1JljJEduGDRED1cVe9GNvmC84mBdr6+gD2ineJVm+tC7uILbo
tukEW648Xwba5ZBeiv3CrH/OWyqk/mAi+3zzwy+bjtOGI825R+mDpmhXid3GyxFf
iB7UsRWrgWdKXAS6aLmp8LLMIBNSPuDSUsTkUTJgsuRYXWbcBCD7dqcmoyXbnifJ
10f6Vw8AEHxFp99urlDwmDqyHltFvU8F48llWqT3nQSPvCskYoPDrrluAZZsBm+b
PuRbW38sgSTspQ5x8EUQgaf14mOsRndYFmRn7O8X5rIfrsSQdQluP9WxJzduRman
63rlWA/NXc+DUgV9VOtxpyNHhyyytnqatc4mXM9JA9OWE+Vn7SvMYc5LSReKm4pC
2iY8XMSPgErvpgQP5FKliqtk2nk2Q1Aa1Ehe4qgGfaTe4qaFQtJ6I4Vly9MQl31o
md0lRA7uAt9tbxg9kzfByhgHB5AHrtz/MXyuKo8W6d0gViVT5SGKLSuyH/vfYglU
s11u/mOVlmXkXXxJ0iCXEvciASFnzYjS25FImucejPo+XAMGWg4Ry2yLXh+qpC+z
CQ+2E4qWfYqUmaiHHbZlVEnrIBb+mwHQ/WEXtUAS1jzPJDosMqmm4TDNVde+cbcv
mhQQckCrFyCzfrO4DyUo1Z9xHps7uGYFY++VhQVegQMeyC+OAhaeaCtziBh+tT/e
3y36/+XzvcWKdkZZHT9q40MH44NuNIo5K3HQ0ha2vGyyjLo66Zy8gQDSPCK06/f9
15M/utWaiKt6wDf6UHrFWhYWQYnwFWuDF8bIiRHoacg4nWquXhU7F6HB/WwilB1G
CztsJ3B6ssWTsx0bexel63YUOo0/QqaZ3QFErt4UHeVNwlTZ182naL1PauAZXGJx
7A2ppso9PCtqZOmCqld3ArgHPnoF5AYtATzg+0Lm5UsOv5aNdm6jgjsru1NRs91j
exwiiGqNO3J04Tid1zTyaY+N1f70QxPjjQa1GLZjiFuMRQHZB5MBiVLDofjz+NJ6
mL7VI1FRD6SOD7f6oNUabVNcl9RqlDCW+u2Co/L+1C3eI0Nllu9x4rRzwYfa/iad
Obr2zCeR9WFQbLScaNUFmPtZmbA2YBlbrohfFGGVcb73AAbWffAjETANiRMkK4RI
yWinh/by0Y/Z9UszUG4uXV5dL6fOGmqjq45B+qvoqJJWsTvJR2Sx9vmxkyB/Xlsn
gZazJuae0jEeWsA/Pu0+Q6w30xbEj4/Zk1+FuS1bXh1JnPzGnFNUS8+zXZseQvdc
4on0QbaxKdzpHjDDLgMHE4kmyc2kbtQz+CyHO5fubRts/zHmP1FuTaNKyRKV0rdL
DCwT8pfmV4QAxpQXVy9JglTlbHluHtwUSNI6Efib1vDaY+5aBhTYcixI//r51HZ0
1FuvR6B/ZZy8h8Z3AIhaa3aPJu3hdnsYEkBJjKIOpxIreefgE1RKCfLJvkMt3zLJ
XEcqpbLVeZ8FKnklyUhcfNEBjIwcHDpMIaenkjbfbwIOWOO7Lv4xapnEO106Oe4C
c5dUqq7TXtkPZQUrKvZAeb0Pc+j27t6+s12I6zEyZQ9mnCm8NiN94YfC+0ReEFLq
Shz829y8M/qZWAS20sR6pPCZ/lFN+cymuZUpipBf63jWW0rm3hhDj/sxxEPqrg7X
e2oUeU9x/QJBk/HcS2doXXuJPgosRGXtcWVecZBUpEHLGDwIXSGKDSKS8C+stdAF
hCPmeioLOuTh11KuhjOwV26TH2ElRDDUzC9HJ2hxlxpm1HsJtz7EBDSiDl4IZzCZ
7yQDaPRh/pJB/0qyZXZPhY+k9ac6w0dCQz5qdZ44WNHl64hz6zGOpwCIvtjMokb2
GdnnrO3l3cSgFyZFiUaBZK6iRd4Q+t6AwZgM9ofceY6yjJMhJrgzIQJd29hPMQ0n
+krroyEeB7BSJQa4t0Plg94gLgMpLf8meq2p1+KIb4okHGmiW2xgNiBXeXm72Am4
NK1n/nefyYGgsbw3ivfDfZtHu/1Xxss00Der5Bxq0hweMLvcRe4I8C3x4C3m41Mc
ve+heFcgUqRGlkigw0btfWbX3I8BMuO8nyBndrREnb6Ic1agG746g87J/NxOvRlF
r4diQMJtSuW2ycGXxkq4ctk9MqrB07hYmtrHSkFz7TFhZS1VGja6yfal8j++dOc5
7VjDu7lITdMCJEJxFfZDs8q1GSGJFBKbblBsCczoz88NuBJY7V5bslSuyG+Z5E5y
jSQG9A4oEYQ9Of001ZylEb03DANNUP4DBWwDcAbeURWvexsaktsCHoN0riEhG5ca
WyPGYQ61w6/fqCXA15FFVzLIb4iWdaNv6nZD4MU3m2aTsNUbcO6e9affs5zUyIAo
ZDgH9U3otqKkHOGkLpl/c9B9IVela85pnXEE5uyOCRXry1cXzugIw7U1O1mn8RQG
K62D3X4CXExTw6rNaTexMscbRHUNec9nXTJJBp5Xj1TBRiOETYDQ/awP69CsOlX/
EVlzRTmDA9GEku6a6OzI2wvPd8WMc+EOxtNK1I4lO2Z3UNP33idt4NVzWgyqmOMk
SLUXkF9a7KXrirVWYk92GgaIGr71ITD4TJt2j8IHM++pANZ22guXRNgG2N41X5Kw
uLbTZvrHy387NNWnCOrnA+wO3Qo4KgXLCHWSy3prf6g6/66fgoAx/EQ5fBhSb9Uz
9EWemkxpLk+w/WlmZtedftR/mapo/UyAQxyOHFDovaQSD2A2E8pWZHIxHrTqT6XM
+xtLybWNEqQoV9/g0fSeSnv+t8+0JiJ1XnzUMboW8C21NJrq+Qju/8Y9EVmaTVNz
lkJ20vjLpxILjxlnx2q19t2wa9zaZnC/BmPNY8bjXnwLMp3XRb4/AiGGvroAN7Is
oqdL+OKK/MghbJRlnxqgZtXfRrbhhT8km/2lDa9h5XswyUC4vFKwnj35D4q1srr6
K1QkRwV0cyPs6tWLoNk9lnkXXLq5Go7t+fjsqm4ynoq6JhWpiDPXyiZ3pjBPl3zu
t6vFfOGPLSL+yplNq7GCHlVsaqnhay+frt52om/nxVG4RY300yLFMd+LQDdbdozr
kF9Tnxzk03GBBpxi/qve39qujckIi6jZLwawzYVrGCJrrBF9mwKtF03Qio7Sxzgi
8IckcX2lFyYvmQqYsXbqP4HD+C2Vx505XQbktc5NrItj8sSdf4V2G8488RyG5WzS
yXGGv5ccXuwYUt/4GTWKM+Ok2fl/fmmA6vFUUbnYD9w/+IU29OOU7ljBAzfWMNVB
QoACywnPpjIRdKUbkXTWAocd4/wUqszszoIIi588rsXzugHDHBJmesctgbE5Sd3B
oT+0bhry7syPMItY1c3Kg1YBJ2w8gN6/AXhdFwF9GeTG4QVr7PK/RguUi8pbBWbA
oU5Ufxpn1yCK7QZJfStRpU52R98khJ/wqXGFWDJpqDKDRq3B5dtOdPIu7rYgTuV2
EdjZt1DnH/NLxcDTcsr59eHEm4kCidayB9y6n7jmO0FfUmnU2Dxj0fO+7CF5H6oU
wKUoVcsnR0xhTve95xTjVWsEAyDozGS2kc9bTnP3hcs3iZy9BUkxxiToFsBhMjtj
6zSUdO6Vgm2pBR1DGhRxbOIJ9BALBAiTxA8BNXnDuK/MSqwiOxkNxBg/D3Pq+BWe
7FteCgxDH4s/vgUIXXy6TpTQRkHJ0WG3QDcuA04v5p5BVxZZuIwG9+HWP3lO/GJR
UPpRunlepsQ6zuJY/UKWCMYw8tJnmtLL07E5K9+bOiJkNjYqgCV4HuK7XLZF5cZZ
lh/fzS+LpiHfYRI3hoRIW8lj4Lm0bJwxhXUzHbe+OZgSghpiEmFI581JmCQWDef3
B6YURY5GnGBc074X+60jWXSN/gBmybkuGR7Vpr/7GqIxbbILA9nPDiOOiq6o5zb2
7RzpW4zVeyUujJW8m/hxstAQaWl4a8VKNZ5O9V5vDbsCzPcojkwomUW3RvS7JAVm
RvDtMSwqEHDZ6/OaQAPrV9/f7N4gkhn4Pe3kcfaEiK6G01eNuIONP3ICtLSTZlK5
a80lyy/BMNwIh+JvjshVR8P61DEghgA41+nBlkQPJxewrLMKFqigmPGBTbgqP/nq
yEjUHDlKOk6TnyYuVtO8dmKY54JmIFm3zDUB+6nfKPi7MjSKuxIGwjjWZZFhLAGM
UaFfNcYNz3WEaI4Tn6joLHhW1Jq2jaFos0WuvCMLSDb2wtlsPv4TNiXXwGGpArsy
jp9KjXySi15R8Bo45pHbrdRO25it3JXk3nzaW3lP1GV5EGUwJgVcyZbWZD1uzxf8
4wXkQDz9DuLvlM7uAFZ0quPxqYCDphbI58b6JEyWo1+CLAvsHG/xWR6bxo7xon0W
Ty+f8RqnMBPfHQTyOLLDwx54EyVcQq2FF2XtBRlx1KGqFnmoINOuwOFSrSXXfbly
hE8guQfuY+MvQwSY6nGFoH4c3r0qtQy/YQ/KD1nhEls4tBMIqbA6d9E+jeCMfIVf
vCkpbLzUDpKJ/J9D1WhvPy2I7qxZ9/R+M+EUCFulq+03PnXsj9IrYTF3DFHj/qrj
YCrbMuDR12gxF6zlTzi3/IH9z2wEsFWBCj2vKTCxPR4pAHjAjfx4qOwkd2to5Ey2
8IeIbgDiG6xqXFvN1tin2Q6QY1DRI1k0yEr7M/WWrSj/F/Gk8t6RBa5Oa1jrit94
oz4uNeseJocJTdomwpvQ2n6/jvvXiR9Vakxq7Q5eT14HrowlySZ6peT+btDIWKUj
MEuPVB2d5IsBWftdkLmZ+8GyQYLOkvIXvK944JvuDKkAPxpavTn/pVgzOh2G9LE2
KxDfAC0lenq530Im+aAUnfxFlCdSSjCeG/qgvCqhfmdQ1KP/SxIj2k+z7BPw1Szd
20kJa4FSlRWZ83T0f4spXLwJwEyzQnojXC1FKIxT/LhWG3rsB1qscX7IgMqDjOvq
6UU5Lj1Acoohor1VVRWNTp6guMwph06A+aaoEU3RlNU6ivftA3YmLDG8V/MDupv7
D5xjBIwUBUF09uwVFUTH+vgKwtzxHtk97TBP+bwEGBQ0/f7M6A1RuUk99aqyPBH3
VM+b9ZuoUkZ3TEu5+T1Jti62F86kCA7fHV/1kN0/VA/erzvqiQbXQQbFtu17rX9U
phEyZ6hve82/KTYHwiNWM/YuxGlTkDrPL0lR8rly3prRmn36b2AX3p7hhjDLlbHx
OpPZg2713QWaKY+Uq7uZb41d0neaSf7cjvn7vMXJyuGWSsVHukHkBZerLUSEmuTh
YT7Tk11kR5UW0uBaaLo4tBb+btso9x46pqy0BzblhETuN6Hco4VfVr54Rn/mLtzl
09mrnh0rg/X3tDS/96CgL7HJ7slJU6n89FPGMC93drzfKWOCL56Caj9G3Yhzj9CN
0oOjcYRbbS9nFue+ZlS5ulicqyVFkxcoIvIp2ZOxf5rGXXgDU/Hl8BQnhLs7jFFO
RuzU7XU79UNMR8/dpz6THmaIs3erLBwldOpllkJv5FUINqvlo9I9qnsA7triQoxc
FsLVfTx3Mq8LPmVP8XWIoc1mYvLB9ww9BI6IU7DIkZefPwdwziedQxSNBe2TJMek
9h0vsk35NIJfl//qDC7KtF48lZZuWG+6KQgQ110E/MCRQXw1ZW5HihxPgRLtUU4a
QDzdF4kikBKSmalL27Pl379aWOhIGV23qGLHCRN7s2q7hVm/VMA3M27e7ls5LyzX
7OZoOJMHKwOihGrXFD3IFiuj6oTyUpLlStJxQWG8WmcsXsmtiimZdGieGnT0cEgF
I9DNERqr4QkY8kL7ttXuG4ueuGlTu7X94wRxnodwpTPpOryMqTFWC/t8Wo8grOIH
mwSQ7C3pqQHH5828KzMlxUp9D6gTQL6E4hJiq+LjwiJ/rFuaCIE4pfcz8jrC1Bzq
d9FZod2N1rxFYEBU6KGc4zZwxqq2Lq35UA4wKF1cJjkTI/fZx6/+OlbLdqUS1jwm
JBUtJmayFcw3omhDmB6g0ybmh2kIfSLZDVBiMEDZASM+4oekivTPLDd2poPxded5
M6oWRpd2ovz8xAmdnQawcX0cjL6Fx1bqcbrSg7qzIht7HgD2UkOHUeKY5AN9ZBbX
ZlJYFzVR7cGfjGuU9rstSKIo2kAcwFcmw+CO40hQls1B6kDIyvUVcKmoV8JVZZHc
hmAvxwv9gXIWi5UlMSxJNlNrGfxeZhRJ8BQ7yTCU2M4OFfMXlYY6TOFsvL5BX6yr
U5gTFuOvMp+gQvIuzPHWSjepVU0QFCOLvHK7/nAMxEscC2dzvUpw/71CZZ2OPBVw
Spy+v1ZTvFlsy+bH+KWrt8dI1WuuJIdncibK8JuuC7lN1gyQoQs+QwvcTbl9UQ1Z
i4tYsn3R5QlWts28GQLoOvJd7QsOrLZ1Y5lz89GZItLcsSB14GK+nMfW8vUbFtcv
6AvtZbKWjx+FVgLJuD6vgEVaCLlBUv13s4WTVsznLnB8rCqkVisqGhLD4OSw4Ach
Z70svY1Iipl9vbCw6iTYfq1B43e+CLnyDFC600Stcfwgh0xKT45FKYQeTHQ2+xFT
5kN7wotcjBDit60ln6j2jd7U9Uz19t+Bqo06+AZl5n1QEZDKnuy6c7HibfRFU9jW
7f6EpKKPICBRTrT0qcWYq1OI01NdViSCufLFnr03rgqUOKYfdt2RLMgOOI0OexMK
wgwRtlWCgxWL8ncfkCSst7CLtvtMb2f0+V9v668c3J56CRQS8IxyiAasoMnJrQGQ
NhCV4FSjztee+CNW7QaP/4E6ffsWIzLWhFfSRpng5dJqTHgDRC9mFdHBV2ymG4zc
jlAYcOiojBr2yZGmBehDYJrrxYFAYLGv7tuFV4a4tqBwjz5jtZkljSdrrT63BOH0
gVgzCnysksFCRjl4GOu9jvDHNl8+buXl3bgdwoo1edVY19MgmYkRrlHZwZYUfsIO
vnnM/P+fdicYb1Rh2wbsTvjrylNtEIYPKoXSqaTMkw3a3PNdEbzxPdhxpf72XyBj
KBXlxaQv0UnkMB6+5T/kY0knpGYghgNVgZsFR/hnSBOJ5hBcN5PtBqC7L2B/UzQM
QAuCiZkKiIKL8a10edDHRLmT6Q3DwMgU4o0CoG2HbkYcw0FA7Au6Se8PMLZQfN7e
18eDONVwKbg1e+45CadahItlYf0cVLnGQpj3Z6AsFd5Vr0OCHzmCHN4ZX+m2Swn7
83w4sqOzXsRIVzwe63uYwb1jNPKllgG1kDiX2V7cvnoopb9482Pcz+0G3MejqcN7
SHHTcoPtlJVhGlB1kaXzzllqO5Ylm/B4kXd1YJZs/OpxQH9j2qDcMpqzjGgkDQqQ
kD/CMLAmRlXT46g9Kcup6W1iQym7s3HE/J0jNepPY5XOOZCQy5Uz+nKPkmee0Uff
qaRDc6Wq5ZDrmWHAxf8E2oZmLqzrT5YYUK68PihRmoy+//r4gz0a3IAXEy0iR9Jo
E7dq7xcnikgPJLIxkl4AfCJSwE5PTvpojlh2DAAAjsWizcT2ywRhMm0/NpK0mNvC
ONMkWiK+JdqyKS7jqVGY314SiWr448tXAWlEk4UmWkmxWYLPJ9Q5ppWKtbfycw+n
I+sPrvrkwpCPerjmx0SaXJhvRtO53hEr3ktj/ZNr6k57UOfh8ehrfqSpPctq5JHO
NsbcyclJRb4kO4JdltAYxrGipY8NsZJHfPHO6oTFfYVm8nhtpz9cNMCM7Me9VKwu
UMzhupWzKP9dM9EylGVtatqoG+ecuLMg8M4NO6WqLBSNqm6BIdqF0PVDyYJb65sv
jai6H+Lb8xrsqLQ2N3UT7FUdvtUbtOZpB7kQZ2XOHrv0r7r+R1NYm/vI4qvppEpQ
epgrgR4M/5yhGo9oJ6m2ll0DXe92gNnRhSpUFdxBQ6rnwru1+NW9gs4fsBBMHcKd
GExVBOJMYoOt1G6StlQ9tOtL26oW3pi6Z3c1GIp88rJKWbwwWMTt6HV+MaO/YP87
cEZmzyI9NYqSD1398wC8eHjjEfOI+CEiQGLJGJuHaNS484uNkFU3gAAthJRfZB0j
rhmYHaCqmpsKCyIAA4uKBHs9JhFmEVuMGyRRO1OJFGPkb3wGauRH0Yj/j/vWZpHP
wSCesNvBPsbVAWvuoAABnSTKdZLb0rSJ0CQs0U/Kyhl951NI/OM9HIJTOURtOf2o
0ax/4A/h5Ik0Wdlo7kOHMTK/823muKAN9AsqbKnYbGLqCH1COxg1jiYF2b7xVi9t
IxQWipJ5DWB58pR9CC7IQ+VwF5H+ei6v0ER+HZQ/OoDnYfNHoEF9e3ZrjQKrk2BG
0Zeg5QUgD4FMSsavxU7wMCN1fib0JJU4H+OypV4gaes/Ggyt1Csicm8CHjna1N0e
zbH5Qe1NLHOGQqorNk2+Cc1HJm7hg7kUwFz75VGVGYq4VEQ8CpoxHGEtkxlkN/BQ
3vVVuWv8T/b8oo8wEEPQBY7t6oZPEB97YzYGoHDOb3l6lOynTrhc/gZF8OqDJz+9
5k95jyg8Tx3NvjfwaltGm5qsmoHuhDumK2OzblUwPxrJPRlKEExxVskzHMMW4K1d
It+342GTBWEtbwmLTwGy/yGVnBiAlwPLuUkIKImit/SpXyCv+hZ1j5mtnAQGufkf
piB1E9M/5uzeCwrNzSt2sSYSHXNcfTGg7jxPYKohzxlssIds+CskirVnLMvxFnD0
WRi2cYDt/+4tlAdD16hYAAoOU5YegJh/VJQ9FQgb/7c9e2ym698P6ZSLtzHGTqfC
mK9q4Kr8mUGFMxnbR+ARPUKijV1DBPT/NpKzC/lTbmsZFRc1fNS370h1PmQhqF/1
0pUPcnKOQurgiD+D5Z2NWmn2XILjPqiF5w+EPCAchwG/a1fPYL3BxMGmrA/8yUu6
tPh86JonAO/oPM0aBMtBhKUFvI9SBk9XcagtGR1VjjoaeZ0crJmg0WEt9Wirc43h
WGrMRtVErjQ1vmLu0ZH6nJUXFkzFtehpkpJKZ1Su3cTZkxzhO2REWRy50NK6VWyK
uXCNBQQ+NmekVjOIFHvzLwNlp/UgRcitLAfYiiR2KF3fDN5c4hsitNZyADXNPSdW
QbjQyfO9CP4zreXxIDn9luiAGpVX0OhCzoIq0u7NlRY+XsDjFxPArUAz2kaehYtp
GLIDYCjtivZy2pjUr+49avhRvWC1h4UhU/WJyAOKJOXR3ZLs0hr4MNAx8tH+lnXC
InvjwLG2h9qr4xzoPrdUtU2fPWPXIB5D09cjtlqPCs38+5A4AHZ5+i9PSJrZCJ3Y
Zr7oGGREFhpUp19rQmd2sAXUEiS8mN3c7lI73Hg0Dge/beR8JfMEYh3QUrVrHBPd
IAZrAKEowP83J9HUu6yh7zuwPoz0JN9ikqqjB8MflmHqdner9VL1ScjHDMqIZEz+
QIYlBQyj8BIKR2irs037baczIJAnELeY/Nf/Cr6j5WaCivakjLTahNXlYc2SyW1g
rKHQrQKuttjEUyo/HVZ/R2AXpbwU+eipedy4+CfsTI999rJrBDpX2W2IvqhLaAVS
RDfsoqgvJJrzjkPrMXMBn0cPhxRfJlXl7RhqxAbif+2cmuM5ZYsZoY5BZXG6/kRt
QNLw//1N2kCGUQzuygqICFzY6QLtSawH6YWKlKd+9aHeTqHCjOGaWe3ue6wSttsz
NDdkUWHHOhjAjl70b0gBjp9bxq0QJZCF6H+vPCgp6YzFAwhO5isbBAa9ZsdPAFve
dR9yf+roVAkJiG7XC8DMLmrPQVxm2jBujxw0TividDCq7dohmp8POq9iyAXSblyH
O8QG4Ii8yvnzU31EL1rHNlZ9byGmjUcqoS7/RJ9omZWCGyLqZfks+cO6lj/3UEIu
mSoPiS+eM3M0lEIX7IF+WWH8fJ+P3JimbQKxQ/cGkhDA8GGJC054OQzkNOkRvz/y
nqMlcXuFddUrvtNnaxiZkZor1wknw5OeDrvAlAdL3Prfud5Ob6KyC1EbROuwFDf1
UF//r/rshZBS2c6lHNmWfP7KwWtk9ISw/kMyBT7vlO46EnrzmlcD/dj6hp8B3nwV
jjpOTPTyyO6cAqpJ33MS9HSMqTBBNSPvyfP3F7TGloi7VxMZuShAJPvBrDD8WjFD
HqOMMsYq9k4VguvnFbHDnjo7Lg8ynOgoMIVouh/0qGp4dJ2HCH32JnWd4QSj1MfA
RFamGj0jgC4XxQtx9TfHplWZtjLzv6ET3u7SXG8ooD/yb6WLkIzyK4TLou7msCvI
vj1pAgoODmw5IAgfsb8QXA2wIySmTo89MwTuMECl6/5/bcPEP93YQvdUW5lz0YbJ
OM+8wK/h1mfRFoedJ3aIF++y0AODgHChQNVhPM/OU7nyWBuIoh/Fq0Yz/sIBT/Ut
DL/lJh3wvULhBakA+X2qQqDXeJjbuAMtHoYl8M3Jq17DpsLP9q/igFsFwhCtLy9E
B4jaazJ6kQGvuXSCCAuFVFyn3MvfqA5vOP2Qb8PEGlcZinqznPGZOKuGhO1n/k5s
/cWE5e2tLptqIERRHeezpeW/a+Nxf1EugQgRtXOqEfK10/3ODmfC7OewojXyD3oq
ajAhbuUBQ4bUOdjWgvEIhjPkoDC3g7ZKetxRTWMKxkWxh05KhJiQFOD2EEPa+qhH
vVDG2rqPEHeM9q84X8eMJiAiHH1okEvPIwR5Do9IHB2f+jXstTAgzftht2aum+fj
BncwXklWqMZQCe4RUyDwGf6M4vCPl64Zfb1ajupkhv10pW1MwB79y6H6raEbbu0L
jn1CMa3AZZLQZLG1TAPHEIx5qpLrKTkiHGkkOpUreti+VTDYjDlfcZB/UCpCrD9l
MmJmCYlDXgSDZMHbCL3Yjuc2GizPNcfAg00qPBZjYZ0+Kw/jTiSh3Dt+fyhk6+uA
d5+vGS1XDKvnxBu0Zqkfo3jP0ThyVrl4ZZaK2ChtZ0eCyN4Sw8OrV+K38ADpDqNM
7M/CTGDt8LwURk4gLLESzTXAgwQH8epQjQmPQyNDiunOinyEiZK315Rh8UsofYtk
clHWugUWzjfJP4eXDQhjEP2j4ayj7cAasylLf2Be8pPQBohUWsEHLYaq1sJJOiv8
OgaNTy44K7melt+LA3BXu3spEKwOGDJF49bxbqmM2vw2utsVKg7GCZfuT9ujOgfo
56Dge/YroTU6fAGbgHB4+YsoPECz1Ym0P4bQWAljc4C4Bck7syqNTxSANKrTZYfs
COZT3IaN4X//mqlqaTLTyaa1eVXlyde8Khi86rUugK1sbSb8UP+XhtxMz7RVKkuZ
gw7c1ZaKZ16CpJJTjUxXKDbrHb0pnOlhXvTe/zKQ6L8OJh+058dPnEmuSMqUvDwv
UR9j5EgtM90hqznHdCQJfjQPuzLhMoajBtLpJdMizmUHkiO5qdqV8P6PUuAIqu+S
Mjrk0Pj83sOLdWB7p9ykuXcZUUSzC2MlKCXRP3H99jxnJvoNHMmZrABgaIacTzNI
eSF6KZwjMGOUZElzbmkgOf46NLx/0L/jR5usKgOO8Q5MAr2XhvkKe4Qrtmoe0Nuk
9WpiIwA3GZwY6JuUIfNaimOrZcjpRsD0zBWWBg5VWfw/nqIspV7SuWruoomlTAln
qSSAKIoQbr5xQsH/ZnoOJxxj3jTCvY3w3JxPXydiE9r9xG5H0rgzsX2Uk+3WRx+n
OP23w6J/POdYHBRROkzmRSzeJSWNKQMKgs/bPQ8obCLCn9ZfuRQT5ipu0PilyydI
c9ObklG7cxYVeCTYBTwEmkZ+gSJ8VDsrvRBl6PVkdJpWoliYSBzV3rGTc9Wptkzi
CwMGlT3X4oGK5KUm5UuAQi1R7M+JTAJ5H9BSj2TnUaCY9c/XHiMWU2kSweo8FAdQ
Fm7g6KRguUfWrWBAVaK1OzzvPWozdsUq6JubQLmNWKG4vhD4F2PEY665eMnlK580
LImqQ55v2/A7+QY6ceyDqONdanuVMa0rCyXr+YaDkrZVo9FS4/FWVHeM9DYYikF1
cb70yfDjQYU2S9B5z9NX6nSQGukkBKhW6pUPaBZsOnCAyKftAP8HtISTrtS66RdI
AsbkxKahDiqH2ozLWvPEMRH/F0uNR27fJqxuUyvBY5Wvly9FVfk1G2WIE4nVonTi
JAQO36bOSf0+wxGKaWm/QgxY4YEVSXhLOKZEcqlI/INmM5bpBpEu0GmZxHU/8ND0
1MBcydOHPgd5pK/PQIIk4IpOphnpONtGSXu2mC2ATY5dRv4A9WD02PYZaVn+CF5o
7buTewUOjA6gNIkDelqs4oAJWmOAjhkMi+OvO8vtaBe1+R4niZEJwVNKkSklweZ0
jvxwzP4St5u9Q7dRP7AUSY5ubhsYFRnDxS5fb7UDxFlOoQe6PVx4xNjvRQZ1yqOF
/+zuwPM90oK7mckmxf7EuFNKFc8xNlcgsCF2/qZQ/xsfjle+5hDxl3kU0LkxCPo3
mN8RqGGLNS5FY0bOyrl2PuqYMASRp+MHb6qDYhcjSZl3pDpsAG8Zb1ZWUfcEr1au
Wz2UTTi10ih/rxAEZiH5/BMVYfyCo5y4pGHfA9m9NbH9QhFH7G0WYNVfdQ7Opi34
HqTQ29H45ivJz8GGpcrqEZGywarvqpFDP4yxVsMSi/JZ77WGnpIJjo3o3wecMuEd
ClWvbZmjtSJIqFXogoSNeEpRYEG59ie32HPwxSyHG3wKHj19Xz8gZTG15njHUU9Q
fdhGPqMXFPytpZovzcvjHY7hlB/27yx8Fc1lkgK9WVtkGLP4jCKyJ1fCDjHI2eBC
+wP9TM451FgAGv0IooLaw4cl/g7Dtm+io80etBHwqkgbN+M1N20V5GeRB3/TRi+R
y+nnd7fBHN3tLMsPM2O7Ta+mEGD2fb/Xz5bTYWBFwb1YYjkrG2XDuXTiGQAPujT2
KHNvyq0velmSwT/GPujQDV/buqSh6CpwsGrG07nkdn5do3gBfsdjUbVGUv5Lm3wI
jffr9j9CyYpsnHDfI5Lo4viStzqgn7RshYwgcahhcglIwBDZibaKMeU3FP4PeFk2
HFZk+dzMYVDcbWNgUWytHBINMBuIBp2jFUPWbdJFca4DNjDNzrwKJTcML+xicFkh
YtqnMyOyenqRW5KnTX1Wb3+iB8XO7jNj+3WbIx/1Scvz6DaRbTHtxUAwHrgLB0GE
G+E3bBsPoip1N3GDRyS8//F9FJEok9LF6dujQPb3hAlR4ZjJ4RbRU2PvyqsAOxgR
uBi2WXqmE/U3EEIaUG6VOOocfQtNPYlcuq9zmdmpEeuo03d2X7CxF1e+GMaodzZQ
Zl0b/6dHQJ0Sk6xLfxj9hFlX3Fh7TG80zlt+jdBzf/jTtE7JHtnI10RYg3kbD4y2
K3EbQKLCguzIkQYPZc4EAwIZ7biOZXHCxPEC0k+TgzlFaQU/nfA5pCNd0jRWdcKk
3zk2UBfbdWA5azXLuCwYxEBXFuauBgyLQ5mw7P6tdoFCx7jymbnAkm3haRe20r8I
WBmsAZNlRSyZWHcFWzFdd/u44fg/cZjGfotI9WfFyNvMQ5Z0tVs5CgT+9a8HJxUl
TW1ke4wWun6I7iRDamlXRgbRz805OR1DlHTA/wbAG5IFInLJ1R9O182QwdqqHaAR
2hYEPIM6OgZ30Hcp5ApeScNimI9k2dnwHsSLhxQc6IwEGqq9z1rPXKYrksXoeep4
ApF8oBWAtLohXzE059Duh71y7uIW6RdGdUFVeuHV+H3rpkXaj8v5QLO+gpSaEOkC
0rOuCYkvJwSjV6cOBDNUYY+M3qu454nzL1dGnCTDYxKPeFasCtQg5cbSjWlpQLFP
kF1DmnuxnxGW30t0C4KiJGHh/ETZaeXZhkq9Jk9gwK59FzAWY7LBNZXz+g/hY66+
zwzse8QFj5zsLDFTH/oU8Ap8GpMm/mIamzxQbZDSAMoguB0+M0JkbvK4JaNQeO9n
SAPaMoP37gxP5CB2e6wYOXNj6DeeoTTuUbDRhkIdTW61LLxAYUOxSgRR0Sg9g9Yl
fAyWchRuKxFaDLvqp2iQ90Oxx+vAJnSs6OM2T3zeS2vuq1Q4dO08qvQF+rrHISvK
o6KVoDA2v2jU/YZhibTGwhVUKBjvoK4aT2MG6L28oAclwj49cBJUd0M3gCE7yNg9
RNwWsAl2JOgGrs1lUt2fS2K3cvuxO2+xOex0WlKASIrEDiWsOUw/vgJWaHpPGDk5
FwaS0xn++IMG+4zBpVH6mt9xSBFZr4uWsY5aZ1Jqvmqpc47o/Mz5IWdavqpsWWSW
HMlNQvpuL8xnq5tclywhmituaagEObB8eNOoKTGnKRpdUegcDbgtDOw3RJW1GGYH
vs2SJE7ZUO4hMItG8uuj8dVDQXU/dsPd9fRBtQ/mNJjLA5a0honsx9WZ/YtoSF19
xVvRdW69tx/9npSQunuSZFxpuq66FN1X1DYPCaar/iUPgCpckVADsYm+OzA/12um
Dtv5hbOTh6SdFLuVyunn+XGbjNju1j91t5xCIS0KUQqSwYHe03VM7r60mCFfJi2s
n5iEwCBaWunU1efdL3IJc7z8c+u0LOuScZ+bROt+VwvWAnGZ4lWDTI7WKVG1Su5G
ZNM9JOfEei+hjUXlVdokmj/yBU6C1wygv1aeN46WGBxU/q6IoEf1NAGjmN/NdbOi
v8Z4phQ/Xzf5y6b9jHUMb7nTI0wu2e7aGRZQyVWrFPQhhhBFMFRs/OjyE4gkomQ2
3pgsvwW/4gKxzvOIDAJTI4j269IeeZzoVf+NKEm5LzqlfPXmMwaEAbsZXXAsTSKx
S+3u0J9RSor6ifpHjtgxtr8pPEo2dq8x2HRjY96BpiHvcJC72fuW+GBx/gUJnQRT
dUJO1q1Zj68FQioLOmLrthDAyuLKWUiJurNNERS8OOfwnp7AjXeIodPcl2fAWXJv
1Afutw9AMulsHjgJxqg8xYb1uAmGkLrdbaKq1s0/cdKHR63AMzrvdE4KGF/vDv/7
tn81XzvpbNOLgiBrSz1Jrs+JuGNXZJXugTvPVh+s0NZTojC4Le9SXNAYYHJRZUSb
3mDPxOtN7PfwZsiwvVqUKsezJmreD/hnhuybx1G+kxIBKlrlaLTR08c2XurHJoc6
y6TDUKY/87bxeTfR9rv1B0ohgu4grZQJD8Wbtr7Jw29bjJ0lE0JyQO+Jxy2RVf5A
gkUPgDpsEqsyywxJFPn1yGcV+1W6kx6aeCKekQvZvZoJZ+pNPR9zYEVcXIiYZ8HV
qsYPodqrcabuM13YZ95S7xIMC7IufkeMnFk6SWolBY9Tja+a6agnGJU1kYv3dQOl
nw4eJqZOUSA/8vsV3EhMCPXl8wDqB/cCZ7ExRCg86l8THsFLH8VOvSgugTuB+LEM
PzxcVHlEriaoWVlOVAF88xqPUITKoDpB/RSIOp1WATxwE/FXREnopO8CSjDfpFJV
etsjGCiKCD3aS6vDc8NaaOgarAeWcOBOA8HgqpCAVfkc1nHagqm+jdFg1cyQiD1O
Dq0ynRlYr45ezt6ceOrGqMtx8jWQwMI0jXH9ffwQobQRK8IWKMXZ9j9kCcii87SL
rR15FFl+40vWB7sFeT+aIYktClq31ql80gxmHj39Y2gkszBcgeft++m/RGO/lpDn
mIIFBkj6rbnGHaZewYuesrSVVBoMD+bFXiyBMkAPoyxJ5b+g46DAkOpSJ0NEZgrB
DuNTjJxWxz9swstswWEdz4aVLb2LJ3FDGwlCK/HEXaEub9KgM5oVd8CyJPy7H+hs
a4uLjlZt3FECsetXKHOC6SGMoI1seumlnr0GC13waxQmIi82VPAsVSLGBM7Z7k0O
C5eArPkUe7DRLBMVzOAdvSYzYmBZ/UGRmVEQhs/W9H2T303SN0ucgTlZ+Z2gwGqx
kyYIjCjfCSKoWiCBXbTdpm8cV4x9dXhjQAkYPmeEvaUuov36CO8ojFJHE54aENrP
2kq22GgZjVzcTbcDshytZtcVq7zwJ/FlJoYpK2YfXvtGisE8TB5lOCxCXhCApDKc
r76op0KXDTfd83TxNLwTP80lCuOyahA26id85Yi+fu/kQAf+SqyH1yhDWA1TOun6
yaK2SEsqh9ovoKDiqOpKRP2a9qUuw6IEAaZ6zoSPsy7sQ8TcARkOyUU9qQdF3h05
omSkm9Hz4Vft6you+1F4yU0XeARsTOdcNTxRH4rLo3cU93Tg6iYfbxlyNB6y41qi
Ssx+ewyx3zytrPngmMTWUeFzctOvEl05wMqYmvXSAhGjU49qOoD+1S09SZfgkFk8
hsMK+1u/WSpHgKuTdCy0H8Re6rtk9AcV0CvmBtw/9cg50nS73eYWvku4i00PfR3d
NsGB5uBogVoF2bEXjh2adEDUH0wjD283bauSC+XnyBOaxzFHiY2kDtTZKu50Nvpn
Zzv6sb4GVxMwZ66tQngU9QHbXlt5bRKHBPqPpODYpkMNrn8LPC6rPT1ifdNQlOrX
gFIOpV+/o/5GJmOpeiKlrh4Cd2j4HbHuvCUcB3116VfxKtSY3FxcumUK5HutE1VD
kjjqwN4EqTMOB19IrS2qaa4bLfCEjmQrJh7NeY59qDEJlJwEPcgwUPGoIb6ZEnwX
xsPmfHqFiHTOoq9SpJe3cyASV6d4h7k0kWSE++4qkwzq4AO7nAxARAeFwVuWz7Kl
xMRsUtq1twzQiZMOW9WV21cBZGq7CLimcI1CPGCfvNxcf9MaAuzCbfV8NMubXRJH
3Q0v94AoMF1PbymVhnTD8HiNLj2DOGnsJyLVMfpQ9pJl+J0KDRXH2GG3r48Gepdj
FxP77CQ1YBNUB0NXgspBz5gnF44vuG1n5/CFzyM/abvg9hqWn35/UiL0eKF7I5X0
rHFxu2f+NIqCJCGivqA/w9BMdvIdG7RHDsNKQhgtCAvYI1EVJFNM3rBBu9BXjY2I
/K1IwA5Qi2shV9I0NwNY498Ree5VwEm7Pr0DSbHHhlcAZJepWamJcbxYW/iM/Wao
ZFTWYGwDO8zm/87jyi0zl8LvcIgDn2VOPlcbc4VlFeB1tBtEF/LL3AZWWabfcDyz
HPGG88VWcx1biwRTz+dAk8Qz1aAScpIE+e+DYkvKERRha0dnBYdX6BGOIiRU84LC
dfCdNeSh4JGL1QetxbjnbTV9R23ueQh70fcODbZH8oygtrSv2iXSBuBh7KhEYcko
6XSSTlIAoj573wxs6cR/tQsEU8o6VH/6Hq/uozDhvLrzyss+O/TKu2fLJVZZwu6g
bemuXPeFe4/fNwLGEjXfuP0kLEbkjKNpNdSG36iHwjzWoIDzBvYk3w4f1TjFIth6
xXD20K5wOFCWTQXKLj8PMfT4xm8iw3Yh2zD/LZ7PThwPVvNicmASzBTsuw1+9Imx
o+rHAU/burEqfwGkoUm9wqq8LWol+SSTztADQc1j5yg69xvLi2aMRhzCkInA/ZFd
+07yEM5S03LdVGEII9F81AS06GlTxSs5/ZUR3h2ZbvqL3G7awwVuU3Qb1e3BEjJ6
AIy88c7/Euyl+t50Y9dHwt7UlWkc9/BFPii1py85mcqfDL6rICvIvLA8fMMhGlAd
Q5evgeIMUVy+U8MJ+DMhB07pmk5ZQvGA5FqZrCiQgtj6vMSrdzm4zSn7xVmQ/+S4
jZs7NswV7jl4skupn3g8u6v3cLl0zwdD8yVgdQh7oiDyXWR/jJA7H9+wseqa5RJM
+yjXnm/owmufL7z45rt9AFQfJPL+1g5bE/b32A5VsqM3vTbi/ZCmHyCUQPTm6fjL
oWcIFOQaEP0ySD74bq161NKpjCNcHbzG51fXAQ9OwYTLN/8KNTjxQOKhQDsPgE6u
YpteDvju50cQ64p6C+1+1UwNF61SYw/1UrOuCrhrvYdQXpRakICwhA7U0FYh16kd
HcABs3XcMFJAS7O93luYp/bjIYf/A1wqTWDs3rGxE+9vbGzD9QFUNRmC9bnbhjXE
8FmVlZG3LCi7I7CpzTF3EtRT+9mc16pdgzA98BOQyTifCk/15Qcz86da+HDZISbr
fBaqlPd277GnX76CkUHvPYVGs5Rh6/sz3kRVzPeQEe4ELlEPgyQsyLyoP5mtTL2v
2gVX0Gg4fDbCsMgfTrmKt68a/GKB92cxHgI6iZ0SYnen8vzuXZbLo94m41tBHqug
rzSmomGpuxG/Mb+lCXVHAdjbL8U7uZSprKAb5lm448//2/Ujifke0ayjYl2LcK3/
wj2A0jSF4SmZt3dZSnR4YSU7C4u2SWr4CkWKH33MLTc4/S0xYzqr1Ox8WfqUABh8
+4XeHWfiGQ2r1vTrt7A2rPQMwsNwphwsBShj3HEQagGYDDpMfsQBmcYu+ErMszM2
oih3713X87yj2iGhNwm4pkD/y18G+YLFWN9I/CbJSb6SFy+eGf/PxymTiPpvkndD
NZS8v8ntsEnZeGqEylOcH2VXEFPZJDuxtYVdXlodjKaP6H5MTpVNGQgArnMNmaZT
9JBFJqqW0N4r9BmYuS3An71gCdbdsf02Zw6OmbPK6x3RY4ClNKujgqANXdD/gS5P
zE0vqgbUI+mb5KPWUcvKGk2RphDki20BSfkjswuPSz8WXg4rL6Lx6Zdb3i7qckPV
IBVSaXRQBbKM3xjj++VNABhOR7MlSsFvH+3c0uNlr1J2vJAV8zh1wYWbD0t/5BkU
gbXqip+rS1cTgNh01GprndwuMVzrl4ESyDwa/Rz1kiixXqC0WNWU3BX09Ki6VKr9
pt1clOmsOyVsj3bHvZHI4w8xmIO17vBHpbw/0Pr+ufnmSbk43vrBB0NdPnu606Z2
8LDnbVriJwzjvBfhccd0+/14krud/khgpDHEMFQAll9E4unZQBDx1jzJlF8j5jrX
6ctQHF5m6xqUx2EJKbdkZAxKtu0nrqWBqIqzTyOoBQSDlB9A2rVRMhQvCgDR0LpG
1zUmo1S1AUVtniIfGDOYgjWUdSr3y2N5fho9oHr+MRgvG9fP3f9BKKwdIklbi8Of
FIgjg49B//8Ob7qV5DSgabxCEs9L0C1YnLX9eMWMZeoB+hjvi1AD/SyCyUx5iO6f
/DoIzImyG92+jIUNkC3cqYfMfQ7VHSpjglPb/QwwXdzG9RTaJ78Bei/1lU8aipkU
dTaoF0y+AWFif+RwcZ/48r+40+27cSlMlT21RJHCY6c+G8s1Om/+oUg52MKz4KYx
R5Jy7f2Mn0GZC0FX333ikNlgWXTkc9NKoGKZsbfIlfgk6vwEFzfiVVtlAE5VcOHg
sZ7s5D71d0D+471WIflyCd3HoUDR1PrnE3W6reNSkXNqd3ISKfC/Z99bsjTobe8q
6djVrYsFWFWf1O4Sa3DTGOgD9GSjOMqE9vb7U0Ek5p2kTiJ+l4kxGHDdbR7NIrEA
HQ3S/M/k4KWgacLuxl8xjP77W+O3GUVOTznkFWzr/VAvb1vAOgIOpQjo3/YNWzb9
oWMMb42FnBQhqaHNmsPK1xHy86gxZkpk/1NmkAK5UZ/qvwdQ+ENiLr0ydnHoI5Ml
MSgHOpBtHvHaiIitnr8GTVUtADXRlkI16E5WZUQoJLvAQ6u3OrmwU+QXO9Ll8aI8
mJPTJepzr9ET0zel5devLMyPpTmUu0y7JwPs38g6djjT06rtRhL9gt3O45TXENTe
XFSUuZ/RAcj04lDR44vzhiIdSIzEod5gluqaY5NWTTL0h4040aRd8bZefvzkIPZp
NiqSU1x68LQwI2WjhVzAoLe2sVKEK/mwoD4y8rIyWM5igS+SfmGK23dO0kAjMLug
fmlfuseZS83bxLGf8dEx+gi5staD6jf9ODSAPpkqzN0MNZbhRzPvp7wjkl9odnan
M8U5iWnEALxOfHZISIPQlJtKScK88tJCI6+kTGDnQEsruS7n16zDX2+SQBUT01jh
Pv4Q5DBudBJt5t6wp9kQxGdhEqNCRScVeq0QZARUKb9cAjIDFrzkvfRh6JvcoXAx
2Jt5VF1dfNkZnM1PDzvyATcn1nySm3wNTK7dIatfFpOCr7ds+makoiScBWzXOUm/
48hDGB5s/tkavtptpVRKf9QCn+6Db+NklkHQ/ddza7mG73eA1RpCGLBvt9UYTNTd
wyiTdEA2z6e0qt62maJRcuCSv5ye0Uc7ViHch6eQe4OfxI1gkj0ordHmwPuQxW6a
SyJWr4qfMEzGmE5OjF7YZsROycu9j/AY96IPs6h2YDWNkULpaMP4h5jQRglFPyi5
SdXWPvhmKECIeu5IoZh/bSQVfoWvRcF54O3OZ5wldNKwjEglGOxrUa3bJMOenA5R
DMM+TrsPx1Aq7iU8hI8w3ZxvCnLRHDGUBxvK/zhJE1TqBlAJ9LlEvQUySCQCABkp
dpyieQ+iZbfa48IpCPQUmeUbINfIzxTtY1ab66d3zfijj8EPxwo69+M/SY1bh/La
XSQuokJWViEH6Ww9Abw2yOIQV0GhHRa9EsiTwrRbUFoGmGlwSQjrxXQAl7XHFuQb
SSUS8wZl3lh1BQLPg7AzeIX4u+p+TL8GHonWuNnUtARON2CNpd9+DmtP40jrtpLi
YRGmrIyWxSlbAtFRZRYWYIUtwd/MD2K8U+r0Xi4Va854LknVw9HJotXeB4phWk5m
nLnKxWCDMevWACkQKOeteUriZ7XnvLjM4JauE23xg71t73T5MiHfVgI3RemxYMCy
4MQ/kVoMFk7k6Y4fVlQ/yljn2IXZ9Pzs7243WkYeE/tX9TQEG3wvyslEULbtVWr7
g4QafRM9LLb9uYijw5UYHGwlwEVDZZAbUIrkc5V9TP+tjyz/kuV6ac8UBOdj+3h3
mFnFPto1jHdgcT5sUBKwhgLDETWlrwiztivGB+UYDH6f+EiIg1LS+0GFVePmzE0x
+2pzlm2QgR2buzA/Ezc20Tz1ckVMGfDkNvTemWr+hcdtRy+GjWSUu7I5mhopCfEs
YW28AZj3JrA14/zTnBwmJxtGlDoFGQVk1CO8x/8AMqrxu+mrISQVnoJHpS7kUCaG
wrr/EdWNV67i/Q1u1sJgp8KztKIP1+kvqfJot6KnUvksVOhU+BbwJzsaUSA9pxsX
iQmHqiObPFsUBgTvU9mJJaSDug5D9UB0tw/zaXpwaa30I7C+ZBLlxY2JmyerNF/G
NeYJSMWbd7oBn5VaqunCvNo0OC9SGhEehDXiR8TFxpXCsyru/Aaz1lN8pPnxttbr
S4UGD0YxKwJzSbrLLQlL5F9A/VfHvsBAMy7XZUHm9yCgQyTRCwmubwHVmVNJPc9u
WVEzGPKfuYAQAWCLxYDIVDrmJEIhV7yvBI4i/reF01FI3HEH0hWggfy6Cp3N1Yti
steOgvgkzducP8TUJp9qQPw/xaxP9LONsf/dRJGCPmsZ/n0+22C/Nke697WrnQup
DikgvbqWOFKrHPDsKKC4YHeD6MfBYhhTBdZ+qbmPU+O421e8UfnSifqzo6DlDSQj
vt5wbJVxzl+UyAZumWQCsp8n4fHYSavU4jqGZOZKxN+pg7pzyG0S9xJrNppkEN27
uoOA4wVvVoM2XR8G0UWjYznkHwQMXj9Q/SYJewG43CqeqHsMH+f3ffgZdsb3bPOA
WxNN7ex6n54OXNpZ1mHjKAGE0x/d8kBxxXIP7hiyhwc9IZFsbI2gU9KWW4mCz7jA
df7s6Z/PcE4f0jaTeDQM3Rnvw8EfyHGcTabqQJLrcT3fdpqaSc/zstFc7I9KlQwe
6J/v2oKhZOhOY2TVkgdOeiCdghpxx8WKzojTir/EXc6sp6iYl9E4v4lO2bnUJK8b
fpFsIxrZL7XS85na72CdDxpq9h9IdY0BhF8U3zPnf6YdzeyIj3yRReaQF9kv/Yg4
V9DcNTvdAmkCwttdEBLLzL8limddQs5jjaGSTLVGkluBQ+mDjcDOteU7EW9d1v6u
QIcWdjtj7K6FVk8SI2W784Y3PeEZrl4fdADCV0tTkfWcAbkrSUmuKercyz9XclOl
1X26dCB667NqOTBOXMsa6VT2yRSkRjp93zmUi3oJkXmuyjjePsjz9zeMRJJXDZr7
5cgdfKc8OQOOlGcwNIHCCU4I1p9/BUB2vN/5T2SiwnSGEcWZ5mKh8mvQ0kcsKtAt
J1xYAVXeVM5DMW3GqXR3yUWUSUVbGyMBqwukYULVcp4hxYdBf7EwtCsy/Pvt/PVt
MU9P1wTz7k/EvhIaZEE5yP1O4qwMDRo07USMD6QA7g4l1UolYILlL5enhJCLXs6w
CdrS3Fv0Kytcm53b0nk7DS5soVR5jJDxl3FV8Jtbt3i6iuaM+cdQ+JPXvegjKuYd
XNwdROaB1NuGfOAhLhYbsHCv0JPl2pEdUCgfnJ/EYqqZKJ+spSsLkghxGH+xIrWE
X5cMJJK8F3A2Hb4vclEVrsB7pw23Ghf3Lb2+VDcLdlJOSWKvWvWem71AndDQFNbe
nfxE6byJM+hSbeSEaTt+KW1Svm44OUET4VgKXSFFk9I2PxsvNFebiYcdU36YNfhu
Q7l9LuLMI+oXJ/ZJBesEc+MHi7NMpaDDI1txurqnK7fcXxPAuf8vH8SWyQERGyK4
yNMo3tOKd67ES0o7hs23BFx4rbP5+Q8GjrDC4Vm6mmfr8XE4ccLzulxLWOaSdiS1
1f7CYDD7HKbfbv15UxssQa0Kn0F+VcpMtcAeaiU0syJ1DPIZz1kg6I+dAJNLsHsY
FV1mE2alcTFfJwsy7d0t5w7CwewDWkTM+uurrT3S1AMMMCqNzc+mmKHYfPj7t7yJ
itHkKtjR8W+7S5rtw9iuLi/KKCnjI9bys6Zhqnk5567txuMw6smMtXaOjh3snBiP
S2MaAquOh9KNNpIr3cAqlg26Q1RvfQM5vzszRemltanNmg2kFjQHkn2WNFHJNRLj
sdch/EvdlW8P2NdneMhdGZw0NcJIcYKv1/cZtbaeI8yyFJZIO5yVX0KZ2NFLBrdW
CHHmsGXEnG8IHCVhkqxnG/2KthTW1SLXYoKZCKmr12MuCy9ne5eEx377pUsFFTXY
s0au3W/KDPl2Aas2n/K7Hip48YoSb2svPX3j9gq+ojUcKu8/uhbgB6a66rTe25xN
4gErESXrJo00BB2oPBPzszyksRHMS+fmt1F2wZNdvzkRvzDBNFS5gYBhKvEyI2j4
pFZ86W0j/e2nLUGDP+EebrCb67RIjrB16s1bYQzhT/IiyfanJaYJ1ol10s73W4tb
SSxbNiO9MCtSmb0v2v4SHGX3bLm7zlBjkt1aMqK61OS9Cl6ZMb0jRd7jQnI8r+VG
4XCnHQE7nx2kH+m3ycl7zsquV5y0lDrMv6vTAnZEkPpFQLvhEMGWX++SN4RTqSv5
C1k5/RU2bbDUP5r6ALIqs8EHiksfnuUBNzNogSVNyBnc/onoz+WsFrOLT6I66cUI
qEN83l8KV6r1EBqWF8LdI/hcY9j46XuCwKnrZk0yQcKmhuCLEN1nyzxSJDB3kIzS
4MpDfXX0DgeECxp2nmNfzbdW9XtHVPuIf0hXSdyHs/jpkcWD5OwgY0TbQ5zFQuwr
4Xgvfhikb9nUJc8jv2SB/o0KdUTa0q8GhPyl4ev4+tOmkdA7WUo/cWp7j35DSEzZ
vIWPk/0csgvGNc3lWuEAGieONEECPy5BJ+303T/+wrFIR3aP2nUdRE4UjyHYay4o
g7AQKMIrRWIbDFkZ7IAAbMhPaZYypIhlJrzPhVKWcodOJFhlBszwrq6W4o/DZNxB
ljDB6RUHdUmWCfUmU+1frBlH10XCeg3y9odksfadb4egudJdPavJtyunw3/qw0ah
VzK5V2Ok7FTfovy4WBZwrnIoq5Cw6v4Dhp6nWhIQ79lxQAkK+T4I3DKhCT83yNmF
7Rksiq6VyjlOSZZ5NckN1jId0pd4dhiw5JQ0UXTpgFbbptPYDqnFxGhvSyRzsVRM
abpbOiAn2acrZZJ8Yj3HuZ3C3lKlFhPcpaCFRoZB5UoVVqENP1tsPEGwxXkud38I
myyYCtR/twmlMzQSXbXs41cFLlqb0CgXAr3SciQRxSg8Os1ACyhJis8S/PIwRNMl
ZX1moWSojpIwB8gpafvQbyLkQuwPM9ZHpFOTHKCtZtl3ZFHVvGSZTQCb2XlOLMUT
XJNG+RrKCOFfd+LAbvWYwXJZ1/I2A5hWBxJvitYJBCZO79Z0WRl+KOCE/trm4FJb
Cp4kvOsHmZFlVb/zdMTo/C17RDWiKXpzH0AfgnfSMyDsoerRgWZht2RGH3V5SXb+
OGaQiCEQ++GacHo8A3fIY7G7lg58HISsiQZ+hbEf9M0eq6YtPfycz1cRK2ErP/cI
I7F8uk7w2UyrG3Py3i6XHeRqaYZtmw86ejnH4FE5VJhE/VOgry4ckzyXmyPFu6Og
/qwTFgAa+Vmxac23UlFq1c2sGDUJAzIB1QMNbvrqi9lb+VqYuopjmENLuP4kESDy
mMFq7nTRUfCOI0x0a7BwqeF0Q0Bxap81/WgnUrvW68B3GRfUMmJ7/Nv3Dxghx1w1
VBsHLPYPVYntE/jbos1SyMMXtH/FLeAaRfD80n+eAIHXjTYWhzzf2OBkuBmQXMTj
no44owAGpDq85vwHT7g/ZSzcY26eg5DM+KrjC91cknW41IZB4Z4+kxBCJs5M1Uht
hnMctKvOOt/qHuXkx7GLDJSk4EPuDBpYzgoH0SgJTRccmB494VuvJtbeqzZ1QfGj
bGyRCI1oiNtbPeaJP2Nt+/4Fox4fUYCjpLZfPRUy4rfcZlzlEj0bxOUGQvvk+vgb
OBCYdiLSmTpalcb3IJfdBQBBOdwt3XTbnuFix4JpAC+rymklGG0sIXxsmf0bkt7r
f3irprMzeBRH9PXK0zHlKix+4n6J6hjG3k9MzGiNRk0f+FPbPCnMBA+12nFtPm4K
e96AGUIqWAI5wvHFn6ywo583hJsYuOdO432eNoi0u9Nk9kTmTNFTHKaULYrV9lI/
Ewu0V0hEdvNX+R113MdtDWGsjwXHntGQDCYHTwHqWycF4mPzxeJlbyrsb6rGzNgJ
90p5RmA4fnd9BtVhedzpP5GUqwn+EvLkHvX+AOrjq2Y+Qw5t6Ox0YpyKMWBKct+j
5O8mf7R51gDNMZIWgn0nFedjKXlMpFiguA7GodkqulltXjAxpAjKWjEn6+g5HlbR
3la5Jzlm4OMmzP7KSuebY6/5DMnMGFXqJYhbVUigOVRXKrjwFGAZbjv2sstwzu9S
n32V9JsZ8fbV7REe0QpI+K3lAa5QECPFvkPBw5JHjAvh5nzRyHjtJK/7suhSfeMV
iQiD/xk4MhAwWvKhibvEbFd5o9LBPUnstZGE/eYzdojuvSSd7Z22XG4Oh7YZD/nR
90g7CxhrT1CHNV3nH0o7b6VsIcl2Xf5HRFQmHQiRKrccA1s+q6oMXYB4iwUurrFQ
4SuIMsYGEF2KibHW3MOxz5jC5/Zct+pPrt8lACuhaH7iD7v3GfTxwOQxKfnmfWPu
PykHm0hMa/K02Igv17SlvP4pD7LSM7v4om3JkMYI4XV6MRvMgspQQ8+mLa7GrtWl
DXRLgJfmEoIQ8AnwR7yV3jop4AVEJjhB1wXv77P/1pFlSX2koz5lbwzrh+ntxmx/
VGct/+ZAmJBM7OyGErQGDj13QAzWPFzAnXhSy170C67zbKUuwxopm4chGYyeCpao
9dpuiyB2+G5AGII4bYYUKCqzvmyAJ9bFqrG5kXkbCkdB6ajfFPIzrtM5yJtOg0OR
ThKQG/AGfliqzIMTAg7iJ1Z0XEnsyBJBt1Gvi9g8/vL9eg83UVhpGhlvAIJRNsci
GNk1vUk8GYC6H9Wn8/nSewY1jpuiR0AX4kX6Hmm5yFpCbODEQqJDKxufTThKH4Yj
Q11JQl8UmoqlXZzcWRTV5cSmOEY9nYRP3PicflDMaw68F+/kdpNARSVeAMuJlXBL
0TCisPIbQzM6RU6704n3grdWFOeStiR0wUXJ5Hp0xHC50hz6uY2DxDojNMny2196
VMvjB/0edx9LZlF7+GnORkLFqUZfNzinVza7tlRcKZAcrfmN2ezLjbStQraWWI/w
4r2uoDJLTKWGCWJR90No92b5DX994irQQwucThlulG5wAXr1RMEQDE994J5oPFlC
V5AV2eDEuTRUdv7HuRgwI+YZLC2IvEQ4FNldUBAGI6PW8AL4FM8b4vawP4K6cna+
dVKsnmeWbp+gfuRo9VCOM50xsyBPeCM8itGnnBpCvY8bSViEg87Q9gKWK/i9DJDI
9bxoNvGINEHfE4+xbp0Q/kKvcL5xK9nft/a923MjgIozgdn7UXO9C49luxcSKp07
I/gxwYg0zJ4tex2rj+zRv4EfS9jlopm6zlzY9m3rlszZorqzOfQS2Y2z/otSrwrw
3clwORNB8b4SEMKYb1fI+Z/gPgxqalWw/5fIyeLWCQvLomldv2bCSFtX3E6paQlK
mRJtx0m2p0hSN/4AUt3UkSN0/ytvfqWycYVg23Ewo7+3xmwr8GPaZenhRJqtbt+g
xwTpdGGS6W4yqREE8I9DRw0EsMD55HFow7XIX0FYoO3lwKs6s395r/iVFC7xYLp0
WioUVKEdMwEVaslU1BCAHEoeRVfr/0nev8PBwqHf/aMYuPoLlu/RmjeG+KczWHun
0t0LTWcNU1S+tAK2eZbNFRvOSjDD6CYk+bV7ZELkP1AgNCVfz5LY9NdU2x017VLE
4B8i6bO2VPqkEVdKd0X/tTzCoXwXXEiiEJmXsK5WlJ83dHF0CY6rp4Wr2gMrRLuC
1mpFfmOsU1zbjKboGHpkNePUh1nHGv9NmKx6y9mMg5TvKVUL24r+pP9X9vr7vOlf
xHvA7ucUKlCjBfJ253GL6Pcm16i5fPXOrQ3b7T4d2JMMiJJNJiWDdPu1cgCmgOG7
M66d0bNdhCboZ2qN5dHWSoa2C5RD+ey8UvAdvl7Ep6sQbyu19AhOl2I95NYKs88P
3101hJ5Rfsud/ytOFWV45pTMlCxzPopLbII1ZFIuGVbe9Sur4uxCMgnnu35v1uD7
jlDz3U4ywvKMcquFrEWHX3j+TKKb4UXt3ipvX+BaBejUJcfhCauLX4rrXPwXO30s
XdOf+iVscZuwO+RjQMnNLeVi/dj6ER8uY4Z7bcUufTQc9g+C+ez0O+7ADsYT+dQF
DUxJjMk/rFAh4dO+COb1B82cU9yyo+J/KpCXUV0g1tLfG8OdcK1Vi65cuHr13B8k
TcXBElBS/5Dp9Fd7+VTqkDTqMJ9rBLHKLujecyu5MteCT/ZU9bM64Oqef3eNkeBE
K821d1zXdwmSCPgVapt1ho3trRQWvntkf7NAMFUm1kp2Z4fh4VkmMqaNf+x9BDzx
cJN99hSTdF8wvaVa9L0g8f12imdBZYGC3I4ZG1JFUa6nStu71J1BLg4Eh7IsdfHV
OaZbtX8i/zrFiFo1utLUEleiAubw3rAWhe2tydTpl0+E/kAgrDHfUvwIGOfVHZjq
87EGriGQCvZeO+1fpxhlkmuSERSVR77WPaxaduca9LvDSWxY+ewCqfzDBFFA1334
qHCsMfu3UADYoGU1wL3GW3cYdFAndOllZzUDCJz6ydSYzlDTEH6N5Ky0mlRLVdft
g1I00TTVhgdn8NT4dX0v7e1Pwl+p4cK+SJmkOWdQuB6b/g4VK0L7y+xnKBQp1HVT
Wa4nrRXr/HpZjGjpfPjG7mNf3Spf6ULyIldJw9rt8Epz9+blUex+e2VTWuWUIuOi
ZJWCuY6PU4W9ZG103dF+A0O/hsIjWuUR+RpsTXD8fsNyYXhni7thQQJVqQ/rKujp
uRjijVy1wxGs2glA+YU3YAZPVuwg3sdCSGuJUBF+AX/5R1NOdIYWl9nAi2x0qnwt
xz3ghy2uww5l9C8oscP1p29lgP5i6pdHP6AXMbZTt6o0h9jH4oxDnOIq/O70GoYr
rb8ETdRFas221TdxxJR+c0UbOzVcXqVX1A189vHsSYO/eiWbbZaMwlUd3pnNVWwd
TsXcyhkn4kZODXUjmwJI+kKUPVuWmUJP+Oqjpr5ZlLJD2/9a8jwI7qL5diYGbIWX
g9nnHTbXi41B7YyvDu47DxeIdwUmtsuNl8rRKwgpG4JJ2g+UBn+O7wXMCkg6I50A
BCaw76to4YjeLuWrrzaoJw1U/QdC0Ybf3sMm7gau0xQ2viNU53nEohUJqUh5YGWh
KA26C76o52HGYVmxJ++z85+QFM3PNbkScw5/Cy3SuiFw7Ri6myZQXWMnOr8/8mmO
L6003iSVp+BWre2K1iXdzDdJ3a2V0+MyTAyfzpkpXepRkallb8sn35yo1yFhQOw7
fPt33rjd06rjGJQyKLw+jqse+g2rgeMx7Odqo6NhPUo7XCYjEBfEcHtgtmpbTtwI
r8vCO6mxybtavBGiAbJI6p/JFKpI7DWuD6vdB8h2x5Kq/HLmK3COyovbx7V5u7/X
HCxNUsT7N0PsgJSUHjvzo23UE4eLqfLjeage7poYYpkZ049jt7z8HLSJ1ps009YD
HzQCL46eHBJdUnRIeK0UrIHC8dylYfX9EJ18FpRnmvCUKhvowBxKve7WlKBHFJcX
4fzkeNrIwnoxhBAwIBk8OMMjJPt3XoYCL2jtuktpOokRUI5eX7i2NjnXY0NZdINU
KQsUQrrvYVp4EQQa6pG1g5u67fEqfYkMRIHyFPLmfxQapO+jUdzCCXhHgsDcS1Z3
YTwycM92SrTcdF4Vo0U1m+/P+az2cAc19aeztU3RV999LO6SrmM8FqBsAnv94tTn
0MoXiMpUy3Mq3TvtN6dLDRKrnh6Zn1OmY41Kub8I5OQNOl2uBN5Qow5Jfa2UmkuR
fjyOvGMWXfLGdBG8ncnQ2dnXPbIO+gE6GGGS0esHX7zjBMAsewKbKDDFOj28dbGl
CpYfF5qZzLWuf+MW/Qp66uOme3pMj2YhcgS8gOoOS15sbkhcFgpxRPLOXgVShYt/
3SkXlT4WXs3KG0e6c1iI1E3EDCNUCIVdkZOM/PVvAyR7DQ3oXhkj0DPxbr5dj6S/
Daq2Cqwu6qoI5Kdjcgcv2l/17brbgbIP34SrKORuE3+1eZnWq1jEHWfOBsFfWjJM
9s5AapCqvGT8BPkSaYY+xFd+KHPhtfXSQM3HkLCLMtQ0RFmXLtZH6Gj7Kj/uRMb9
IPK/6kk7Fnwf2ofAE+idDB7JOOIXML+OljvEAbExMEsAvzkimcqp6ZRKG4n9xsPT
dBsgf/J3YnGZKcNXthlGwiId7dvCWaqruJULwUlg6q+gnBXFwmtVCCeu48YTLoRR
kp0e9K2zwQiVvYbkZWjSYiDgAmwAATuXLQSIdyKy0uLhqeh3wKCRwAtOuGSbjlQT
gNpwZV1eK09qw6aDe2WZFZWcQWfVWE33Pm1lM/rNUxm+h2ywC2f8A4estqQKp8wv
VnLfNFpD2ozxuwshD8i5qpSp2k7VhHqgTBPl4PFTW7JWKjuoAlquZIX/g5RFsgWf
LTn4aWswmJMetZ70cv9TR5dJgYs1OU9NlOwwEaZ3pu6q+GD0r4x9G52lkbzqpojB
8+3h9ZSMK8wMlnRxeafUM5Trb5lIH3Q7jX8BBok2tycS80kABZ2dHyJhm3A5w1xB
MlBc6gZdfZl1UGJauEh6Kgbj+znliD73LdZmX+AJ5zAeRBX68J6RUTIzdb6suZI1
+Jr1FJmoYCtckELwbe+K8HzgcfRNhFQCY5vnI4AFFLM5D6/BCSZrRvgIIxc5Kcvn
tN7O2YCMMK+JGtMwoyBBLIJFQ5fi5Y1cj1KwZcV1dk5fLVSuoZYQ4uFOFQ7P4X5m
ROpFbjHFLJxlHu3cWhhVeoaCfLmIPzDXAsG1Phu6m8/pBqZ6gts43BgGDy+TvoPP
CHAyGxC8W6CDIe0SoasmfdcipuSE/+cTGuMRhe864A8viJSnIbyCSX5teC1yIFVl
oTZE9dYzQ7erW0pPj3ft0UgKv0JlMu9XQH3pAhTo6aUpAFVvoK3GglceDXn+tUQ8
rPGqHOitcnBFvjLCBNxqkA2tpA6S54+cE6S/Xmdk7Ub86lZwRmCt3Hli3XHZfm6V
zdOTsW2rwzo14XYfN/oDCjJDT2llNZQD4e+itlIVKpqXIP7FEnYzXhyitp4N0HXl
uYCxR6GeTw5Oqf0BZtyIyrUnw80MxGM0N9jzShDDR3Yl3muGPzMQj8PLqlHBSpqQ
FHxdxWDVja3NuhZME5kwGi1yxujANS280J6j8IVIXlpv86x9a2VDLIsBMNeF+LPK
3GFlUkGENCfLrHn2dHdjTQpElon/G91i65dWLu98t1NLnOeJvXADEiH9eUJPH/oz
5jYqNYu0NbnbfWlLYddXY6AF7iuisjK/VWiTVorljYpe7rULJdAqjTZaCHF9Zlgw
9ip5rkRvNcTLZnOnQkUJmoqbSK/LNtl9h3DOvNKdVmTRNqpdU8cOxOMupbsVkVzC
SQyM3+G1xgaFO0oQ0EF0G+vT6kskAKgnNcWjk6pZjxWn+GcvoDDy0okoifzhrGyL
uLceWefODx+Y1k5wIsZeIMs3nwCRjhdTljSMghj73NOQ9F3EJRKqXjRF1iC6u5yR
RNX1qc7Hu5vfwf8M2CbAubIc+sGF6atgA/TLkifm5BaQcPD0/QEjJk7dY982mZpf
wB2XDx+MrixYuNmVoDo1k1Gdg8ZnKntwSVwORT/1fRk/cMG1va8XyYOwrLldZPc5
lsevgkTCymAvT/hmES+d/rMdkQAk7/2f0WtP+xwW37NvveFh/MNAp1KLvzjpRiV4
DVR+oFsGGDs5NNMuQyeOGhmWCqXS0E55vJEvo0cylpNKamMshW5wHXJzMzM5EyOq
6SC4Cz3lj9SeomfEmlXpUYqHJucfXmO1R0MPa53w/iZKujYeWEausFP9HC2wO2OZ
6AAk85THPbfxau7l+uh0QE7Og9tVT7a/HaLWqsBu523wMkG+PCaSka2/ZmKCeSj9
k98o36C0UXvkejj9oC0mqc/G3Rjymbj1CLDcssdm3sPytskKfDiWwLHgdR2Ak2ca
/RdLmPR+5+Zk4VBVMFog/a6+0EweUg39vFunlMjI9S4246UijIHzMX6EqTCJH6L5
8xfneA1A61LVwbBACkIB1AnN+yD/EFz6SlaBBJiM4HOwoP7KaIbZUf/AzPFFT4DQ
emXIUFtCkBQLM0+HEnq2pLzHdxT9q4zbn0zaJfbHt+cbROj2Hqi+PqW2TC+UJnUM
gw0E9OV3PuiPqOuHWVLpGIY6mGwCWOLU0tKuGh6ddjIXJQdAlesPyrTDziDTsPMS
2i0dUG3RZqbDW3KvEh2sKEyJqJDlPg+yzceSIQRixWSIYFDFld0FZBumdOea9XUX
gdCAZXOA/UbRAfPHmCTRUULY/eA9EeDQTJzIoPTUYBCKCllk7p9m5mcRKqEB0egq
ceuGpgJsGCnANfxmiLuBIemDHgfoKwsv/BzoeQk6SM81xWfF3Up85V6SusmalOS1
VQsGi9CC8NE8hfPngqzwyLzRjx8v/lwJKBg3u8qK2jK2t1f6eXd5LKkvZBdX0lnL
ctjZ2IyKcLe7DjLdy8fdO76ET25dmPzTqr0mKjBKc+ckbZ7Sb10PB4IMxT57Sn7T
ic7I4fm8+OF5fTjsRqUp9oskRjFa8btOP60ZJu2o2bh7YdQvXW+MJ0c5ZawXmIZD
v0zQRX8qXIaVMNrKcn5PhzDZxvtORRhFFNrtqb/sExMAnGE/Npc9il95l43xqrQt
1NKXJBuHFVDKYkLIdbOr8kS3ISIifWicBvotbP+ulC1RGdfJASVtWrlXObUWi6JX
c1K0r8fylp6b33HxXfNd2DhnHoZZSOCLfq0q2vr81yP76ETZ2CbuApotpx8MCGAi
3lO1CAqxKJVejCeze1tQ264+o7mdkAd7hXngwl4yh3dXOSaIr7oRbpHpawqArfUw
ALRm1unmax54C2TupXGjwKKYmqsTX2wjAbxiyDnEK7WyGeFuaWO7OLbtoIWOe/R+
5vaELEObfJointkrIPOusgRErfjZlxY3oVBMCWlvI03FojNm8/SqqIk3Gv5fajVT
Jq68pSkMKO+OzfvVB9wtlnkjZOddL39wPObQ1CAqZ8nPU02sHMaFbAa7erihllcB
4NEa1w9oPA+klK3FpMhovgJlZgroVVlgjuL4s4K+SiQQkS5k/0Z3AMs10CaXXE3c
fYbvAHtqCvRD6f10ZSiJXBx4c4uXR5DuP4JBBU9eQk8NMpCiGGmrsAo6Y4K2rfwh
9xVphHjpS5UOPkx/VfbC292nrDdIdFUlZCrbl7tL3fUtCyQ3ucL29CH9+fmIjW6+
uIz6UkRmNWCTI1tQvQmkITqztV1iA8SOGknZ7G11cYt7BBPYcRkOX4lwg3wa7KGN
b3v4IvnYfY7xgfQWmwXp0UMk3K9vff0edVXXiqw+MFLnD8kpTSDVrwpJj4RG0aIP
8lKthjF323y/Au5vuY224BmT/n4TFbgdOwj+JP/JBB+KajIVKGhWHQ9GAxq23Yks
8jTeFowIe+Oeo7uslgjUpBGYhLICXGV36vS4SVOXeyYz389aAHcCtX1eHJRnskx+
jA+eFq5NykjATCdVv60h5u+LbE2S6yqfeE9lRVlbMS47gsdhD0nwR+M3K3bF4v6a
qk+80Obxt2pkz+g0FnJIomSFkChNN9oPsGv1NVYh1aa7HuxR/el5sHzi/k1OL4FD
TG4V8Vwk2rZ4UXPIuJFxbQ/OmzgWf6G9/qGmySZY+5SRMyNOwI5YEmbkT4PuI+wy
BZWsVGOyRPR+7zBmL39jkEN6gPF3DD2NqlH1AW8YGO/tEG8Llyjw4yUp4dPLfkWR
rUJX+lpkQa0PGv2R13ccZhJ4DTe7u4bclimRnMgpmBKzCKU6JkLy8YHB7YqYajOV
5K94BsY5zeILIoQPniaVYTCGbDeZpn55puHltT+X6HEPPnO4z8s8lCm+ztsw1cGJ
VmB/eKxcRZSsLFm+c11WgnnDL5roEWrkfsiDxjJvhxzNoLFLsSEmsRqrrfdtzw5a
Cmh9bJJWeQpv7ylzFPWxGc44iFqxuXkJuZmkdmrtSsTTPbzVjxFYseQL2Ei073M3
YRDXR3xr8P9SwrU8y2Wq17p2uYLdrW9GJ83CrKNw6cInUEJAU8OuBn2Vcqews5VY
4SKgqgdaIi0iG8m9MWgMK3Ir8HL7Jkt8AwsCHYoP/rf6yc/LewNQHuK3JW2BfFJZ
9QQ5NLzN7wd9fQAA+quIE9g0obsty/vZmcZfde8r/rUqc9K51skcchDz8P6ttdRl
/gi5JOteMHcwAfl+snFaM5MMY+ijA5Csx+lBTRHyUiXH3vbTlSlvueLG0oSanUEy
Ncwaj8K9YSrjLOWrFSNKR7YPsjW6D5y6huSsfwMb0hQI+Pbsnxa4idzk6IYQH08A
DGcbwDVHoK3GpOSbnWAWj6JtS+sC0xWs7xKdEKgOZT3jqQhWD3/74iiR/d6Wc0GQ
Hci5z+Q7/v/5XJnPnvaPR1+SvwJYQQgfwHld8DgpRj8zxvi/xtc+KmqsoxVs70tp
wY3/fKRNmvICYxaMV9AiXz90UaWBk3EaerDdpkSHjW/nbVBhVnXTUN23UQobm/uu
1KghI+4uqSOfm+QwUZTSqrSBgPX0vhFffdk/vV0jHbVNepanUMqBsGtAyfH+S888
kZlGVCJ9hwB8sUdJpYBgsZfMotaS3KO628s6fUdIsQV8Xvtk/4CrzBZGV3ryjPFt
EzX+Jz4MgRhozjwIQHeoLbQX1yRYC6CX8qK6Hzk43sP8RfvLqqqeGVmwIcvUlrkk
Zw3DIu5/86+DAOmesWEaP9DYPhrPaoxSLmZCz1TnYYbcIR9kGXOy9hsgtaQM4VtD
LaDNkfuZiAV1Y+T3DS6pLCX64iUxfEcSd4QUNADIxRvlOu42XLHDSJVHVCl0ZLmk
YFmeJtTlwG/PudR7kDCYWFZRDMZMjPTMKgAoIcWaCoayEKyOqoDX7lNW5osfqtbw
aVX16yZNlxXx0z0Q8jmoB132qRRxrHr5HqfNmYX1dLBKQ1K+CFERktRPoMmJ/Ciq
pC4Vqwk+PMNcrye7tlcOR/exsC02mf/QM4LODb+eamqybQw0RQco5RP+3ejK9ndg
kVr751A2IWe+YHnYv/eb+vletbCv92bBCMXrEXKxBRwugNGdZfLb7gkvRvoDmQoy
rZyIXqgtQPPJQh7WEHEOdd60m3pCxvZdOaMOpz7kjuzj/gGdB9M0gPSnDjSBvuC2
mxSh39gjpf8TXO9JW4cvHepYlt6o2SO8q4uR+ZBnhwNhLa2SZIpGPTTWhzYxYnm3
SRQ5b+gI90yjXtIq3jsfV7Fx45cvF5F8tiQRne2Qz+0OWfkald4v1BQApPFGCOFA
b9HG+d/szFFpdU5YvuAXS44OR6ZzkmJv7xA3ET1qiDuteinqVl8cOSm6YBoIBuII
iAj5xq5qmRoujmD4Igee0iqppRzHV/oVqagsBIBpWL8pt9gzs6wbLlHuxosDVKOe
RIQ3W4efBeB6L5WupT77Fe4DHHHQ/k/vWiZR5X2k8Zu7gH37O3eSo5ploFmRCAaN
YI7I8zdLnEGI0oM9iEI9Mxi10fCu0/hfgh2eJNjCZn3hDO3pPHRYoI+MU2/4870C
m6ppOxDGTIuv7lRhJKathAjcBqNZuf9d26JK5xy7t4vOf6U0oXhkv7JabiUy6lBg
PWQrq8aQPLRr+pKV7BMQ5CIXzgVS0MJf3ghdhk5pwntnw2Pv4GyltDeUzAT3q1Id
6hWRGETVqWuhhRX5ke1HzjU8ygGhsGKzjyw+7oS+66XzAb9JPVxY+e3ih3FCPcwN
fhuRQ9a2D1ajoYIICFXypgqRAKpS0grrIrpZQ6M7ejpW03eFF+HGYJBoKFDf8vyn
dMx1bQWd1eeFRTeFxFvS0J3sd8jMMWGIA1Q3rfgQPEzXYhDWB0JK2hUYhlUVJ3Hp
Eljlyk5o/HMa6qP3a1m6f0MWBgyizjXT36ZZSmu/kl4e+eAhuUQn9PEwaTO8nr60
in5F2gCKCPGEFLF+ePL98iQQ2kn1C7FTc0Ptfk+vOXA4UA4+fpyETmKi+cvr/jTQ
l8u1bLNtOqascrgGzaNQxXwJVBARCAC6/yuwDUuahQa3tzos4KvMGwOWhaYeEy6p
FcVc1vQdhNuW/VDKTNHyA3JKEapz3zrAsNg+EY/E0HSz+coVI4chcgQqe66Qqp03
nuQAqhgkjhwznCXBLXZw3vyAQ1KzbAt7NIkfq8M7W2pnwOUTTEBNkxcfu+3t60Wp
0qMEmPuNdHzuu/OlJnYuAfulGchTbAF+FexDCNg787RuX6FkQ13W/dwFAvxNSglu
Rw0TW7+O+az4024MS+J7BYic1RiWZLQJLRKEMWRE9GcmqzksC9z9EjCoegN0/x7T
/9XQ7AAbX426QBt6Swg/V+spe7rflEZK19rxXED27Ef8LT/fhqmY3WRlQ4+jrP4s
Jb2SmnUsU7/okx08JG4PwDA1re6XoyeABVNhpWpimPSHx9R3QtcnEYPNsS/3YVLs
QywTN6FkSVFstsdnt7qEqyK4hKmi/MFHyJlJmIppdvizuP95sd3VBGVmjJ1I662l
zwPDBbWomgCnLQACpK96xV/+lLHjxexvELB4xaOUr6odfw3nmIt3V/7IUJizK5D7
VQWG3WUIbxq943fdD20UMzVi3WSa1sVAc6QVg0vBdrQOjHQDaPFgoL4nrNRutqFE
9Z0c6Ex0CMmi5RhS2Ro5J3Sni3MKB92m/3eY7xVZ8rTVVXZBXsJmiGbyvrcZ81b6
WdYYkdLEeK3J3wM9DVRFntgdUkpB8ZRwfzziKefU5UqPJfkJGJDPNBRuL5m0nqKa
f6uA97UlMNGnli+5zJdJg2o4rat6GSG4m4ui+aRpeJveociwsTrR+NVJ9RjRpcH2
b1o5oP4chh0xeXkPfGm8IuOoWai0uSUE+i6hXOokUDbvoR5iTpeAGxnVx6wy1V7Q
CFzlo+dk1O6HOCPIVAoNNyCK9IirUOzznDeRgpsbukCe5jgS/ikGPziQaGAZe3n4
8+rKc+okeJ6RzB4FIfZjDK17HmRoh2PfcFx9MdbJgnK0WdVFOPOy0VqqWQOP8bIE
ZvGDxXeC7yT3tvY8j31M6uGDeOxTh7SSkF1OxyO5lD/7iEFb/bsc4fyWhEL9R1Bb
duTh3KfdgxJ70LnAhAJhuDZJeTOW1IETP3b/bJOhGMnmYI814+gzwu01lxdOHXYG
7k1/JhPHI7wcNaUx/GI7VN1EgdLXMZ3mCzEUkhAAW//shMfl50ZGpVGhEP6T2Phd
zFCotIRHuCsiF0gfxyXmJoo1sS3koLNtwwDKhOlqiPNNYobLBXTayWdY2OYmalct
WItpfgmH9knXG4hmZog1zs4I5uGR28fGYejmr9D0NCESUpfj9oeQ2x2TTVb0kW5i
86396V2dwH+1SJQ8HbX4Wx1prNxI7926mxVNMjMynuaGOVpRYMrnmuqY5WwZmiR8
enc+f/kQZa20V60oOgBTI1kkFDsj2PIY5KAnpdJqOORMAnsCgGSZx1YmJYfg4bgj
sB6ZGBSVFt0wg5Mmt4Ved+5eVdpuc5wUZvPjTz60E85aMC8Z+5wtDX9UPXgHvvcX
hTA4nSN2e8D2vGG5HwjHjURqNNiJIiZWcPud4ioeboVnf0JlCN2fkkWda60/jZc7
XOEltsFHky3eoyben2qV9diX0kXkbJcJz2tMstVNHtoDQzAq+iGWLQFerS3ufie6
5ph529sTTGh6CGmLWbt4t9YhSxCU0i+mXyCh8m6kmWJrhm23XeBH25dKilrsakY5
pRofn2W3TsiWDXwEZ2wTKUkjM0zetFMvTQzmhiZfnfB3HCnFkIRlkSRxuNUBTGkD
QvX73BQt9vw1zPolkIgoFS518qR+DksYz66HikUKi/xeES/b6wYRCxHj2FE1TBwg
6EenoA87dUSjT676vmzFpAEBj5x0SsmnsRLUkRcvid3PPsBWnSbPed/e/T8zmnv6
RIfRxsbzmxY53tra5HT9Z13j5Ap2CfZgq6MrPwTRH9MV8lDJSM0d9rrTqyPaZQjO
3WTp5sf3kP9FQ71G47MQcMFVKOrOjVnyPqQCQ+6Ep1907ihSkH2sRyCkNgBH+KjX
DWODP4nbxoV8+PcG8uoCNMvBIK58r2JWLMgUzJuu2kPklOKdCDdF4k7rasRZ8qCt
tqcMLq+pSvtVUVyrhHAjFInQPXtt9ntDAKc/5ywTsB499GXvMf2tzDRsbugP/4Lc
m94XRCe3pTdk3/T4ugQXRFGJBAeZrA4gKpq4L7LWlLvygV+MMNc6B1qWZOa6UNp/
mQYzujPyd+X74ER6YyKMbLrJ9ntSK+/xGa5P4g0S0j+rJww3rxtbIVsF42+tOxDM
7FeTQmvcla9C+aKAZXHoU2yRTeRuQx0h5EilsUImYUnkWtG9qhdOL4wI47w1PU5Z
28ubRtLY0DR1coFfZLwAWhtWYdVckwyudsX/XOHY7An6wclrLZe4z0QcHp6BOCjs
e2ZkEbRiIZEMNcypcdHTgnMNzfR+bgeECsBWDCGVSFTJOnOUZuwH7U93wg3VexIJ
UG94v97v+H15Xd7VSz8Ja+1nbSYrBvCV3v88E/XvsuDzXJBVw63HzhYFdIvN72rj
jh+zH9wc9ueMDGkfumMgIT/YKLO5do0bjgMLpCEdOijIAl+6lZ5cz9ET+EhIKmu+
+3TxGp8x6XMPIxBVlDQxlmEcTXQxG39wgGT+PZOom+FYuBYoS6jEgAw8kc2PxI4I
kO9J9j2RyV0ZvNkKqVPRAvT/EoYCSdsMVHIM1oju6fiU3baMwnc5hV4qTSPZ/E9f
79rbAi8Lhs97DfORsU1rnX7qGFUMo9gE1/epy5d8fdrmUnnS5n1QWFQaEMu6aHMU
bVjqNFwY1cFAn/FgTZjZUVYDn+QjIpMAdecmSXyH27fQx9nHetKeR5c198+EZzNE
Bi940LhvFnlAiy+Y/9PBwS4/CBAbIWpFHDIrxFMnd/xtJDPQ5j9yre4FFYHdRmWB
9KyAsDYusdX1jTmjriRQPpPIfQjmfmafkaAwkc7reUZdgjeCYOjDJVUkNPq34Qvi
6JtLosd9rnH9POIAF2Vxn8JUmFaMzj9+u14izFMVqrHI6UiTZcG5km/f9k5p3shC
vL3fRsnetknRFKvPxZKHh2g7lvFyuU/JejXguZ0wPfv/3DasRR7N3hWByhXEWJFc
zFYYi4m5v8R7JwUBX7nMo7em5MRcJ3anK3YbewaCaKONmqK9vPrmudWC4szJNNYQ
nmJaGcTFkvuHywtoSbK0GyCjrtC/tUwEUXokoCjvWLsF4WeOxZt4bOlmABkGftGx
xrWG9X3d+v7WX5tcab6UAVrSTTU9uHDD6W5Yd15lg64MpqzZTsmVp93NLd82vopV
In9d58qyjRW57a6N15D9LdGFCtz+tDPx3DA9GGm8bxC0ro35dNhJ+bk9awol+kwo
MXBAqlTbBJ/LPw6iW4so+8+bzFtgyuY3Agwd3NNCfUHq6LjNpcGmdFddu1brlCit
ER65Qfq8UL3kKdFcTGj7DbXyKy/yKF9l9RfihURw55t5oU3biEDNtX8yD6oAwlbc
SDruYrjxOPiWKh2WOARRlpSvl8GB/spulX3dYFvcr8ljkgLLrBHmBoxZ4qoV/Iai
sUTkUZ3+3i2gl3i8tkvsaz+GhKQ4dTX3MsbKINtVnCiUPdroEsiM9771jWoVLjEg
KBe8XetmnWlHscavDnE0XtxCZfXAX2G+EPgAL4n8DKXJ1nuxd55gqFw3dTVtq5Ba
/NIKL1pJwfxFIYx65yhShrm9kEGASTwAmm5GzZCojqafa8LbAPDsggtW9gvIMVYK
25XvMwkQAqTRrvP6yYndCHYrz1b2yvnnCT6iK8sUKxzN2ZgFIBJmoPwtGCyvv1V3
YQ7R/DApGAjKu8fKSkMVnYBAwFKkIh4t3GHTQ9xnIhQU5u17SxfTTBgeJ5iYpAM6
bccVu6Az7oNmzjmg9OdNmlUqx5yRhY/7GGkqxaH0N4udnDgqM+zvWGsTm+8LEX0R
jA/Vu8N+DIo9yNtws+8fKxFy8r+cWH73G3oVldGk92phLf6oa3jCjoheZSuC208X
OMdQHQyHMRVrppw4QfgFrr468jgwhrtU/YEoGTmQm4KPMpFYd8Si08Lk8e0AEsjU
xgOIGBvxGeRvvrjRuQ0kw7xvCqlcaIe8tVWbysAnDTZV2IxZsxMkv6JSbCkP1jO+
nuOdDKbm/8gL4vMi2+gP+7dQdjDOoclYRuJX/2kxevrORlXEfVCiuVoJmYc5oVfk
bHso7OhBEzQuygHI62Dwk5QtqHaOdradjxA7bFv/IGcmsiBnKTQpssw781U/7C/e
tEG8xXa5I/KLT5UB12UkBaEypCgubyOcReThxRsMn0UxAoVmZtjlf/6610o4arwi
qcnnmJeY7j7qv2FP7JhawMo+IjIGPE+ndxDTW3E8MORHnYBSXbscJ1SvAxWVVovf
2CORqPRzUPESyiOjecq62RDsZVa4j96mj5uvKnCuE4mvyho0qH15vlAjk9gDmj1X
kjj6qCiZPWuyMBtUSHayoAuyzhftQY60EQfzpm5N+NAYWUdgUA1H2CImURijfqcE
gAfmqRn0efn+Jq94TPdD5I3vc5Zm8RvUTVm+5Q2w8bogoXMUsCXcEOKCE0cM+ITC
mfqG+VIdXwm33BaUmYo2ecGUsWQAyr/Z+60ecl1dlko1R6cxliLXyKzVAaQ+YLFj
gTBRCxas7IDMP2r3GXlyaWlZIORRKMxra1TVdGQVrWeMtyXBCnTP/AF/0srdGZYx
DWfF0apld+U29WpA2l80RcyaAr7ew/5DF8l1Gkl9M7/M9eN/dOX0yvAh8fnsGWiH
L+SgQEcA5W5Qmc5mHfFgBigMQjs5aGOvapX9HVPIi1cQKdp2A5HUsi9oftOEWJnt
VKNkVGFlyHWazhobm9IRBOv0UeFJa0VaY6xlq9ROTPNGiKscDhny5GX50vwi+6xH
aCbkoJ6iI2YZ5wcqP/paW6dw7HimJ8BtHurSttOcuRwDiRQO1lMWih2cLEtCrUFD
cQ9xGAiJo2+R0+KQl3ejD0HDTRcYk7TM12RYsqeGhiJwrK+A1wNaaBnxmXcPsxfR
DKed1Yb7Rl+8ULF7sQ3HDnGpvBzEr1MjFHCcIYFtCOeGWVcMx+SVtIQ0CAaTV40y
uvsKOgFdIrPEOvt94mudfo4iv9s3yn18W2e8fOjfiDrYggNH7arg+XEckm8xWnq+
C4w8Sm2FgeFfBCFYaBoi6CKu01qHXwj4tG/EPA62ugLgBLDLlLXB9/fUcKTOnioK
ac24CkJIiZny2QgtYjN/INDNYWNbrJTFXImqmd3bI3FaB7G1OXFi42F1ZSpp5rto
ve46BrF3vq12SAYZv6y02vt/8ChDyiRo01d6Uxs8uKYSiTXUsgK6EJRPMX+i+YsR
aYwkQU2xsUqkbGh5CmaNSN+msqUWzkCF2EBEZwOlhcgJXyz6ytMAuLhlIXEOrwSg
OeUye0qcdZIXPUZ4MCeb1qXPS95Jb58SPpbxUp8toGOumySsuOqPQdb2TpyMwgd3
xP/vCGMswWSdbA0iA07wHd59cK7If7exzkd5emkyKS/jFlTh/gHTIFVjBgnyxR5Y
0dKa9XftvK67EwAgz8f5+z3v42k0oTWaxZNUTv3atOYYQgIf7CILNx3EcDBhDtsQ
JlNpxo7oCQDNUc2Ug8bMZJiJ3LHWdNU+Ubrd6qZS6kA9guWRPivX6Y+8EcJqdFwX
HFwzNHoPI/l62/neQXEVBrO/sfG8lJyB3w0KK0vnz2Zl9G6cFyodjj1QK2fc4wl4
aJ/NXd6uJDRTjha8Bg9NFeidX56AOyj7nmbT7g44qiQoGKU6StxSVOg4hw9MkpAU
srk4ViGi5zVRWq/G5SYSmjrstmai++F+ODxJ1IXAfMtx/khDCHX1cyvgeNF6+F5p
vjpTIGKtESW9l18xy/L3mJg5slGzNdVt2EDNLA9ZfbjzE8KMhqEkedTU5dpd++dx
O16YmB1GuODRnIOo7IkdPvQRAEL/ZfmuwHcb/NveL+dqxx6jTth1w15b+sbUtcqY
eCehXNm+aTBFThU+UGOYmAVvDhIyvXOh1bEsjzX99G3thmO+dATSYWDkPYujsPLL
p0fGfwyTa0grvq0ivTUkJ4N0f0JFOPVPxqidXiO9SUIBminsP1WIzS3jfMRRPC7x
onq/a95WCGcx2nHLVp78nwJHm/++npkglDlsse7GHYPxNREVqv4iwOJ3Ggu8ltSk
tqkUSWar/zr6JteJIT49Difcxxb6wc6JjfjDCuy5pq7PYdI5K/0AAdVopY9qb7Vu
x1LTENOt9z4dxxqJjRtxedR4DIhiLmId3uf4LKUMk9FfIPgC1Sfq+JFYrA5iOuCC
6j7NKdBGdGjcNIE13/0UshatuF8b7YqpjUiJ0c8GI744d/iICAB3CNzSPKWeUdtJ
PTeu6MZUcyNwxb65nuw7QLXynXy58t+On+QMm/MuDy3Et9n85yp9XyrFBUfcllB1
p1zCmG1QpSJ86e7q9lkon2TycP2eDblFn5nxOcDAhGEDljnm+n8VRck0X8d3lk3m
NXkKd6TpBuWZWXNv/Z61CUbQ7UpdtRnmp5HxcxExhgqS+yLiu3iUXRrIWTxNjG3A
qLwUjyzY/o4R1ZjJU15eIDXyemVX56v9TbTjfXnil8RcoI4gfW0/jRrNKzLo5F5J
gcHIkpL3jsJ0t+qX+ayZ/PL/BselLFwojbm0osGh1PNFWjAvhl6NGIp+LyiMzjCK
jS+tobsd6hRnhUh++diC9xlQyi8J3JBEaF5FGaMtdqINdC0YtoTQqyCaVEQSIDHV
4YdpssX6eHyk0p4nzAI2U4usYaiEv2aCilqzTjeJpPw7/gC8Xjfcdt+p5EtBBibm
T/91syxOGN7CZAn4/daw+le3eGirJv8ekZgz/11IcEyq0HtyEe4mV+ROCTxoWIw6
tv32xy5rxclyMYR3g8lAgxSEHsP44l1QHC8Gh0wf5FBennVw+Dgg2d5H79Rwum3b
xaPIAowQu/qjY+8l8BaPzAX/8g4EBt0J1I3rhE2++LFO9TQ38SQ44FXbH9VXKn17
jKjh49HK/5pscqkqv66HlSx2/OxJheDRL3vkzKm01xFTS2a26Ek0+breHYPisE0h
T0I7BaODyDA7T3senCczcLfMxD6+JUhodQ/i1/weEFDC4L4kxNKC0yN3BQUZgfFf
1ZknZZnrgyuEyzbjLXtG6LYG3GMwULsrODa0Q0bP0FneuO2TA/bq5e9I1wnr8O6J
4RhgVPBBb90jfM4PzWZMAWCZ/hQ2VbzCKJaQK6HdC+hM5oJS4R4FtIXnZA1snfeb
y9OpM9ZDbsWXjJ3q732FBulRfbDConq2YjkUzg7hHBHQAOH/btG9ZzCVtevor3u0
/FIC5imv5USt0jlWD/il2MHF6IjxXWvhXf/UtWDjCqNMDYs9FLeKVFMWhEfsleCZ
XTduc8BiamVUiV5JOzvTYkTZ2LVD67zNHCRIRjbzEBtplq1oae9AxHcuaSvtcaXd
ufWPNf6Asprv1//BLkiDslwI9VZmJ5Yu7e1HnUrjx+InlnqUAMJdnphyHUj5ZqKR
45TJ8jG1nWYYCoY565SdKpWYJnVAcDTHmXDK/PT2T6syQV4JrxJqRtLYWFl62A5P
ckm+LYuj8MAdddt+oUWBxJVPGumq614uaLh0+3KhDxRFRVTG1sNUXYGaWQKX8HMh
x3I0iIB9fwMPyIAJGAtntKWhxh74/vD24Pwgc6lvPwTYn7TVd8Nx5aeXS9cXO752
5NA5Sa41eeBguWE+5ul9CzJtSQE5mRgSL8Qtmp+j4y5oiCWzhrxSEUOuhexzq0YU
+elQprt5kzCYoGniKhoz+u/k1xlKv3qjnHKy7RmIQYTZh78oLGtrhqf2KkQs3vz8
JUmwwcPB7ZUlrLMLpaFrgqbHdGzt+Wf2XuC+tnfnN+DMijGOkLrw2vJFjegRNhKk
dF52Bu9wTIvSfUdPAnBsnJRKSdC29/NtUwFzRoeXHot4kBlYcx/adUSJXCb0PsRT
5h3jXdZYVCN+/I+WGlD9m+jSgByBIyAc1T4nR7LaEKal8PFUgwte8wOFzn7vctfD
8GOn2e+hmZ5buGjzO1yo9QVnnUd04Dp/flF5Vc1oIbjclugkbT3Co3ReJj666xNg
/LBJSQ4hquLHRDhFhHBTX93yaqkkKR56FNePSlEHplbcDVIgkj2fZJAhrjsJUmn6
Y2/ebZZR3ieKsILy2/3ZtxiXtdDjqPFyGHcv0j1uc1/iD57E/aI7m8RySfRPq5N9
McD/WcO9kTYM7BUTKzqyeoOOhtkkB+2F57yq47aqv3j8tWqKdjS3htqHSLjpDeGy
N8mzd5f3i8bALxjMRTKQtiiQRhviR8iVNCA7H6GrfZ+twfyw3DTMpNJxZnGLmjoQ
AGOqV12alQQzOoPBdBE5jDFJmcSlO/afW9XgcxYpB/oFH8gAOm4SK/3dK8Uc5FI/
tHxCxmsxwagOZDGfDb9GqT9MhYiCCOLQ0h7y0vogcgC22P3jlNcjtqLOWk0vgps2
CMiyz7JJY8y+LDtK1fCgmJpW1BBBKOjZGVWkZGA5WTLweUpMH3MFEWs/MQsdN9h4
S8o08pNlVFFPE0T8+lAIB5baGRLMLrsNuAdM7kuPctYA50TnwtG9QjJthG+V0261
oBSGgGRs1Dc3pOOtqDFYiBWJHgtgDx/R1PpucXwXjBvTVvHNdufbQ8NZO42GvyB1
KpWXrgcXGYW2cupemn9EH67izMtB3ldWsC+yUrJVDmBUh5W1izV54vSMAiBUmUpy
AGfe+aAywsbIFNvrVJzNXJiBCzGDwsmDFGpsBDZo9PgSFXRYOOjr1ZyL8O7TXeIU
xC5CIN8qFUckHR6PcZbp7r1v5giTwQnjcC7lPGw3758wGg67X0rxtESOh+d3mrya
qD8lA+Z6ClVx5SwjnGNXhdYtM/dQbDnEPXZQbKvNO1MnsO7fs9G6VQ9XJsPBJW0X
LYIU0goWQuXzrFQh8ZZQpLsFEhZvt5FNcIFtE4G6IzO2j2eqPAFdDQdzceSrGm4a
JtgFZIhyx+uPOp07ktxW9yrCdoserLD2VE3z+RVvY6wQrJqKhGV+LosjjfSlNmz6
ggtFiPRubI7IhrG9ytG/AFCqydv1Tyy6qFPxEwAm3IDDtywHV8HfRIzgZ+gKeNRH
Yuj8RuZUttxAby8nO2tFCzifwqY0Ky/M3ARy7DfauzV7mOpYEi6yEwGHrQORgjA4
ORo2BmfhELp9xVi16+LtlrJ5rvWfDc+17rMq3g3PhsjeFj5y5KAMxBTlPMZukuce
v76cDUvzbTkVNBIiCNSFHuyHYzqs91zugIHwKH1oGmevoAe5GPETIsgo/VC8wj9Z
8BwxUhNk5h/4BvNtx3wum72l2Id+EXaHrEISCfFJ1m5nz986OlNZKpPLAWbewu6S
jIe55xmRHygXgwum2TVzNIiPRclzSdVoBmA4ozP6o49kx2lY6L5o+jDZPyi9TKi+
sNtN0iyzWRe8L1RF1zHGjFe3xr5XFb4kPFsnIyR5js/+Ie58pvLicvEoQrrc1aK6
1oD7Qk5Yn+4LicKxctpb1bpyU+W0N8UiSCRhkEcEt60Ms+DtdUUBPhMYPokgUWht
68eF5bSYdwMnFjWc5NQAuccUqUATx68ZstkC6U1xpL/bRo39ur+fBNEZEF8D8F3g
cNXzSedUTq/m/ow9rY+GzsyaLNkwcPwLsLlw451qpJvOeK+kfUax5jwAU1UEVYhy
5wjZvmw068hESfdX9mL9AcSYm0i0VzqjZKV6y8rXyXxvZf3W3cAXjm64wHnqm2Sk
VlPE1otXlCCtEsvFzopELlg1lJI78WIvhHZVaEtLsa9i7nRhX0VZ6ltLSqXTLPwB
wQYgnk8uJTB4LF++4U7mRzPwWCbmUmfvM8kq8JaSnEFodHQ4+4fNBlbjvqLAGdwG
Dv9ETpeSSWOOmwGpCsHmhCI3xZO2biE660mM+4EGeqGGDHgCtex+UH72olyirogC
ZxOcBlDHqo5mcRvrtguIuFhxAJ4/NiVvLznAH2nNW93jDniDl21GXAC3ukBwdPLn
fweIK42SRcIqr2sQgAmxYP2vUWIV5ngFkUI89O5kktqr7J6HrdvMWeh6ZxLnQfUd
I9BrRwesOPrZ5QDo7+uymI0ZN5QYWMTIR0oLaowYz5laRZ0Pf6yPAiRaO1/BliYx
QbHLw0As/32nJ8W3kVDYZ0wq/ZD2hdUDuUyZ+j/Bq85+3VeJXOqc+iGwmSjirlyQ
pA9HuySBg7aETPDRJ81oIwL7DItIiVWEGZf+nlu+FWxuPo0YujUFzvORMkLk3u9e
z2ex/jNF8hUO7iZttwzOVLl8DB49Yeg77dm8zX+BK9Y/Fb3JSqOb4+oMEe3Z5Wa0
19Eg4tjhyadomUTHw/pT0/B06tui0I3tkRgT53bBsJdjDgF/pyV45iTQpATLOAWw
s4T/LIoY8wIsjQHieMyKjFVySi8KQbFI/S7opVOp0FzBdn8Mbm+94+ZUIuBR9n8d
Ck4yqaWWKe0WmhKeidkGKwpWvqFo9xmQAltKnNnyWXCaCAflxz896Z/5Dl6J1Pzp
GyfyffzmKHtc7tr/3d+Yj1AKNhGnS3X3fTxJ+h/NFZhn6GbNOFNHoGKRBWuIPtDc
4PYzQA27gE9WTW954l6Vmh2MmUMLIuFkHSCfmho9bl/llTLmxlfG4CHBhtBY9a79
Qu/UVU00tFGYFyrxMvT6RcojKK88V5jE+/p/FEirXL0U9O7Fb/5gv78EXCHVPqVk
aGkNERmojxtafC35ARlvdNbchngdkiaPOY2dp2d4ch70LHXRga93/LbYMm/FNS5B
foC/wpidwqtUkEy8bF3JWubgyZI0DaTwaoYudR275BEgX/2EdsxILk4CcxkybDw7
BgHFyw6BjP2QgUYDhY7EG9fRVCZhwqr8SmiOX7vYddEKW9iKKdgKVWnV/IQ/EyS6
0R+Md44WwRsgKDVj4BVpJXMbnGMoB3c30l9tKennFl7Qu1vhi9a2+j79hVDaN0Pf
PLg66fGcCwhU9nrP8F4DbwWUo2WyIoa9IkQaa0MyPFQkNM8gbuS1U4znRegUBrJa
JL25SjxeRR1mfXWicRL282Q6MaBB9DhNGiza6zplXc6EPvF1k1SBZsOAINuVdmJt
DuCwZ91+hZGlx9skcOe0+agV9MNJ7QDOMMa39+XF3dSiebb172ByB5Rlo12smC+J
Y2Nl+5AYrnwNcaCOenIlTo9xrVMQ7McU804Zll6qr2XKm56T51h45tYhq5+nm5bd
+t2874kXAeHBRxyAz6VxAur+mzpFIYFY6+YGBQ5Br3aa0blIHP8ON4i0vA90RyU1
ljnAKEpMkQ52bA4FlNWrwgaGU8sIFlLktOHM8MfYovA3xyT5hrXfIWvVHjCusaEc
DuxNE5OnwiyrPMVHPgL6tZGIpISM2drysRNUCxRefWpxNooTqHWrpxPx31QARosY
P+aTW/lUinqOQWbzwj41siROuh09ul5olgfrTbY+llsUzmwxLccSAFDzmMbD1kin
mKOQE7gmHmI9/ul5S3pVor3iq1ez8PuAfSAdp1uxaVey8IQVf3kmk0tImYqpKtbN
Qw5hPke/f7vDz3/HTp+prih/drcg2j/lfubQ9v36fs6u4epNEzfUCchtWQFcL6Ot
cE+KfTxNhxKXZW2pCPD5s9Php+3eac2Tjl2+6pLDcOWy7GIk7srJDZF5FMc/MFZy
BDM3GoXdw4L9Vz+0K0qTqbEM5TgRhsOE5R6CHEtTe6CCXQ4QUgO7rwec4NyBejbf
yqlPUuOCry+EhCaMw5gVktEmFLGuRqEmP4hxQokIMprViTvy8DbzMfV6aSmQtUBp
o6pw10t+eh7YFc6QiYLll8rMA5ZzrX4DPkFpmWs2oBrKxJm4/W/85uXOfgv6WM45
urlJkdZXX1wH8cdVHHRzDBJ/pnqzI2GbHqMclTF+aTzn2YmYhOEKcWl8RG8qEN/x
fUUv6LPBG0tZRAvloxrCM23aj+TgyYs/STn8zvIkHV6FLfeqJ/0t5yPB0Tl6KcsT
6ALEFYTUuV/yz1Mgs+9HF5Ook5AP5SOwufFTXd/TG1zIg/06Db8N9hec0I0XZEAA
gJk86QL4uh/Vc+TWL6XHNexsugOWzl1xSd7/1kFkGP88dSI03WQTo0vc3lzRokqD
ZCgB/KYdBm/BDijJX1BtUX98TaLPKoHFw6pCV4zBxrB30RzG9AhaTmt+Gu3GJSGA
6cnB++OF38xGbvVyA5anwdn8S6z0Zv00JpnD1MdiSBjoYcTgOd6hUsJVBZrEb9V4
aTE23VBn7YjrKmPBMc5sIQoual37e/RxTQ+UywU+jyGTr6DcdQT0wyxlAbUO070o
FZVLp/5Jo/ULj9wat5Gvl1xIrlOM1+F0rvCb8vPzFR3u3WqBtIHNc9QhMtQK68V2
0vOrpYMUXryIh7G7wcVEHPkqq33I0YZOahaGnG33CC4hFRD+ZqjwrRRJxojCPVqq
OCkhZYux0lYc+lKA9Cm89En9nE2g/WXvrYkQUK3fhyc/Y20V4tLaH42zRP0Ox/lh
8fZhW1Y4ohIY7zV8N1u2ZQe0zasONNvkT7zOUJFQY/l1+WKiTE+xrgDGQVfpcyaT
BMeTOLvVRz/3DiK0T5HtxdDO1lxDnoHWRV7x5O5QowVtMWuOZokFpQvookLnUNK9
D4/dWaJy3YGu2/iECE9uyGDMcir2bT2G4X03WwpT7b1wwVWUq8qarB4KN/rMRoGp
kP4tWfzjcFdwKItfZmHHQM1y+7cibzOiJpKsrgiEiLaePNlYRyFCzJvz2psCemSx
yNp0DZZSAXYsmmmmZfl/r0ZxRXEGFVcZHmXjqIhHGnjhD2tv/zTsqOcWVhZHEvXu
ge33sA9fncnisAbM0hRrGNEQF/yq7GdP4jG9Hg6+dbQIbFet9F7RJ3Hlq46kBG8g
I7Zbo7XYBs+rG6KHVmv0PznodKIlFUDaRs3S55eKQfXM25l8yXbIpF9q96g8zNPk
2RdUOSb4KkqZFZU7yg1gvnC3wlWPvvEdjLqat556UnYpIoJC0NPl3ucYlDPkjdiw
J6ZaicOX2kUhaMAAnZiwNqNm/gv4EZ3rkBYfhrnNllyenptNwGaILmwwfmQvBWlU
Pjy/CDDsgBaOhZT4mEOHGnWtF+WroqB/gX0uaj9CXBba0BtUiu4S15PVtPVhdbhB
/5tHUUoY6ODPy7AHV27CByjgiYFNEgbvdmiW49Y0c6MTm+TNlGetM6wmvQGAABkY
1/XjPcQy3moMMt9YV6+bxt6h56flaKJwiCaSi78ayiNx6Da/k9YZdhwjK65nEtcs
rmhwh7jU1bB4MPxLTkK2sgBdgAct17yJXmb6VM8TWIQGr6lVEEM0dyRYDGHZzrXR
l4cLVAOcv3LYn8NMGbq5evKDZKCaNa6EtRDeKIqETB+UEBflx/ejKAr4c3Bcnzpd
l2xdkSDWlCQawbhheGli2lqKDT1+NpByRVZm4DoRGfSnmtS98g047D9nvSPrNZ+y
NRmkpg+lZGFXgXvBQOy3/CF+zM2ypzzkDLh9uQtQRJcLW7bOsAwWRX9QL46EF3gu
cdc7TW1RaOKNclKWwpE5NBVqAbw+fWOZhfNqzwUpSE2jnNNZ1E4oMWmKZUa5652O
RJknxRpYMJtVhQyg/+ZviO9rkoi6O8u/B+A522vNtQnq3Y+EUYGrHuLhAH5xOR4e
oQw6yCLhWO1tFAC6nQAQAv2LQnX4MYXn/6T2bq2tf4yjmpQt/yOZwlDnvcUug7Ia
nkXvpxceHbue6DEvidktSk4tzROtYKGpKp2aZ/ROloLrERUT89UBl8vjkSsK4JHG
iUyY0sWB5mbuwqOnzGcOa8KnTsIPN6q9idpv0DEoA+aIOPmhAbPhE6UQ+hAGoebV
+i4pKBjRky/9AE7aJh+qrve6uTYxNaEY+UxRhHTSj+65D66/8squyuxui9ypOAJj
d44a5n+2+lRKlYNsYCDtxFvgbdLwmGjWDIDM9zc/yVDvx4g8Es2+H14duHZvnNkQ
H/QyOaw8IPZpLJNv2L7oBNbdfruhft4B2GRhCLgE5U4HXkiomSevg9VzzZym5fAT
76TsxzrKpc6ecHVU8AegVo3oyOn50i5iUzNYVEVi7ZFqH9jxA/I+jPnpRNgaEQv1
89BolKvZnavmrYZT6cZ94vPjMgQYLmCPBsSI14VWljJWTWaA3ooT4rLy3yJqoff5
e22O+s3pDuMWZXKMFAKWUJyxepZzBlE0aTO1C4ezbKEZatKd9Kx2zvI0N5knIqQq
69D/r/AIQc8P4RG6m5SyX5DulDMz3ppA73eXBGRDBQRRJ5thhthwFG/F2ePiYmJk
B6Yj9h/oCuTGOQ2SLAZ+I72lp6K6SNxHlnW62k/mIh6aBFoKM4iUnfebFPkp+cvC
qOh1wBELz8CaKQYitTDXo28sArv+Kl1fAPf6R6gozLb8eP4znXZ/p9EU/78pxUXL
lOV98u36KTj6/O2DHdNALePfZRJv/u5V+SZK+5BQf378AUJBWG25ukT74e0W6UqD
gJzWahRrUTpPEJ4rVLu1PHqiEV35JQ6YN3Ab+/v3trHSZbbsiEZSBBSbUEIZNi1B
Ejm9cpLFCqsRDYiD8IPQ9alhjIqOCaR7DF7YS/KV7T06TzEnnExRaAEaaUSP/KUS
TSq/DCWVhzLq2NsKtol1YnA3DdXbE+WBC2sGV0tcWt8m54X3X7GlvTf4GCZHhurN
KGALKTXvjAbh0GGkN0rA85rPOZalfbu1ECN/zHwrI2Wg3xCXb2S7PMMYKfVwvs4M
yFnlCV3Sln6f+iqPSARxpA6sZwQzz2msrvx/ykNbuRUTz+CTWNTZDxKGActnjtuq
DWFMEUKcqQinRlnVgQOEy9hQCc5zm7XFedyGsMXhOZ2adSxpM6f0bUlgtLKVT3eX
4EMbjxdq1+n3255aOY19iNS97Hu/b8tmfVHXjaKxrSukZwHpEwyeCz7+LGS9hPWo
8HURerBdJc3WE4lSFiP0L6hcHnsWsdsvcr8LzmQSW2AU9Yr5GFpHZzRbrEoPSO4P
ZQf/Gfeos6WZk7jknAVgvXIFVxiQEdGv7/CJQG0JTugZbzpxAzSeceAhkFhQV+V7
MosmaJ948Rf1LUX1hIVuRebWXxdiPzjOGlcs5kRALsErVdWXKAZmgifBoM+VxYGI
9XFj1sSnGVq97qb8fKMDDTr8IBWsir1c2e0heBXCMDl9xRA5d1o1VzupPlobBO/x
GPb+82M7kha+Vj7DNaeciayvmmFfmrp/xljw7ab1Q8foHe5K9f6Hq4A8iKCxw/Wf
wPHZdnEXwt5E4xDS7MTr+jbsCAJUQ8pcliaOvGhr8KYpTVTPmj3B4g99sl42iv91
dyUnelab68Fzs1EPUcSlBYFmRoe3ar/oFt/bilr7MM3+4+ZD3FHDk3JhQJVl9UgO
s2kJtSyH+NN/O2rHwE+97gM8/CKqnFWB0TB3/ZYaOz2xAXsH2aZWK1+qAAwjFNkr
2gDANo84dcJH7buqb+pFdtlmzLlQJSP8Z5cAgnowlsDOMgmSeG6w7Yidp/9CEOd2
IChO6SZIX4FNy98DFLJcIhiUmj69vF9NIgjsvOfO6dqfopB0g/mrPTwkr+7loevN
mm/V8ZyDxDpDwJgtDAGGXQVfYlG7YSSGcQP3d2+nHIiSEWlQs1H3BBEq2pm3o/3W
xeETR2X+64TqcjMij/kmDHp4ilqNr/mQe5iAiRFyrBx2iu0Hh7iwWfc2Csts9E5H
vP3IPdxDvjhV8R+7CUY5epWQEudlQTZZGeUnb6SMhCTAfYNdI2y5AYvScAs9bqEh
+xAo8GlSdieEvObMMtAu4OXygx57WV9ed70bHm6C6IZKl+nZMYJuxdDjeTwETxSM
SHQ9A638MUIWbRg4AoAfjSh7h1N3bSpHq40KnxQYzm2EAC0sXcdKE7hG61eEj0IC
q1QtWeNNgmWc/A/cAe/e/O7SXGgU78pYwat0VCxZGYwUTTJUYvQsyJEX2p7BBVwZ
NRz4bQDTAXFzq6/Z1qr7YdOGtkl2XqiSyo5CM+dmSffiaQsL4osmt0buNcdv4D+A
TBB72TOml6o8l/T1bk3jsYSyHinJXBZOZ/Za3NjL78soQI3r7RXQQqyjfOYTIfdd
mdv9VGhONcEnLsVHdWAZ91M/x1yFQdR9CDq2MT23jth8Dg5suq6JVU/CaFF9qmnq
myU6TEwQ7AiHHX8AImosyfdPtCN0jamXNioRcxXcmeVHXvkpWY8tI3EvcL7VgjzL
CwqbII7q+0dg4CbruaCt5NohgKWO5apkYW5dWlBZBZTV4FR4pHyQOwonokAahv1g
4PfptGhZOnhnDC1vmRlmmdb5CzYtOdiOoYZ5zWU9nwqM58f/pEBCRE/DkiXsTbGl
9Iqfq5mfh5bTskX/vQITQBo6UsR5q4X7zY6xrgCps7PIVUdPWCUcxV84oh/WVEvB
nQWgdfSwoIHxPz7YJjdkt68ypjV/ZGkN9ggzdN0gmwByLugUrSdeEQ7FJbDjFytp
0RRwBYt9CvhNydRCJSR9jRWBaU5lvMlwZqEgazkfC+h7x6SoCG5l0JMn6kpzG/60
ftGTzi27c9KkpWjV1l0N5gkVtJvaOsMObAYe1RllOnrMB8u2CmJipsIV8kVjm/Np
CFyEehHQ2Hao/vgi0NjRtANiI9LO3Ymmu0hjgkP5hnoSej9u5SKzyQkwSeYrO3UK
6O40IXjxa7fJoAG1pWz9hJiBwwJUDwe94qAubHWXVOP5lColbahufe9Pa3xCOf2n
sxzYU/oVc9WFp8L0mIBSsVCAiyg+zfUoE4YvT2FXiH7zw4P+NvJmE4Qjx33sqVEQ
Stu2zKlPTxL3cQvPytjO1vw6A7IgvAiBUMNZLlNXxefDV3gQQ2kqGSP5OGMnIEOn
Qs2gFLuJEdxIXsDHt5ph1vVlq6B1cW83SdKWcxYNqDcnwFC1kiI06uvbV+ouCpx+
9zNkMJ8BKZIHFw3x/rPnwRMT/N3/28cjjZmYB9WBguR5TaJiLRDNQclw9S1p2WoU
0f2nsQkpV2TkVins6jf+S2FWV9S9tHZHOFVjxN0U0Ep7SPAv3RXfS/65i5MpCY9s
XMka1ebgo0qCr1rHRu4ZZGICiSqIXfykrJqcI+y8wXtv0AOrsITEZ5fXBP8GgsFN
QkCRG7SBWlAuixXcxFLxEs4Frny2cODCYjNpt9aJb6s/ga4LEL3G8SQKFu9qNPjE
m7UZ7dTxvo74byqrSmhlLnE7lDKNiZeWAO2W+6GznVz24xHE0g4POkhHuV0+Atxn
bURFkKDuzMg7KFxPenf1j994OM0axLoWiJCAhZqf/V2PWceiiV6z7HO+OwMTQY5I
Ahr5OZnWMfQkYeQJWAVzpNb9BfYEkZMHtwf9j6Zph+hqvlS/OZLxvXlloD7DXvO2
oPy/AC9ItPWyyk66kVnXBMb1jx/OOQxyIlH82WpI+nU+UOhznTvKO9vhgosTVASP
kop500xvUOHxadyyV/Oe3N98AjI9Fpke5LNcBU/8bR4u9Nzu+RoDHy8XVXZ9sKi3
DTMtSB5/Efqcpcd0WZvGJKggZEUjB4Jeht9GNVO3cab0l5l+gLHDoU4j8bZByHFj
uHkk1bk33TwT4BayoaDBib8WeSESu5ccEyxLytiMyCgkGymvIRtJ1v/dHFoLNc4N
4xBCH00J18CzepWfyRi81P+M+uFv6dsQsmouEq0FMCqTzoZiMqtVp/HoUGaz8pC0
piLnKHI9GTeIHkcU0OB+qvzOlAC9VUMtjRsAChqkHwED4AqMp32D9bWEKu/AoNjH
IcQGyqlWKBMWzw6E0t/izE9bo7CzE6L6W9y560eYgBPtC7tkyZ13dFDiEbW+5uGm
EOvumErsjj0FJ5mYKRGjO+PXMuTPfDM7i7EFVU8fniuCWJhmx5zsMs45amqTTM4b
KmZ/5rcU2NxoT4yusLFWFhr2TRUDH1Yv5ROAP5Ju1FHq2CAvwS52mOvdjhNbDYIw
fLmyFLnLOU/A+RjCeEPlxVbxpPNmZhCQAAbuPWvMQOVeP1sCxGW6enMiNvc8VlRK
qnnXwodNBJX8w3mAJCCHRkL3rc9agwUO+qcyEADfi3pCG+kWBnCjYPhXxskUv78o
KMucbuYtC9wh0c/TFA9p2Q4/g11gRFbH+me172s+7/lvWnNE7oKfPJ7NhM8MUqLH
SXQpqVpPX/GwMDyIHNHCKm8/lJy/ceIrPMGi2+FMRytKst5E184dnV2BNezOzlS6
pWmyj0kdqbCKE3oKS7vH5rcbKfh77RPltSY3Lgt8dq/GBeqFx+uVv3YaHxvKUHf/
xo/YNqrJggCuyJcNr+xd1LrQZgg+Wq7Bx2Idyz/WXgU6jtG1ovbbBC+fuDX57SOw
/eTpcHntobvYCDHzrGOfFQlJwZtHwJh6NSkpmeB1i9YPZQNNyuC6/xmS82jCFxu8
OSlQ93WJPj+zEtJnPiqJQOXQ74PRpPkqiQzA2Q9mkwQ2xA1UNNngOrNU4CJUnoU/
D0v/9SS6dglBn3g6vaZBLvMc1AtLCP3kPAQ6+pSvDhgVYmQGY9nKlqcklVrknLEu
22Dmim8xD8fQ0R+s1aSz85z3ragg8mhI0uwHiwu1tmoWLv9ZkK1ggGSGzXYhZsga
fGnFDiDkCDpkAAheXerLO1UKogX6EjGP4B7MbOmeGEBCBbz/m2UmISZOC0iUCwFt
DiwBBLGQIyt8iHHu7Jnq1x7TmAGZ/+fcTOJoAWfaONFIrMKwpKylPYvzCfO/q8zc
tewX1ywR8UTh40eiVhx5cI256Pl2+eT1VWTw1Wdhd/l3rh7lhfWdhC53vvN7nrLD
49P1UWkKG5ymEIs9dTajwC6yUrHFZjRjIzyELgU9dhrGKAcXkoTWOyUf6aO4WRVH
JhH8+IjiVBFIZ3jO2/fBSXniiTLTvaUm4UuFOMXQTQhXXeUraNU1wXdxJXyEhgw1
7RfGX4SGnqepCc4WXTvXeI4LBew3mOGAQlNDgqPAbkd4OrH3t/0XylsYkac4E/TM
nfe4907Z7yhxoiWQKUh2qpnq5vik9XwaMdhH0lKxqNgs6gUkciQd279S1pVU/vT5
I5YdzC7bmHKK3o24Sbw+1ZPwlGexY4Oo8lFEon9A65LHDkiCHNl7ZKNQDLemnZ2x
E1TB7r+o7PvkD6TBiAn4JsfLEnlvSbgQcQKO4eZ+3eHiR6Pbs6LfpO5u64Ltr4LO
oiOPSvfYaG6W+iqRfBW8G/5xcoHoVS/JDIGkn0wviWSwilOb1qGTutNEaOfOR1Wi
zEQBaupCr2Zh/s4Z0kMJWX+rkcKXZX+bIG/gavtlDfY/Q8dJ4Z2oRlGMtZd9cyqy
ZSJKP1nVM60mV/ED3yLEn71vjrCucsg8HN1C4FpJ46I6PCRDDv5tfcyoWvZrOIVI
XBxOF6U/1zxTPs3VxYDWR2ceXwzc35IZp1jh6uq5wL/iKi+vp3r6aFRv7dPFA4Sr
zc5Urq5G4TMOtFke5rA/DPYBlQ4vz3D2w0k1MKo/+ZYPtD2kXUusNot2iLxssqR8
WuICXFXEPB9rr45SC6MA9ub1FtTl9hMwGaEC88hfbnbqa1tOmxLmd+/3LVenU95i
rqXAioiZkbCbCdZkikDF76SpvPsD4vFm/LyFm8Tvz5nS7ovqGVtzw0q16k4hUJg9
Zw5xzriQ+Hp+NlGlK+6iMJtSh/ZOfTalE05polUjlSX03hrh+4ow6wceOhf9XSX0
IywCBnqPDMhnZbakREAnuWeCJSAgj4nIWDu9gXpMUqIJVjIP+246p9pZrVw1eVK6
O2ilG6izJ3x86/8dJSfLFrwciB9QtqtfTfoWyD1zQtSMiDBvb8jTO19vEwMHzAyE
kf8i8LPeHyYEGmyH0/yA/m5J+jt5NSrNKHa1j5ivE1YMMnIQHRPJ7rP8J0h443J3
6cUczn2HHzbkvpnKyRBICaMAbQbjYseVrVhCOHDwRykxjWnf5PQzHsydq6Ry+bjR
qf8/YYqDARkaMCwEt5ORsYRYPmrZ+SNy951M6CivsT5NEUQoBq7vSjc1xSiodCj6
n1jT15jmHJ5ZoPqd/LBhuPlC0ANGn2DR/6okLIXVbl2yxhgOAp4Zowl7Xr4oQfbS
DXryx01pFtj6NEBArfkRQo4FOGa09+CysrCpDbDrOmJ77lm0ZNFcJa8FQTiddaUd
L+T6H6vwFGvDi4ZBTr63fDmPeN7K0xyy7ftYeBPzPR6ijhrzjkZdVWaGD0Awgb99
fOsmunxeGj7ORjQRlktY967la7hWat930dzSI+2zlC7iBSebcql1TFwzNEh2eP6r
IpyVvszzwV4vlXozc+87zsf4V+onrCFr8AcJrVZ/viOaObXb8E1of86L4PaX8o1w
0HMFlirY0nBdx0dbHuAaJvVBSLNaR+dmW9gLnwzasULXVBl4ytSD7K1pDF+ZUDlT
FUyzfUrHdpqpHdziS/ZbEBNYvhsRpiHhlix7fxkHZaARqwDHhf+j4piRqTloUXhO
nrEPNkZ/Mnxrdeq0Jxg52IvUxPR/4BFpe2eJbUbYyocqaK6tg8MgGV2s2efUCHz+
r/3CFzHZz3AE4nM9XbRlVZzWtNoOAcNO95RYRCwafgG+9lzaDdg4wmZ7bCSkYNY7
VZaTRsS58/OSUtp8PCpndN53PAje2NrtbPgmAfm4XHi6hVM73YYWX4+92RqU6Bxb
R0mphzR+LrdtxiVLPViNxjupNBMfLbfsyL1r2uxrbjFc/PgRKEpB8qrCpgVJNLJA
kukKkw+bKbjL2Z7bwgW1Y/gqex0frDPG+dNia7c08oNAVzrojPLkv7rdpWwtx7P0
8+WVEP754Ic4zVvOPXdpcBDVOHtfmVV51x4qvebAtFrS6wVmRqY0GylM/rM/+Iwh
dvy6PWdAm6nXPpG7tntWsF0+h9TAyRLWCgzlmF9D6sa50AG9nG+O+M14CLfiGEye
Mk9Gndx/cUDlAdo1g+BTSQO38cUmWYPt2rMLAE97LKCOBJYw7FA9c8UyruQqR/b1
GIzMKRjbvYjQjD2AC1EQrgQCYwGWY7HQwuZJtm9jrXJRB4aTiwgqKRq2exCNzDMX
8i0mY7lr+mOscUIM0fQtRoGk1n3Kz6xhYmgpRUutASJQ+mI4GdWxNpmMqnZoado4
bXN7Xch6RamRHksAQtrRFgT/FqQomeYPWWYpLYv49ykImVrGuW81ANY6IlYwy3sd
WVJ1ujqvlUXYY//DpRkTjGq3GXnj8RHJ/Tj7DRrwHDevzWBCLFOi2THgKpvntQSR
splrNGSY0TiKI7JhjHol5IoyMNEnm+Iv4U7IkmPL+n1XpGm44qqquoTmWBh9GQ64
e896LR7RcTItmChwriCByTR8PPNy0X4H/9R9vAjyA5chGIGUVUUzg9Nm8R0L3eZS
CvyENl9KVIIV0pHi9PH2dduCm6yXyK3mVqWzdT61aVFxRGlh2jbWmQpX4sAPZpdr
Hlfy+yo7G7wJqOErdrXYciLmN1YxGd+2J3by3yOppOcYrRIug33l4B2CYt8T/9Ok
wK4a82Fc+D/X7OCVPkcRygrIhPHpA9Beph1sNYlkuh4Jr8AY+r2a7Dly1TGiIBYo
Dfm6QS0n8kEe8FtAV+Dxw9paCgWeBs5jYuX8FLabKHYXOULlajvVJXY87dl3MyRp
HvGmLW5Tlzxj3H17VMmvJ6+PdF7b2JqDxBIE7ZCNgK2BOG8fMaNl0jmX8f7AnxJE
gc7WJSZndZYlVkeSJM+WKTKyVPmp1EuJ6xb8ssZjo5QcDAbYT/KUJDLkrT4rIeVY
kxaebQ40VFTklbpC9yt6BXGLtj2eyaq2Qkkg3zKV9wcXkLyVSxgv135ezOfBfYAb
Bb4hvHh9M9CFkJm15k3CokJvtoxwOOfipWM/IbiGDhWXzVdD5aGCsCJ9dkpyVyQj
y3g6foVgmDPlxAXq0bjv0cMdMtsuZCKqy/isYy9HRjMYCrdc4epF5VBdi9Xc/4ox
nWiBu14bBGZAjRkpJKpvN4lTo4pFzF0SR4G2WNaVjhVPG/Y2puvIa0Nq8JKkvxpc
X84K/SHwCUHouPo6kwwRdzK7Ne6IgHvS6LrzLRuuV2QxYh3IBTq6B1CYGwHmDIbL
9zRWjN2bXadtp5wAtNiCXfKWci/ewAaHtv27fr2QpDpdGXsVVW781g1IaJb1JE31
yIfeNbRYk8S7E6MuEFbXuE3Zv0QVr+g4hnY5bEPEynBz7xFN4fW8M5HCVj6vOk0m
Lxg98mgyDAXsyF8Dl8XMBGNCU+ZJctW563kh7eEgvOYgB6D8UNFFkSwuYRJXE5RR
WwbKP8CzBUGxI2+MSF46Dlt0d3pJ+ioDO0ax0VJMX21661HGREKaUEFjeCeF5blY
xu6kcz6Q++QUKuraHs5NLxtfBvEhWZMF1KONm+h2vP1tWB8CbAMcVyfgKMpPdKGL
qdGr0j8RoKSg4+VzYj+blKwVWkg8MzJUgjvOjQDqx8St1xrQL3VD/k+I61Iyzm8W
rZ9uN1YaVRh+puB3K6XWXvCPZvnN9OChn2oJsGbuGBoybEpFmjxJQ0SAAukeud7Y
qM4V4m9epPpOXBRmBEqz5u/XxCcQIp6KADGcBayqDaOI4Ooep2r4Ltw5r3ZG6B32
B1I+ow+ZppFl2caZhUZsvM1qIDYELCaFZgO73tY9HFETFliVhXZtxBw5iWgXaSMg
ITOym3KXureWnYs0tlGVeMgc2MSTK0kfOIycgzf1c508y/HODENMJ2GiqgHeh2jM
XCFhyYaqTYH76N+5Ncoh5KOnaVV50f2+fiiLRTWrrHY8hDhTGv0PYQ0FXWgl7dd6
ueHWiJl5VPl4FBLgVryeO4+E1J4QSTRKPtbpTGV7ig7GY+oQ2JjcjWi2hpMxFG+S
dK4lOHTq3c1+Wlti8CNphFfgBTfrA3+x8Wk7NzS21PtHbiJshdLQQTb83bnnwAWV
aogBkH00xDKmp1HVZw/DlmBGP4inOeAuw4A9nQIDD+py7QLs9yvfi2a5q9nBRgPV
W/BbKyyf80oN6Eq52D7T8eZcNBPFbvNQhTLW/VRI9qEi9FMWm1v9lbeAzOr7og7h
iFZkLmvsTl6srZF4mWW/EktBGKnCyQ4SDDLYB/dX4MPtZpRcPq8Q4sk/4a4Mzg8r
Qq8aiDqHrHKKhByU66nC8JKYI6gD4spBlO4YMl2u0ZfVccOq9jFHiCo5ELHcOYbN
fpNkR7Y5ovO4Haiu59bMaGzb89md030iaxbFZYPg7beFgoGYBPhQuOGAh6VSCTMo
+qNpzgXlJpVIHup5oTWZ10/aEzpsZwgO0kHP+/+QS0ILgq3f/S/UBr205BKiFYPY
sfvFLHJFTlHfXcueAqfM+pTvm34TNNZD9AJfA0h7hvEUNsLgvtXFEnri6OZiRFqj
uUtYRXCE8Yr2ehGik9Wu6yBrsjPx25GZ5wx65S6sPb17vwW6Qut5HRgS7KRqBTKD
RgLW7lb0+wNTCZwCh2XEoA14Ma0yWE4CURmqzMFXdedwCmebVjdHaAbK6LB+QPsk
pUC8edLZV9IfpvfCsMvrcB47fWDVnIc2/Aiqlt3Bcs7wkis7aLnv9BMj3KQDlUlM
U9EBSiozErRLxmxWFRlgye3N1ipF7o+T/6ev+JfwM2xXw56fI3nH/3OeizgjJHHy
IWkNMA5/pH6YyI0nD4WqGWPd7M6R0REKSbPOOk00vLw6SEYTZXjEMKHc4/6CwvBK
xYyBg2PyCzJbV3E8n5QP+kSI7FAljHQ+Os5rvZ7WpLFxRldU35zju8PvqT5hTUk6
qXqd1byAhih02cxpl2/pGh4htSLVxNWveS6i/4mf1cB01hUfYfh269b8qmZQOkpY
YMeNWqqSjiFDvpzZGlkbBq4dKSYSGZ4EI4lax/Rd4jM+nfDYsMnl8NboC0mAGDkA
Uk54DdIa+dV8n5lFwuMaFMmhpWYoCbIBg8so4A8HkgrRGEeT+ETcHDlhkXNyvQV2
esetr7Xyxer5ZYfcgU6n4OZ0Jqr6iJeipa+WHq13lGCy2bWeWJIvT26Tn3HoCWP2
t+Z/2rUggyPwNlMpl709712jJqSxHL993N1rMZo2HQKBoTGpgv53ycsZ+njmaV8W
prAs94cqoDF3su5WLCRsSDkt6zL+RihvgGRgluHvaw8plXOsHYjLXwyUjq4fT62v
BhANtuHxI7idtSbBuiaDCk5gXldpqVXXo+vsSZDgHP2DYGpTARsF2doafKtkIWks
gdeQgFDZ5QaBgEeb2RjyrNrzMM6zJiNs69JelN7hfG1Cj0qbqfjnxREnM76KvXle
NRoKTsNqRAQ+hOd1Vxx0TixVDlQn5RcosY/pJOhfhwJrM2X512eEPp5RJePMs1DM
OOvCCBlSaeTCBc/IktILz1s9QumP7xW2xizRTggAKTvXa6thmNspUzUXBhYP0rc5
HhO3jopLlj6+RnlQHU6ySG33/jOULPPPaSNw2Vp2TinYzVrcIo2LBDNy7mR+2TAE
WL247XdR8Y25rwYydDhNYZnYv1KEdQ0B3jarHllo4w4qSVR/gezdeX4qY/orRWJu
Dwzu97Jw9GsYuYwDMhKgfE1ktYyQ9cfhu6paNaZrDtpsJVbdSlDbP858MVskQZEd
wS5u2mvOfYB6NWMXt6Z4FzAzFZoTsgzCilwqhW8BUV4w5Kic8wVXiyEWk4SwFLhF
x64pBXuzWa5s/0u1shNbZ+DIvoES8yACq+BB+tWxBna7+/ngW3n4APK88HHEixSL
e584wOl57BK+JspjbMKbsEoudu5hliMODs8bV/Rs1T5yhgYFpoXJV+AJL+NcFG4/
htMqrfnR9w/4lGkSlTXFsCD03KSOqvP0GeYQUlcfMCdr+XUb6gNyMqg02oOH6WJe
IP7qe531RWtprQZYd10Fk2Hw8HaXwOOc5G9zxn2BafGYIut9XayzV7I2LwkVqONj
9qTMOatjuWAT/x0WCFJkdQhvymT85Mf2t8WeOSMODy7e26I9Y0OYvSXby1vn2t9D
9mEyIwtwH2lGuzMhLD4VcH1ydY+wPsvzJo4h3tHcqt9iJt0SfoASsB+iJb9bYCVv
tQD9ZrjhbVUXT+1f5ySGYQCihEDs6GLDgqBTE2Wt31v2Bos3ty0JclNHJJjkshGs
WdsXzNNG74gEINCcWQXHzwG9i/KYHRUfdnXLQPJ1FcqDswNxsVojcLjrzh8Ks2cM
XULwwRhic1HVa3jOcnPKkW3bF+P2cV4DzsU9oABYy1v60wEGBxHtCpPKyXy+EE0l
329Dh/JcFwRjAgINM1n4SALT+BpfZA/rXAAxuZh91zwQ+JxGaK2sdYaonnXA2uxS
LCnpLDst4T1ZaINCUgmYyd4NuoI6T0JBtma80xZMrnoqt0iTu41pu+NHQI1EDipg
sC2gAO2sekp0TTIf//99ApXqlWsDMri4DuVXPiLeEkqL2n3Ki4XBtQjMg51DX+W8
BEM7crPVhCsmvDoU3CQ+HABHTFK0B4ehQRlCw5tmeTPOUkt+QeZPfyHaoPwueE1N
WWta0DzD9VE2OGoFLfWPfWnO3wVsmN7mLoPA2KkzBpio+bLvC/JcA6jS4TGhCZF4
FPoqH1/YWEyUVvPfPDI001+kRzteJoYZfpKFoYG5yvNgG7g/olrmqJYJfz7/VVm3
i6DSEjBon2ElRjajAjvrSnzlZ8VtWEvl++HMOUJvuJYih7tT6KPxlMBKzg59xl0d
wJWNQdaflR2rgP7EUqKSNLRjK6VMukwNYsKb7n9mmrctrNf3oDshQbIv0ZT9iLKv
hOvTWktD8zi+fwyAavkQ7UF/16/U8qgLKBi4JAi16GcBkfOW3L+pQcEfw9hf3gVC
dV3lTN5ymEwUdbFflgvFJ6x/tQdsqfBAfaLZxZATBY5asnzbzAUeUbQjjBq5pLCm
Bt4/jmeyIFZlLwiC4e/Wez09gbp5BglmhqA8A/H6Azxx6cJSaQg3l7sHDq4WZTe4
ZRjJi+NQgCXL+UOdRfhLYFkEnCvLOLqDs3MzoeBtA4lgWAHjvhmKifkPPM9/1ILK
EKqkrvKLlpQX5jabwuD2rwJqpZ5oe2ld4AHU5gM/8NImtjth47yfXIMW3ByPCtXq
qSRkJQssk2XGEIi6ODe62eZAxFGMl+GJ19kCUuh4kcrpLIK7u6TzkesOkGoTobHC
zGNoPPZN7Lfgz/lfaGAL86KAyU7ZuWKA62og/C6iw3OcBChP9F36CPVzTVDr0sE/
emTI9YMJF2LxAdpXyc2g4/dnkxDJsJHJzWAX5qYcVhILQIa7G2IITO5o25EqM8tB
46zKzbYL+i9b8CdDoNmTszniGRlwV6GslDmPkOrov2uU/6UdQGy2Xgy9v0RhxDmI
Hvt136Dr/Facdao6vi+e0PbZY6DyZJMh1GGoD3ICUNUN4UkAZcQoDDBse+xpaPgt
s6JDHFme30dSW7/syV9XmLU8oX2EouhkoXX9oe8zoiQFRn+otOd+Wn70PqBAkWW4
9MeNrKEg9K3BPD5Qcs9HLDl+hbircPpEpx5mGatCWcz4F4eCz/ckRkLRE7g1Pijt
0TdIBWbx26qzU1XqwW0GGdevb0tL7KbUaok4p68Oey4eD7BxzkRMU3ZwVsNZHKJy
oNfN7R/FDeQIWuGWCazY9ZNJCknIiS+HSL65+4/GUZ88cKUXkoR/hZOG1umn/wXS
GzUGSZCPauuVbXPySWkhtRXtHsk1Kvi16rHP3UGmVjO1Wn82c+SWC8ASrCoWKsJM
uI3cQc278wsSOJMqAlLQ3mp4z5E3f5HZ7jNfLdCtkFdQDr18q5bCEsIDMTFOtuW0
/RELRPWREnznV/yTP8aBJZpr7+y95IdZMwNoKhu1N/p/cOPTbSxrl1RB4V7RnlWl
4ncArxO3ERud1hoLTzRiAB/iecuN8bLch2hgqEnCzRueZbe9OmIRkem36v1gFnhO
pTBHK4ZYge2RaoWRQNfnA+FuCeZr0JmgB0uZBRicSQYC3Xc85VVCSkJ6f6ulanKm
Yc8I61mO05LU8ZQvhj1rhgEvYUk8eyaqPNKbTfdTl1eoCjRMDyg89M3ikS2KgCI9
KpXFvzXjUtFfKZ6BV3tYWXkmC6NBOBO7Ml6WnGN2XSBcWHSx/7rkYHDdKLm099Lt
pnwH/XlKw/Sse1YiX0echxgbKOkOMj/Q+0sknI1FArDCGkyvlzsQN4Z6WPuEusyf
8+OshWwK2C3Fx1rV3It+l8TgOsy5o7cuZtxG5gAVodOiEgaLt/h+tL4fa+Nr/j5G
YZiglyZjGddu2sAt0+0XBQjFMJssuXMXiMkzgNzqFkia1hhr8oHY3YJufmMF5pHw
+jtZxGTPnT0I4OP4sxToHHpvytnVF8i03M/tXYkfMDDB9HwLoiDUsS9jYmBRVt/t
/Y/2f3PtRwSyqL+f6DrdVS3S01rxviJmh3ukxg2Pbu/MGu0APrWF3JW0Lk4m2rGR
hWq5dGWTKX93FKlNiU//Rx2ZyFO37StMX14lJ5LZaPdWleyq/Vly/RjG3MLAP/zm
du0iKruQAxmVdWbsR9A6IlYGNJLb9FViyorGNYdaF2bkqWJLAkwMitvWONRCJcag
YBocc/2/aDMy/nNjqk3wQqGj1zwhU1CZMMoQGWfOeexB6ouJNUmjcp+UycC8XIvW
J8RpDojPz/SsMamTob9TDdcQ8cVXqyTQNAK8FNCLwfDp9NgPqvF0yiVCuJmXTI1m
4m33D5bvXhpUuYuhUM05OD5gJn/PJjxNKFlmWiwjbLrWMRmtyKJk9nbSb8NwxUGD
oLPKy5d9fQ7EwRFiNw3s0p5Y6HyqPPD8cVxX3WoGW+p9aABa+gT6W4Soszb0aKqp
aXK6Oun5KRLYPTMfn6LS9q1mfDxkvxl3NsjbZTfd+KMFhvUAQkBSky3svA2IpuhQ
hVHU0CvPSALGjdgjhg8bKJ4n4T5fuev0lzAqr8RZtunpoqq2sjf6d+J2CKQ7qwvz
0pJyptJF/DD8sAgXHJYtJVzkfhtwNkCHE4gyrHU1KOC3mM/twplOIZjNQj/IuQnf
9lOt+ahEMq7bH+z6FpPVStFs0RY09rcUCdSRNOdmyTGn3JeHk3ytWH5O1eEcczXh
jmMaebZI+rbVfuH8WxNN7tmWHAi1o+5XsCTlcTnAm3eHFaAD/3jlSXL8Ac1WatJS
Ya9QXP0cyteOvgswCYa0AqVW+zPa0sY0WjbhahfI59rZVOP4Otcy+sGWS/JrfmpD
gUCSpWG6cyBlkr7iGiP0IKEeF+fkSmuSVmKL61XNbBlrFleaVgknWJnuI1Q9hUPr
3E6Lzjf1iYrypQM2gfa9lSBZas5eCqwj4PIN3qcHfMevcS9gvNrsrbegk+hE+ZYG
LQoxJPVjASRxW5SzwBMM+GmjgHZLvGlCTueGz2ccFd6cw0Uqe1UUaKfWUi6Q3jiS
eDEvU6zkeHVetOKBHQMZYtQQ3LonePLqBlCBFTfx0UM6PXgEn3XWJM1RC4UYDV8o
TzVGVkMwM8cdPJ44unl4OO//2y5aXerPnedOnrdlC8qsdFZWAuoGso1avLLdWdg8
dLjCD+0VEKUD8TbKah7O8qZYf+MtMEmOrIXPMrWzxSYgDfGnxcBiTsjeE4OGAmr5
p9TgLcON6ujuM+kleRj9dBhhkG8ThQnVLfNIpGR/9GRCvx5JglSndXRU1Z4d14U3
df0M52aVsmq1fkTX0SIkvcOShdbvcD065PlVCV7q4nPhVkApPIuCOtp+uCSw2R+N
h/SyBOk4gFVL7PWYHB/8SeQ4RG1BoA4V0mUkxlvOswwg/eYguypeZDY3DhpxGmms
tmqBA1p9EruGSuHq6m/Gs24G9tIFu+p3Tb5CUcPp3WJaPc49vywqsKkZvjTc5LWN
es/lofkEWJkcNpfI0A9RvC6Yiq7ZNHUrkV850iJjWFWad1OD187peOib69ZeKwaX
tfY7fX0lY65NrFoLCQwkz1eK0/a2sTkW9G24XwczdswLs49ZjLAOPvjIZxUDPw77
DyBdFuMJRiHsB3mv5jpamO/bCVBruG4PMHM+vzFNEjTfQamKOyXKoy3bQo7DQwXc
9wMUPYOrxqsQgFmPox34hlMBlCZEBZweGT1nenm89BWVOf0fIeBDwys1T0xJJjkG
e85ZEm+kLnf/pkKwvOm0fMoG8lY5Kjo7HZY/6wHWGgbveaVco+4SaDvfA5KKkSOT
SHT8x3mLSVhtUWGK5qIrhny8jOItWp+ThU6j71+mwlpSW4mUTk9OkZySuYs8Mipb
e2vDay9WJgsIE9/y/ufQP6uHGnAeYo+mRxLh3F9rvSsyebZ8w0vQxvU/HwT+QTh8
nWVz5IiRRfEpMiTkzKHvnKNaolZNp5MbRFGvFETUbiiNQO0mRXREclgtvHnxFOGZ
SPU9hBbWhESyT5b8R8B8Ty6J3JkhHsT0COXV68Xwr4W2zuvnYcMyFBeh1UJoSWhY
FlVF1g8uCNQdBJIStLQEVfKsV+niJYRH4gorQpaTavNvlTF5uSLXFpFl76JWedQC
binSaOtYCywipry2hq/PxOFY6KblWz9FKGtIs8eJgSSP4W/0VIwKWkcLmgb2mDnt
srfmDT2djD2nUbriLXLk4LjOK9sllBP5PBXQZw3xWidAMe8ylCPd+6TLkbKqQwut
O8UJ9fSIpNUB4RBJBAkRhoOaKMhgena8ca0cbMNSDEz5g9uOAfNWHY4UoIL2mB10
xteREXLPeYSWGEItQQhrQB+UFUnd4hu145Z66ybfngxxN3hTDxQRw8Yegb8a1azz
PUIbpXHzEIj7MNcQnR1Y6GpClaHajbbdlxOdHRoebbmmxdnDIYShh37b0sTqR4GI
KwzulYL6uXwTmzfwMFdgMRu2856X0Td6Urk74AwutyIhecICnG+G6D0GiJgYs2zY
6FSJyWw22TYe7JLRbkq/bnti7n4R4ImtlUrxFvKeYagA7dh+cAqmZfLdtd4HZXov
SUaFBp4Z0U5/H0mnbCOrLUMLOYLVTyZuW7E7ICZLHTmoIIxCrcAvssvfrFMr1lkl
D37uIpVnKcZqZIvdC4bZ7+EQ/FpHgWozY/lJxNnjFiSBmbpOxgj08Usuq4h+1y4N
YxlC8PAzFiCbXD2ffmx6RjxDiAy74uz1dPH4uPgbxdn45cQgK87B6rgm58J+mHJo
TcVYLMuPm483gbuTRD27Oq1BK3B0VOnadzNup8iH4/oiBNzauuGtY6bn2Zj2Vir3
oQAVQoQKP1HOD95WtYUWb9yxeozvP/h8MUEzvbO15YdX7Tb2TP2XshPJ3Wf/X5yj
jqBXb8xfiRBKYksaLiKn29LmWZ981mox09+fTkYlXKhMHseqd07HEjjgYlfM8Xc2
Jg45NMCE4CfDm5bJLat1l62o662RtVNBqJkltVRm3GrdWjRUt/XQ9RlOxzJOPKBf
dUOBz3CbtRHOC7ufvaLAynbyrjaQwJJujOzWbZkBiXfLswgbUySN4MRdL0OdHsRP
DsC07DMDEZ5GMwga8z66zIIvomNEUEltWoEth7RGbXbXCWkxcqhabssXdf7qnUyq
ucxvBAuKr3BiiVfC6ivtQAY5Gk11lltYJejG5Wfxeu8/V4R63lCiOepiTm+VWbdz
ekbNLIG9GdhwHvGI/z/ycz0K2ubo82xvDIg68AEMJsJTQtUnLIAUKve/rdT40QT1
FHT2lNt94L1h+uA4h+EeAHs9hYI/YWT2Ls7kXyjlJbExPn3Syl4buCfl75/ZuMkg
Y+/1C7ldEBLDFJ2ooq1+0rEsaMHnIVjLwzi54XUN9R/valO+D8QLYKFFJl3iBF1f
4it12ZpXOBZ+mb652gEo8a6reUYbeABnmth4SkA/8OZXwpyk/e80ESp5YSm7tFXJ
a+ekpnQQHgYaJcS1qlDe14Bm5GjxixLXHFD7VgUhpeEBvIBJyktb3Dk9e8V2HF+J
R0p7ycB6gRa0kFIi1uViK+TJvrgPxkluCuvJXMajhy79vu51CgBzGMcdxJ5xWnD9
/PGwY3p4TuJAemtQn0sTa0hsbuRnDQWL9s9Gxw4z8j8uKKZ/w2WL7JyUOEMiEBSX
tPuUAVyHAnv2WzXOXRfu9JQUNVdDhfK6eFGuswnNmn1hOLJaAV04lbsbsMdoyY1q
BsPSKLE9jSnSGJOXHkhjI0Jjf26MtKXWMfgeEt9ZPavFZJo8Oe2oLL+dSwt7FCwk
ZgWap0J7POvRtJmUX4Y5OXsDJ7GpXhCtz9dd7oYENkOAbEnQj6LY0sXm8QWLgn4b
kq9XujCuSOTVmF0/fmVoeNGn1ecYyNZNMapqNWH1kRcZ1LsFva1Rg1gkBHE+jUrp
JHAD5ILCDn7tAcAiAyEfBrYFdFNmZ2grc+mByWpUfZxLb9CtCIF85NuLFMFmhOCk
WGHNI42kRe3svLOTmi05C3RUAnNjMgwR6UJgrkIsRuDaFwVjFBJcxM3189cVsEhO
edNHctBhGQ0ciQ8YiAGM4cNWqVIDSl7MWvVtlE5z40q9FmOUDCvurp+4VqfurTYu
aIaPQM/pTxbxk3r1OSAUrkZoq4OOmNn4/l0njFWYiKkvv3Eulz8KSx69mGF4psxm
ib7lDDA87diBgA8dOKhw/mv91QdheQasxFcYH0g1IGs1rHNl5xHU5eSJ5Cm1HvHP
Lvw3kasIu8XDSQEILKEAxqtlMzBgYBIICQERRiLrMVMhVfV+ZrEHoutiVWti6USB
EmrSfmtxSxylmf1BkmZ6nB5IturRw/vU+6zEYT90AtY9fh8gDHD43kpqgvmuDBuA
iXOHU2aFGfkUvjn4/Qvy3Wq8eQLmPRELkQ0t9i4Wl/Jd3FwTRmCtiikplQlYSa3N
91OOiIDhYd+R7Yq+uqJy9UYdYnJevwRdqpWMkXhzaC/MgVtGoLLeywHdNJjjUkwb
JaqhCo7QHjZJbH/Ly4gVN5Q8bgoDl/q8W+2PPpN7HXUritAvvFEXCBTwkc15y8aG
+h+HmGfYRPtTMWs+rZdk2M44C12uGmtP1BMyEFn+dQjSptOjR93M+lfUFN5XbA25
zBHRBX9QlpMWa0p54KgwgHw82e4o4EJDY3iL2wmen0ywcCRdIiXNGb4tquSc6ZEM
Qx0gRug0ri+iy/mwCdjbBnDWJCURuRaJvpWA14xNuw0L21JSoM/WR2pcWrW9sclL
qk/96cDzPWuDvLWse2SHFJUFjqozJu+oHxQ7QkOcM6uSzpGgR7F1sMDw+G4O73e2
+H98kOkQz/pxO7WnzdZ8rMGgSZW5GnpMaIhiv5OqwVevodMumtQ0cRvecy1uWnue
+kwdH+UQBkK7sCG2asw6/pafJecTD2AWwLL5xH0zZJrHcOtCurIb4d2IJqJW4wEy
dK9gD5CU/FvJVVXZkhnRMpqYwUYa+GwNBjFKHK1xl7YOAm8wg8SxjPfJHpEO4L6X
Zf/xLyugCSo0gkncfDOL+znOIsdN+W5J33aXd9MOl33O+8owhMpCLVSUuclLJHNx
+dRnced1PRnyc9WxnWF6W4z6Afg3vK4PhHeixlShi6KxPtpdNoK2xX8L/24KiNVn
sPbTCk6G1aM4B8npliJTY9mtwpG17QR7IkFA39YS/pUX4ql4KNNu0XZohop+c8bZ
6GSRPepyg7vZrJHC47azyBV1iKFNFcNGty1RhIeee3s1uXkjba4mMQq6QKrnohF/
Fe6au3kXVFlzDS4p/819LARHwV/Q5LTzviOcNu2Nw1gfxx7aSMgR7nZZ9stsfJMy
fNTIMKqbD5Wfrf72WRXZyIutbZ1cwOWFuDW+VPvtQ3Thj14pPW99wEte43O/kaU0
1JdwdcwAgzaUm6wxyaWLZ8WqywtRP8GddrAu8LO7ag3SR9xgaPDr9wYc5NmMOQGM
wMgdybWzVzVaiT4AzBSEZHsh7d9eiO+DZxt80nV4cWCL2pAoNvKmiFpUZuw2N4hA
wug8lvqVmxaYwAecNtPlnuh8kW1B63lYeyDsBzHxzmMVuwAefpWigOZ8BxNFoHed
fMB6x3h4IXshClxWfiTd0RHjLNJFWVqMSK1g2X/SuboTuw8Pv2qQ2SuEtScXh+3Y
1rug7IWAu4uzTIAsljij50QWoiWcNfKBgTIWBn2R5NFudYFNjOOzIXv4ZvGIeFAg
WPX4gVesavUkBNppAGs54JfmSvQGqxXV8r6gN0WqG+S6D61fAPOpkEK8llC5h8lv
PhXuIjSXT62v4HmsVGaNw4fYl5FQlmzNDi04+80bwzaSWTnwjYq3fGR3rjNsdZSV
9RVGnDotFq3SyLJ1/OLLpg//WbdnsjO5UKGUMwyZbQtmiqnScYokXII4caaK7j0F
Hc7I/ZF3GPJwxKKNmw22NcYlFARYsBC7NEvA5eJamLGCdI8rV9Qc5k2fJDdWjk+s
Yxo+nLotqBzWsL7C3epISve8JhPzWFIGw3tYuQU0WMtgpAR2uCJY5rwukHZli9QX
lVucIipG6dfJWSJkGhuelqqabl3jd7kIo8kW8yBnVPGeAFrugg4g9qg2EUa7P1Xq
yXswdv1GLbFHymwzcQXKd0Mf9Z+7r18t90XY+LwdgEi7We1aDFOHpfhA0bhABX/7
LVm8Csgx+JXtS41pLpeWk6VGoQimt8NtjC783qrv4LGm9aRoSOTY68Llo89c20q6
5naEgXAeBDkJITJchwaKuVoo3KVFGY86jPjc44eteM0ran6uyUPPaFsiEH8/C6EN
ZjqqrzudrF4xXuZFmsn4nDs+Y7nbjNkVgiOoaKCgIZjGtBJb7QZR3zHOtLWQH/w/
P/fQboU0d/z+X2Sxla3LUA4GAFTZQJ/enjzbm4fjsPeVOfrmxbRfM8rZ9IoWlDNS
QcfX6OpUgXZzcBIeEcjyqUZ3ON9bDbeVwAlJtXUmDWj1oDkE3V2UNiYHpNABbKTM
n8r2c87XeWClEZXktewVA7Jr3OKdTTsKBWjRqlEcI6ocGGZnll/OwVP8Te/eaT/T
88RfwIqvUm6RxSK03Ewys0u/ftn5wx66yHCKb1Z3/DaSlB5IZarqYVdGCvDtbAwd
Lkx6ww0yiFxphZvqDcjgTeD9u/LU6cAhvX3iqGw+fVQVuUJi1z3pibOFLkmZTHPf
L9+CNdUIisNoWfH4IYszv8E+blp9+GX3VBF14gf+8TTRk+PqxACOtNBnuKnEbBBW
U8CL1a0S81Jz8pa93WuJb4Y61gpdV54aQSYwMX7Fce9leYq0DAypbpM5mhJzAQPh
UUGSLx2jD5jD9L/Usf7eDXKWxNWNv5timkhq3KSn0lO6Er2YN974fgkrNvVMVgs5
LjqLQI4Pp26X+LR1a5pn9xua9wMpI654UNl/zl2xuvfyZbajY1L1pkNWkPUJpmcb
MExVvrBxZJjqHWGRXIDqLbpHcNrnXbZgF2+iUTXhoJcgbLI0uOOAxtQcrS+Xzb0V
3t4oQRF8uPuYYWxJ/CuF8Etv9B3ckG81iwzzW5XXq969aZttw5ccx2FPfnOAJZ/A
Q8UbNbQfKPFNKU54qruhYPW1mjtFfHVMNM+wlp5ma2m7+P4i4abVX7JMfAk837fS
ZJdI13aBDPuNm3HeJexlsM+YFZ8LtXyBwNWxbB2DHi6UdByoB6xalDwxNPp6YidR
uhzEMn/FboPX7QI62QNfDZGHMQrcRWs+NCs3l+TdiYyAfN/SneF/VNi/iMvq4Aj2
P1On5dZB3yupKP8wy+8Or9Yfd2OPDR7fx9UNttEfkHBMTXPKNJtu2p99sHaj51A2
22En7Q7qQtISmVDDo2q+lFZOEsaSTi4IKGcHkwLdp/Kr9PlBHXsxnTWaPV/loGZf
GWGRV5SDPhQXCBLjfkuvud4EOKUeGvNRnzlsrK2ceSQznYd81vxLLel1Nab7/kGl
yqof9M97XOxH/ioSrCw985tpX3j425RsJH/FGvV9E+3ZW3D0cLBhacQqwMXYmKN4
DUZRPzqABwFCN6o0C7HuiD67mX8S6P2KtiLUDMwr7uGgVgYL6nIBADaYMqDihKY1
FNNZYTw5s90Bc4x+EzZiJ20/BNiUFvOLAAnyt1MpzIRfxqgNEW2FfCYI2jvIu1ox
8YIGyKs3nM8/G8XwXz8IvVzwV47wDaYocpYEGuIISkl4jVE8Td5AFPU83BOweBUX
F9dQf4fxT8bBiU6wldwM8qnBK+BIYZM/Ngo5v2UhGpesd4i5zBhsPLpkwLrLAhO6
xeD4NekaVQgsP9k35vSVmPAL8qsxUkdJGXnAynyeMAThBCNbC2+9QZAlww4Cto8o
LVzEpfo40m0Uok8fQkTWpRM+96uqaw3lLYUKIvR86GGqUoY7fGKbeV5msv6Q91un
dZe85YX/o5Evanv92BimR2+XQsxXXaEKpKgz+p3Eef0lGq4G9CmPnVkG/9NfHsYl
ik61/45nwZMTa9C5ItRlstKkEHF9izef47QgDes2hn/wOa6gc3Dcaquyqj6QFq75
Ef29g+4JmeTETE6e2mIESrHq72ScjkAq0eLCfVvdrjw5lAkiFjS7/Ge1j/74ADAX
3Zq1WYyak7VPtyNYuzKkbAX5TlZuQaFFnObMjsb5sZG956WHANauu5DnkkZZHR05
8UCax/wwXoAueDbfnf8anTNujzraTos1BZWc5Ic7+tvPlvzG3l2qSlSa1Bjgg+/N
S+SdN9eou47ipJRYh5lxJkv/8cMX46laqKnfSH78wDTq2WBkFqwJmDhZ5UefXj35
3quLCPWjXF85go4Rs/iYpQd1+iub+3oTzx9N5HCzsx4DtKs9gCqVBTEsPDqXs1Y3
JPt874KRQr8t8uyUkJ8B9LVF+x1t+5wbqJEWi1Z9wqDudzZSC8pd9/sSDg4NUksK
c4SAMOFXabb5TgO+nvmvM0RjqjshSpZ+cHzBceDUeCEyL8DMZhHrVGn7WlWbKlGg
cBZ+Y1+ZIIrhLYooDa/zAsSGKMFAPr2hcpp0WIFwPlL5MH7mZhvkLfEy/LtnLyTb
MZlQTNuuBMHAOhtaLBVuadIpgV5nGGpmrPS2XISChG1/4kWL4Ax7tqPv4awPj4pJ
v8Uu7LwMk6S4zBDr+A0nsqVZISpiIIjWiWO1T3RtEwPT09dXHyHU2ukU+tEl0OQ/
mJZM+GCePQFzJ1XPNqBRC/4n2Oo/I7pJoNy//zdj6EW5orAbMDb5VgvDwrTKbnHQ
+srJfzFYXxKOQ+vVdHepN+kmH/doaHooWULQZmmxD6+az1nHfy4CbyCjhELIT9I0
0vcIG0nrXcKc8T/kROEf8etOCAm+bYcDEU30akA5jMza86HV/1217EHnu8K8i5Lm
tifMCCgscKXNwYqtlzjTC87ehmxlWgDDHMW5PO8euv/JXpiulozJCHLOVfuY541h
PlYuqTsVe2ZHKUAFjsCkGQ8k/Yx6dArMlckc5fUcLJKuXn1kzpfHKI2xuwbJew6o
AbioMCLaWSHz8mk6Mpo8Gx0yJioaJBMfA5bqReoLQt6tfHrz7NUM/IBRZBuLR0tP
PjmuwDLKzla/FXu851pM7kuNBkkDkNoklD/J3cZExEyJrD9loHEuyhmvmF1/zKsY
m6360/9T8Q1lGmFa54/rv2VNsrFHoHO3Z2PMSYDuB/+HDV5xg95rUuDNNpuMRojx
7GxeTaSZPXnunqkOFwbFaGLruWudnBjMlBh68nUybckeAZklzqRWq/gAdZYehbyK
2zZ6Hk213NVGpmd9O0exASewVqQ5jHyq0p56g9rihn6VVonlcTZQsKmYxRK0c8Mm
zq5P4vlR5JVvJqeoxZoq1+WjHlwImPrm7NWqYoX92tFYeEqIBqYZ/dbgJrDsmudg
2bbyAFp5wwFoL2gC02SaK8nmUpbH7Jgd7WYUiDWBHqA2UtNrPfjvMHLgRzNlFOzW
vNzivH/hh3anMoA+UmnMCrVGFxqq1M+EetkZKk3DrQEwYqpP8ucEHk0uyjfuvsKy
qp4aFqiQPuYGroAV7cVIcG+HNJe45xILC1k5mOjwZremBqSQbnL0UR7foq2taHHF
ur8jOKJGe79LAIZ2PqtrjL0A2wzc2HjnLqaPmpxoJRWRdtrAIuEibULx1UuHEb4R
1QIeNInBDyBskbOF2ydn09svabNIHU1e9QBMAerhK6nl4JTBcBvJ6LgLxgkm+Xpz
lF6PWP+WYFF/mnHhLVkLephNpVCWSxlSn+76qxUKk2B65VCmzbD1a47l/hNQ+k8i
i1hvQ4ZnjfiZPv9pmf08Ok2Wu3GTCdKIbGFMP4lf6g36LlQUoMJz/xycix6eOL2p
zz6l9FJaMgIWPS+ceZEcxcNMQcfDontlI07K61MTvk93VbalXdMKj0covUMMGbzb
Lyhm8vZyPbxjU6sIL358lXEMZhZB/Sx/rA3bEB519S/D1Ef/pT8TyBjawUKmWDI8
JdorKpydBq/+mtJN+HCco8R3+srRhbEO8UlkiSx3pHkJBUr/64nWHjBJ1fnfrzfc
aLeiveAxbD6HgeD3XD4qCGzP9ifqjxti4Ly59mibhHErTbyVW4FIe9QP+o55AUOQ
tkRZuZmlun6ffA91EIOZD6g8LlqbWdIYCz41CeI56eBMuGG9QVYXr46p1L6gWJOI
Nu0nykWU+lUKgLUtjOuBZufGKiNTkQpipwzeLK7LTeFExhtthL8TYKpQyvq/57hW
qSPZs9WpBcwC8hvxq4VU+cTqFf44meQIrE40Eza77/BfoPqcm4moQRud0m7vaiHb
k0l5b/0sGuTL6AOjSuQAMRqFmYj8/7YS+wK+rFHWyaCiGv4ZRkEy9U73c/WYPxdC
Bt2beujIOOLRtda1f27wjI8Wz5rzcgoVXoqwhb/eL7c/1wKESiCHZ2pjNKfOicYG
JkSioK+5TNILJBHDzGVn5PUVxSGdXLPrYlpxgotVLD1ZSwUELhYwBZCvTp4S7r/E
pePBTELNrCLvCUz83B9BZeObZHzR+ujvkPZ5bShMkZVVbbpebCaqOwdbsdh4HWSp
s2es7N3Z0foVDLoNYnazjdFq23IE5oq61PNuqV2whThhzZ6ZXy3KWFDqBN9PWqkt
udgBroeZZIFFd6UDHAYBdUsdMYRKYbZUpbxB2cIZIw3+G4eY/GNp/WKFSJOKiB+x
SZ84+HZ8Ku1eZNKhvWFno2Axn96d8wpXeqRfDYYFGpi3WamCtgTvokZzE+3KEYyV
TAmZK49CfTVDw/SwDDAUy7lzP9kwAHP2lxdcLU2qmgTO0EfqWScK6CbfmOg33VOu
VnT0K8lrRIETrh6Wd1R0CGJlfzxNZnXCyYWEbXYFzxEHijMOqfGFvHzPvL3vbXJW
a0XnK+HHJ6BwfduSoteopTQeigOu2W2qwcR9ApUinuws0omiDMkMnCQqUZBvayjV
vxXpsK+pe+w9NSXNnmJMBHlOY3GeEXJ7xqRDokwmpksQ8fUapDL1Vpzv6mYaYS2m
POsiuZezgtd9g3+OpdQ1s0CVwN4O9JQwpYU250Qf/0Zl51wVVKJPxOpD+Dls6SjU
LRBNB3OSrI/CzzbWvuMmKu2Rh4SZzPy8LOmJN5pbyG1ajpi0LYpMxAEyetfPxDG8
wsnwVy7psWGOcFgcpJlF9ERWNshn1O8DFd3TXnuEx5Td3+uA/YDc+L1MES/6NG3X
RdHQHNsLhmNKi583VUxDbRhHnv+4Q/8c/Q+F7I8Rlhtk+K2r22OM9sb3XegTAPZW
az4euHChbPwBD5cOWJgkDlFm+8exiNKZ22rAwmBs8WdUQzPYcWaq4oyfJOLOMyM6
I4tkrC6uySCqcczr0d7E0UsqkTCJWvZ/azXO98hwV4I6qZ85QEgmG8HlVheamV19
C9vbRwOPAp8cIt4NMyJyMbWe3clFuuAus3OKvINQ7Nh3hMDAUmKQCJPFb1+xaA2e
9DoHPKz7t79qJ16WRneCWPXFxVNpnyWFS4jUidHE4i1YoB55myc4l8jKWeaGjW2a
L9gEMzy/fZyVuBkbt0pfrrxWUqDXhvjoHcy3DIdin34E9zPsNy2+MXtqmaLzkHnr
wPV50wNDj2Ucxm7UyKBF6nBAXIeIzh0Ea6n57FAVhVywgq18b4S0cD7BWXDLLsum
3Hcp9myDIcVoRCF2wU/VzH9Zon9+hK9LBPJ72p8tg2OveUgByXB6FiWj0WG84vJV
D1JE/W5qUu4XoaCgXt8pJdIGAnskykTnQgcds1nshITUtdnn9gYmK67D/3ng39i5
/Nlpf0vNT9e/neATNiJD5ruvyc+tZvn5ILcix2nW4Q+d8D6Bc2okUFH9GCJKI1YD
z7u9/GVdF1JkGMWddZVDh0/HdOc6yp2eNUtvIGFDboMpJJWQRi9mn4yEF1YybmGD
INfl6R2+z4m6AaLtF4MU3Ihum4X+gc6cEPfdxaVDC13La12UPUM+Dbr7+Z+lZpAQ
j9vIQrW/rTZal0K4/73Fwjacll3JklhLP3sB7ZYvhN33kdkdCoNI2L9LQEpjUoxY
mMUPBTej6nd1zHjTS3RzR9afkGrW37zmkMYTn5HWbrZmFLkurmnFfy+3WE81LanJ
xbswC4GxB44AaoP2CLecLfsFUavTxWJtNZltK5KYeaZZKzu3vZSZiMu1ndGE7ln/
oWwlfA4+bR5AaWoV37IMgb9zIIblKW5eE3fXSjl8Ef1PwkKUNfDJIzLoxct8IVxP
qt1WGwGj6wZALuhH2fgx4+BabvbmzpWHWW+LIaXr5slObUvjB3PwEZnn+5S8Cdxe
WQL+EJJa3kILRqWgK2MiLMEBqTRmV5pr5hxwgb9czqMWsAfrD3N2+zY+EY8avHYP
cqFPeFtGzSoJBeyNBB+FCE5RM34Zxp5Y+uyeJMkpdxZZCdIz499z22JnZ2ryOIQA
CDnwIrzNnjT+OIpJq4QdNZNJGkPGYLesJGiCigcFJbU6yv2i4ERjGUXsTC8q/dyl
lTF4TvQI1lApDoMJgSp/EEZgeG4t79jfXIN8a91nGIgKvl7UZt0HPmsmj/Fik2z7
O6yCr7VTeh/FY569FcpDwWjFZ8e+oNoBv1+pDbSB1J7ArWEwX2T6F7FsHXckROtj
HZgr2nd8w6SYyzu6K2tf+3qUO38ndq5754ydLi11kdqcvQFjhPfGAzXQGsAtAkJp
jjGPnLHAvdZRyVMUNsXM3dZkVKWLXNHG3viTn8mgCGspyxq3Iu46uJC+7VlImO/p
tfYEDatWWNUpkDH72C2EzzDXo0XxtB+R3kCIWAhrZwgspJU+ekWw78BL4QrMWJKN
bfHKqXSwj3czI+csXt3zMBXKpHGgdn6VyHVVikJXqPq2AZW0mYuxeXA9tvve840L
iA65rQuSUWExi0z/3Y6IoHuFxi2GogwObIqtipytnbmkkcomKvXoRdrRCS0SEfUW
No0kOZv4fL2RQfhMt/XfISrU7asl/EKO46fKnlmo8qbTjkuXYfb1ld5mmm/QD+jP
DDTJcV6Dkh2w76a3GcPyOnbz3bhGm4BPYUrtcR18iwyBoG5E7TJs8D3Y5Q/WAtyh
frhr0Xunku+/DcNlEwx+y8rWYj5uC7z3MnXpHnLnKQUyNJsQ1HUJEx7Pmt+ghU3r
XLPR8gD0BWYSB13RXlKhWy7NGlQORPtxeesGDPtDpT84PaLwjwGjCsZmI+lnoL+3
7zq2YjqgUAYAk3WfbbrlC30YFX2CGB8i5EppkJJ0XntRrxkrQdHuJzElJYlFePDS
NMiukBG2EZafmUQYgM5JA8Yo6jV9q4njGZo551dY+MCliRqw673vLoyyj2LgsXZ5
TRbcK1FJEk3pYOqpRYdNH/BmxevAqTA8RNuAcvwrbLVATCIpkQqzvwLKLO5UkNGo
cwBH6o+P8d+3y/U82tGJzSVb5bnEX7hw2/lIkEv0z4q79cjc6Kf9q1pU/HDJQBPS
Dj00fFa3rbBsvFld7Wtc54oOoBN9/fmFAcAq0THwOr5fEWgHOnKPE9msSXT518Pc
UEOy0bJ3kAXedrLkkSgefKxst1kNzkeZ7sEMPB4b1vJEj6o3SydpUXwc16paG4gg
yXobskI5iDXb5eyc13nURwrhqh7gfpFVlOiU7z3FzkoKd3m6jeY+toe8kHDnjBVI
cm0asNTmn0JIIc648STrKKxqAs1O12mL+towx3gkp/txjWVzB9PpJqCgy1DZ7Mwy
Isi70GSHXQzHav9hRY+LJoKhQ6e4XwzuBGrhwt+so2RC7KnjnwqXo/Jevw5SYkRk
JzN0yzKIuNs4wjjNxBuvAmRHnHedChOoM7TpIzRjsatpA62g1YP1XJ8eigzSWP3x
SQ9Nesrbja6GadgQ5PRsNrqV70MyouKnqglsI18FDMIm6k0za5cd8OPomKWu8bRJ
SAUGtHtoL6/PPQqGHziWBC5imjMejpNuNReR4INYDdpCc7iGmJcFf6Hc2mciuSct
Wu4FXfVnVi8AEj3yXu+xg7qom4D+kWQSGoVMW2FV1N4tCB+l4gA2qRlFGdWvZn4I
24EbTzGPp74bpthBCjNmrDnYZ4EE/YyOaMNCerHWOf2Xtk+dLhQn7DfBgi0NEDin
Zyryy+c/Gnwm3ngfpjFFOtVccNIe7s85e/QZWaCvSfz9yS7FZiNv6KgJtBr32KO3
+rgTBXe7bBp9nhvQS8pfEfBAe3vMI8HFeygPKTRdo23LQ//X8t0U/zQgpbRhDIUL
dhGBz8NCdZC2Lw6HZEfaaMoZz/2+IrjJJZZFA9Rg/l71duUvqarAg4CcA0TQ14l2
miHSDCTEYmpIpwWHf/OM0m3t4s8Kn7hyIwIJ3vDwNpnVXylBhoetPig9EV0nCwHQ
JoCN1SCSCw2IpRMfNLPYh3R7OTn+t1iMJ1mmgwrwyfJpaV8QNbP9NnTb4ofJpjt9
Ah2lkG9HqYfcxoVGnZWCcY7S/nkn2nY6D3ZqtRv9lHWNYtvdtY82XCTBZaYp7cgA
eQ6a8mKUzt09PFBytDUPfIs8OMor6al1PSDCroVE66iRDsDinjKWM9jMGfMK53Zg
kmPB9FiAeHeaRUzZDkmv24cZF3W4PqActPq4Vy3eoicLPNTmzoizE/xZqUR/3B3P
XRg3d6UFhLRtPq3liZ/mJIfkPv3ZfqWkT+snD21QLirjnDV3kTcH2BJ9afKcVNNz
4Hx72ONG+qy+kdBUqpC5VL2+j9u6qJuMI+XOV7qXu6ZY3WQaE6X9pg8MrnajnSBo
nKxTOrIbV+EdkfVWou/gIqWfGyuY8HgyZUwkr9glZu/UmzeK42O0R2KITYGTGfTB
q1nCv+EStbYgGeSWwxbbmA74/BEWOOMbsrW9AqOIgdls5BYowruE2bG6Q9Lq00p7
grS2Se3mpBPpruSzXJHIugKU2bMIniIIt3fxNg2Q9+eLLWy5xSHuRvlRfiAlCQnU
p5RVEyydajcH+8BTWfHxfazl9Ofbh9JeXWat2/U9xTympNZXRNcIKjukV2CkooSe
vdmJMZZghzvbCEvHuwfhAoIQTuXoGk2brIEgauI1HBCmEs363wQ4i/vXb3qZEpUO
fSXFkwRrQZ6IkLN1LIpGbbY56z5ye9vS3/0zhsaolzVoXTiiOLoD0CW/fGBp6vuR
qpbYtD5Q7GYsGBo2RocwCWdNWcPHfMtIu1Zg1VQIk8LrIoSfygde4NzB+x3RIgRu
AmwFFehNeYHlXGamvN/lVecNbx6jBwe69+lydoTqItBkGA6Rt7V4djtP4bkjhhCt
Wp1Xn+yPRdby8+IGB4GrquuC0pI1CEauQsrF7s2DXCHT7xsH3GegFy2hG+C5MBmf
ksv6tyu93bKvI8XV9liR04XCINHaDQj/q+w6Utja8kDW0VxPWUJgMpkeItM30tgd
oKbIEiEVUdbBXnoJIj4LrcPvj0UVyBbxIUBqHforrvaoFYLMH3zRmJbPQHAIBrmw
3+mZvf3K/dyweyV6ze9dc5mlMtTA2p4AGhmL8ybeCKUmQ73KfVJSs9Z0X9n8foiI
yKvZkoLyQdkBUO6oA37Z1SAHwyyAkSzTrXu0USiIqXaC3SDZl4RYFhxRFtxNj3Mz
nbg+s42aVJVKEzrbPkuMfw0bEec95qKx2Mosc9fTFFwoF1wctg82RpNEH4n1g3WG
aYnCQ2jRFLe+4Y5Ntl4Nv6OhTRQBI+a4m310PPoaBrwy+AkujJrFiu2DI2yoI7O1
hDdOaIXXe3vWyycAeluPeSEeGocX3b9x8M1wrLqVEhpfaMVcq7mHG9FqxxvnKnXF
tdcfui01Ioo6GCJh4N6DV3C6wnRt0GER5UtfholYTs/tX3qM1Ph5LoNztQpW6f0D
SAIqqTzyZEgrkA+DCt5S+c6Dw+hABdv9NaRqZn45z7ZRofpl213+0AI8dNWsmpV8
p6N8dEsweW3PROxfl3PIfWwxl1pyb/8v0cUswgTQexvDyReuk+0flITIymyNITxX
bNx/XfyX5Lri7TgUBNvOvPwL4qkHBoxMha7o/e5noVn3l/3X3B2q3S2ia4xk8eF+
XcMrwwCXO7FsBFfVQGywUoFSRLCwEWncClT9NWeW5mPiHDL3876tgMN7GgVvdCmT
eIQbE8dhZsbK0XuBwpgaI3lRfIR+vcgA53QWR9OxZuT1I5nDBptG1dr4bJEzEB7+
Xw4pTpQRWvBb9NOeRKW/Ts0E/cDBUHDYUru5RBhWlISVTeyNlWstKqMABusziNK6
VZmipEQcAloV4eAGmnplaeZ8m+5kY+ghamDKvg2p0xQttilboJbYepdhbqi/UOW4
z8CN1SjEJuNw9W4wqHoDgudrWx7HNpspmHsXfYmyA5RV+hXKlojm8/08Kqfms/Ap
5qa/LuXguYTZXGgsayEmC5B4jWFBhtXpmy12Har/k1Z4V9KERNi9WqblS87DsHag
zKMhDAg/l+Yfzot8ZTX4UR3Swb8bgxtoJx6LVu7Ze7B/aaqhnmocHOrE0gtR3nTT
LT23iZjVo7KVOxmxkeA98tP1aHrdin9+VNMeFsJU/VQ1jFGNco+B21ETWWkIF03p
RVXnf+qoeyzNlsPbAg8nixkQLcyQVWqiGWHVaJcli1yqnbpNGIv3HuqL84fri1Qr
3m42yCHEqIrqJ4TccGZh94xLLJmiueDDDGHb56lsw4KD+K6Hmh03dBxPDr0+aozD
y7rCgtxpSlL+2+2xVJXBkHP41E4fYFOfyqZQtzd736fe8lTUZbH894ucGyNTGggS
V/bHbYJmYYH5F38+s5FBwnwOdFhIbGoLEVF3aTv36KR5BJWMjnU92s+/G6666/4Y
CWbL1JPrxsEwX+/SDhuoT2yToidM1djE4aSQmDyGOeaZm2nsQ918uMgxHK9+xi1J
tPz2uJjfGq5Kgyk9S9n6WFSREliGUf01OAeigS6sbh4ct0QG011LGcr1pKdH2ilu
XUjXOo0k3QAFvM5Nn0fOps16+yLUxy0vgDc+TXGM09IHSBQpmOIuKGY7FK1HejzT
XatCmL0/Oz9TmvYhX2MBuGBfmoLhWDEGyP4NWpSO6U0UcPYARvzdwUsuxgW9b+xI
peuQ04kk5cXtn2HJ2SkAK7uH+mITkyigD34Tan3udMw/45JbGJy5ehXvvka1xOP6
YKBvLYbz0L9NgEDeI558LSoGJQdoSNgw0f0f3IOLoesE4DwADYZIBlOn4nRfBJOf
7JetmaAsIAJfzb8x18JVUXpeezE4QlIfgImqRftgJB4is0C5gz2bbSzbX/tQUZGW
1++MeMq13H6l8wCkakwpxgcGAuT68rLO4D+rN/oAg+AuHXw3eAIPyJBMD2T3PoYb
ucVVyewhzB29WLry9Ipk5S8kYm3hrJL47O+FFMHAaQs9iFELmtYRnvJ31CHBHNUL
jsfM97lQhQDac8bzQPZTWiszHK1gvVZtXQXNmfYcyQLIFVp6XdGblfMVWHPY+t3f
538Vo8XROW0GMTLApZLxhCEoTLzbf6u5OFoBAOJFb4uLDnZPQ4WUhxMApZmAwoW1
RNokwOyVN7VyNusMYprJe3AlI4BgHp5aXj/FVBryNSDN6Q3mUmTG5FShqmmLDb2B
zNeKEJKx7Dnu/XzPmHZxKMScVqrofYhVUcLlEyxTQ7YQE+gigYtTYgmO7QY9Qw+x
P7uJZRtsqtU6StsC/Iqi4LaI70rtyUiJfVKlYR//YWquaUYVbbEWFi49yqcgAoNP
tOA0QMqbXGzqweOuNQk7psWCk96Nf2P6Dr9XmQmx8uUrbW2PV1YtVpIHC3hNxl6z
kBQTd3Y4mp3RamAWBTqeCWWX5RNHNkEOKH2jjtiYwXKIu9ERQl2Fj4DgiwMflGbC
uZdcNITRHYV34zSoADKpNthVrusBYpfaaDiCLl/zrTvkfHR4KKxQkHsMJ/l3fTkt
+A577KtbtPlT8r8Bu4f0rBDLrP0nDFdmfqx6wH62Wwu52fyIlutr38Oc1gprn58J
ybEN3QOaC6HqT93X7MUOamUBBEMGLcj/JfApQTFBPaMhElDZEZC7c3NDmOajJDe6
0d1Y3NHq9TB2Xiec4JoVZbekVb82tNlfRzrJAt6PhjqdLz3scQ7lYVZAnfmZ8mSO
HLNqDEKcgrKXb1D2fGlISCQ5NXwUqdUEH/nbjszTTm5w4bKxWVBMY4EPCAHmAQny
Zbk4UWOwXG599IsbJpDYRqQ/KWCQS9JNHQModPE7mDd6Y7/h4xEGFewMLoiOuDCX
U3UM0wLGZ85ddCBTKcCiCSgmA69v+gKL/BRsfr+01spnEd/ylpYmMFhJ9ot9GexY
4/fkdo4ZqHJ+jQX5T0kA0zZepQmyPEWIc0QeWmjeZ8IsDjgO1Rr/m/DKty5+vw9v
66hoeXlJQVWJFGaOYSKHgxC4wA0D9NSNxdtsDfez/vu1VKjDOdQrCNxbadkO3RfE
LSF5m5pHep3H5d7i9pNHmVoQnKv7PHLXLY9cULs7tOfE1VB3xnIft2j/yLLT4w2R
HVdxTJJHlMquPmzbNKpJZ7OfCzQRbVnhd0qpwMlKS+ijEderN8K9QByXN4/EjVXw
1SmV38jfvHEYT6PL6AxNMhBxoCuDxg5uYX8VZsQkgsvQjdhI6kaKPTx4PwZpFjuA
PfgKG/KWps70TEqbGguzNKhFhfmkCkVvw1VtO+Tdgol4WhxKQRmkfuBQKnYOop+X
kRZBsSMSD1VqQicSvWG2EBcJJht6gigOUzk1att0ex6RjiUCUz30TORObnO4o5+b
ZfK0CaJg5JBWvxfbgISB2BF6LV7f4zMvFfRZNrhUuzxVR/w2w24iaph+aURdcMMZ
q7eg1UPFqeF1Z4CwTM/BpSnpCcOQa1w63sBKJ1KAK7OtNmA+Bt8XIIvb0fo/i94e
cVvK97JYQ1JxXX3BY74H9Zy58M8L+cS1zQTOvNhPaxNY3RIM+MUYRqvM6/0Y9p9Q
deMBfEuup9BOsVKtfwamtx0EvtzNkQ2l4Aq9eccwkjm4JUtEi2lrt8Kp7yAdCf2t
hNi12JqThcdKN3E13CI7v2breGwPKe2RNdd67e0+fV4yI5ku5PpNm4iaYmJblkbR
frS9DFC4flrw8bQmKtmWJyIbDGaeiIAEELize4yAi602ek3rAhX92sCCMgbZOOPO
UIN8iVkG+067T5sQy6Sx9lzT1GU/LaeyHVp11YO6BuNXCKrtqxlvjAFPRa1B72hq
+gj5YaD1JnJITHDr83si61wHWVLescMSXNJjagDcTz/GMqD1w49PpeVBAdHhN6RR
p57C7RL4oZJmUF5d1UVOy2JjETa9ms+RFDlHBOd8RkJw8FvYlhWKfa542+ESHrju
jdOQKEpA8PrU3cZ4LIug0KgHC57JPzK/GU3hO8idKFv/Fr38DT7mf2TNUP64/t1R
cmrW+3i2AMn30KTIkkUKj/yn/4faCA4MOVyllj1cIJymObHN71mRvskBdPhM94rm
zRwRyb8tI2+CIH51zmQNj05ojZI+zuEzPEhkrOeRHe50FR4BtHfoABQIURS2+BxO
8kOkjN84DPGrxoSE9rupNBgfaw8Sy8o1r+bp6xNxgMzkR0f6vDogZyz8by6nlDLY
9VX8il7SL8NaURofwoLiiLrytETHD+7vHEPW5Gb05kY0ZMTPqLwtCVtCAAZ86bA8
nyFJLJfB8shTxpfubedu+DPxg3LaTexzh0HnXPF7yr+m38m95u7Z3Tan+S71ytA8
+ZfAr9FlxACy5NptWVvhzUSNcWMekf6kw0sxOC3wZU/KqmIDlDAM8dAIZovxvNJs
pkiXprA/qNSEVCbMndJUjsmCiRL7LvZNgJIu3i5BjAbHm3RMkJQC5wBoaynslru7
UwYen9w//SasW43/0DMzXIZEq1PzM9c+1XD0NYUTNhruoH//F76vyVEiJPe5qACJ
VK3FVNheDKyxXbX2mK+GAvaDYeIurztg3r7eMt/Ru6H4bPE1K/nWlqlchduoJgy8
2PKgK5qXuxc1bhIwZMZISZnL5EaunJuMLrcL7HFOgDJ9iGt1U7SaEXSQLwuZsHns
7yzM3DJaZqvWy1KfB7rvMcg+ASpkCsHQm8xLEJQ8FwWruqudfUbbIZ9rCER2J4VL
JPpAL82E2leXWnCXpVRrjaiqReC6QKZ/XIVawBD2mrZVBrcg4C3vrE2P8JhrVn/z
JmVvno3hjNeEOWuMJWltkSjSp6lCHz3YRvk+MP62ihwdC6lGBItRDRyxvoQbsRat
xaHhxmhTD568z6qKvOgqGH/6l5xnYnLXCTX9fSNtWkA9rHmBjET9CRhHYJ4lqO+z
z7Uq60+2hHa9Afy4+KcJAl3Kjl013FvPx/f6ZVXSOZQq8Cvou28KBzJNcyriAB5A
Olbvk30/N75JnlWOL5xNcTo7YIE0Uf+aRyQokbVicz7fNgqgHvDCnMOLbBi90ZBb
uYh/FzegyzLpEEmCqqniHkzucwKzhyyodVD3E6Jbp+FpJdDHnK1jyIhflY8WJ5Wk
KD+D7n32QmKzWrqsex9cH8txJxEj6eOvzqVsGfEIqe7a00weGKTfy2NNB7z7EBbF
0NRo42P8sWn4Y8rEJI0GSOxSn5jnsrET/KajrCE7bH+XG8zQ2cMslUjO4CvuAC2b
mxvEZdzN2U/+hrvaO/V8zxSu25erAwRDN5zXKF54P/s5+e30wes1yRBlgiDdgywr
tuFp7o6NFogblJJ+V1jCjtpZLSqkB2RmxwuXj8vf7ZS4eUN+eVcWyuLPKWcOTSyB
Yjweg/Jq5m5SKORzfd0GDNx293sriTQ08Lb9Jx2z5pALaoODIhpQM9gnL6A/0Qwr
AzXcg6cvoXzlZ5MdbQ9xEAtLjr+D86vKNHEUjL5sTZTstb1NbolumEWqF54E6SvY
+dTXqvTJykmTCkAAH9rsRcGv08mjBQ+7DRYm9SiRcry4vkwX48DAp6hcc9lGkTQb
DkAYnLAMTx5r8oyPxnMGI07sO7y0sFYiP7em6uES0Vio6fC6hBo2tPJiZF1NJDl3
pEtAS3/MEUf06l7FCTugVUDccymU1uriaz+ZrJzwz+EwaKzi8Ab+xZ+QlLpWcXwD
0zwVSudq/UxvzDgY/b7a7AOEWfVmMiEpBfcspbWGklcj5VPZ8UXRB1O3/9+ywmz3
60SPEci2EEKOCJc8nbyrNbY4lFmsqYOdrkA1Je33q10U+z/TvyoJtofSBC1ywdPm
kUacdRx7UUcB4AU19v/ISAM43idqZQyrIuJmeGHJafTCEOBggUnPtGg3QaHPedDi
uV2ACCpIrGZIbqcR9oPStS2IX5qPSuCUKr42I/J7kU6QPs6OS+eTEANph24e07a8
Y7SUbjz/P0GH1/q1DmH4wuaQSkTxcULz/S5y5s2rtGkSkCjt1mNM/YHP5Zh7pRyV
Uc5UpGOZEt1JQ5tiDs73FD9VGhiSuR9qhR2vLaD08ioCT5ApvFuu2WWKwPCnmYni
H8O46R/g0mWBajCR4Hbw0aEVs85C+rT3MUKhzL3HkpFAvXWGnHDf1gwPmudWZrds
qxUKybVzd56EbfOHDtUZCdHI49fK6NqmYzp9ZUchd8BzVi0682FmEeiZGHWvPn3B
KlqxQOzKxolMeteGNuoFhzQkrBsTOkgdMBy7/i9D3pp1T/fQHX6d3LhhxuDCronN
A1YwDSvpv+T6j4enGFbxjeh2nsZS+ZuJNwPHBtEju+3QDBs+X/qFggIaOyOWcsQq
08gxXtufoi6K2FJGfcE54TRfUWO1e1dlx+Mou4y+CPX/OgU8H9M8q/PjEO5NYB/T
2Fh/lFa/SFYcNqCNGpvCz1m1jnI/l9OWonDp8xhWjnqi1yv7rhCOGtF8Ck/695du
jl9/Ukx2fw/bLPRpoxSykHwvzmIIqr6VeO9h6vN//11q9m+vvzvkq8v29DkUNUMU
QQ1X0Y2VBLVhIjEtwe5boCiL/LRV2QJ9oaRwQHK0YRkMUAlfBipp4z6Jbe0v4wyW
brsLeap0UL97731KnIxuM1y5yJX2v1gKJ+7muJX0U9pGKBF5HaVbaenWGwBehvKC
oM/ZcpgtpNqFC5uIcKctDd5ja7y6ZiuoGBQCMicuJ/d0ksfUZBG+0lVLFxmOMzCX
X8CgxKzQ1CNOWbj5hqMvLWQxH1q7SppGmwaLHi/Lss/PHowqerxL4XPNPxgxStrg
VTrNwnFV84sBw+W/nNdadjyrM0VASKT74HWmj186oYm2OLNLEtR5K7jt8gz6aVd9
V0So6yQYsb0hJVzdaWQPxVbZglE0pczqPBc0GnridnRGLDY+rBjR/q8i49qkdf4/
XwC9cu8cavA3AjmbAvhx9xzH8glp1lFUj1+2NWNzyRCR8yin9ryvA4nR2lnY0wA5
f3ZrgqGcb3fhOzwpIxyvXH4W+660BjBMK8trfgysz4fj1z+77val7XwCkxbjhA4Z
Jj264Qeqnxkl/T1ITTTL+b5RiRcWPN4w8kxyLcsR8sslWzpba+BZei8geXI9vTTH
e2++6+vdkpFqSGkB8XwwSdfjD9OhvJysZXeuDQLLfOy4CuYRi6EK1VdI9Udw6WiL
YZ9SQ9Lmcsm4IXVXqOjvOUtJxeMoyr4eLXxF/Ms0lZhbTQms2lIcmLciWEjeBzQ6
L40N1xIh59pGX++WdzrXYJJbdVty9zNTePpgFRyy8Xc/PhFjWaS8CPuKtPD57YrZ
aiCUwcVWDGkxXqaY+wdi7JjXYobSVW716MtX5D4hVsFSCSAHYLhBtey27dejkicJ
oXUFDrtmAimGSFbE1AP5/UV17+CW+BxdnjlMMXnREPc72IMX4FmJaqKhKgWQZ09e
xBpgebuRp54vgfgnf0XMQg/3T3AB8jMXH3+Hal5LZnGJwBqGgSXEkgFMhp/0xf2n
mpQ4FXfM1psKJioizQh/P+EglvEDxZQWuePeGgY9Daw8onftsd2OeSPBRiYDPUjq
YdNRrkUup4SFyqvm2fETy9k21y74q1JxyBJM5Nq7UXsgT+n44F/j2nfVwBYUASJK
fMH1QZ8pEF2PzkEoVNwaoudTOv7Kk2e2bcW+InxEQwIEBHoAiDons6KecXUoV8gS
Gps5LUAEs7+YasAPEuk59Mz328qF4gMw4IIqbshSqYXl81116Vt2mnflxc9zgVBN
1lB1D1JZpEHIxSXzfjd+/88rUgmTvbMnDwHc+0Duskf0a/W9yRamk8aAiTaLm7Qd
LIG42TfNMvoNwjPeyz2LLfZyT3FDVA9JkB91/InB+pY20+vObdYhZgjQjCC8ITVK
HJynCTREdj9Pf5LimuLfESTbEfMNumzLZ2NTp4tW2VhBkh2VHR2qDdlLkVcM20M/
tKTKA7j2uOfJMV8o34wBufIv/IbxFYPpxM9GaF08QgIxN0v6RymyxTrF2fWUiYQj
Smf2hk34OjETGZllBwqAGhDNQPbR/S01ZFZkFS/S7px2lFvQHT711jzzcSbICLYs
phk1NhpapXhPu070TmIONsl65MMo1ez4r1QAcyjCg2N/TBmsUI4ipIiurOD9JLQ3
lBxazDL/nUjj9nx67Gt9xn7gup4VyS9syGqcpbgbHpURsgh9wVZzJZASGj5mRufH
LfbkD7dpp359i3Zx1B5ZO8wO3tuRrWzJePz8PejKBkrtOcQcoqp8+w42D7MLHE64
TapuA79AyaGNbfguQuHUGJSH+0W6ARHQPaR9vuvYRYNWtufXbSc/XEy5oq+6X07N
w22TZoy3U9YrzXfi+HQNmyUj+06T24uX5IFbhYFOzkfKNPU/Ut8tzPGsffaGs8B7
i2C1gc3p2/d1ITEslNBsAVn9D8Zdj4N3BUIY+0prRyXnHzm133iyXWtZcNM+9yYb
8ZWEao/ZFxpQpcgy27tjh7chzWiXSmWE+HN4KAhVmVGsu4t2kaxv/oAROkMKk/Am
z1L4YtdEdJ7wNbBi0X3at7pYKyMB6Vy3IrfUqoG3s6rX1+d05LLt13pae4a7wgz8
ql1ZKJESJd4ojsUYFgvOig8w3N+PsYxF1rQFnrB5dxbx9resMHGnVDNibAaljJM9
qjmYKKNiAH6Sugssh9pBDgd4/JYzdtfezGXCU/96EbzhiWV9L2d2QuLVEcpqrD9T
AV2G+KcuQmgiD+DqAMN058n168NOcxjgDdHjZNFdY3fU5ElQrILbfbX0Vl7p3VK2
gvW+/EsMuEXGUS1/Qnab7oGkUMjTQWf47iVQ6zhAJ/Ea2W4GEp3xD9zTXRbfThin
DZLzgfnA2NV9WJTcqHKtXi/JnaoCfW5Fa9jz33OEdbd5mnzBfhe90quoAB8X3sKM
9Y3JS/9WOjtAPdvRTbv7WeZrwnWS4QckkLCZIiXOowWRCJc717tVIqtauNtl0HnA
TWi9Q2dJbc3RED1uMSgyQpJaf5WuvZF8Flukd6+MwI0g1F4irjj02ZtLRwXQiZfK
/ZDvyeiSrXXOgQHlmCGzjrgARnbLAPZDmoc8erLj4IEGtCuip5mLS7ord4LTRx7o
/LayDKkNRLiyGb7mqwneziQWYqUXzjD2Qslx11b7iZwmN2Y39YqF0Y+zKvbrTeG9
Rf2X/rE6nqhMEzzSStowNElspOMCpqQR8fke4nG0GwUhCSvxMrogY90vKdSUzMZd
dSWZxruq+LlheI/YrmPcFJj7qXUKnpgCeqIJ+SwmLH5BbFQ3o4yL++Y0M8jnYBrO
0fNHAw7a9twBCCherW+Mcc7wQeGn4ywyBR/VzgFnmk1SJh9EZvssBkTAs60CE3aN
MVxNstd+xSOr8QmdhLRWBiY/Qet40I0UXUF+TsUN83LRKob69xhor+1pNUlCzDu1
67m0lqayjFzxsGh2JKDl7X85OrwU8EdcNm8V+RHpJS8+FuZoPVR8QvPChh0+5Bh0
FHpgn8hKvsFtUY5TxVW+wdc7IjoV2ptP/0Yk2obFpQcwpRq5RN0LWrP52kf2E7MI
uq3Lgd74TD6kLr9smE74e17qBOU6CCfTKhQoFnHpNzVST/wUoxSIqILsf3tz2JjC
gCRDlcMzg+A3LiwEjo+tsO2MmHgLAClsxWQmdfbfRsr1jMeQJupwsOe663QIU9YU
uOrvOPEtnNlF+3dJ4LdA5tUR9TML4Xh0c60KEc1h83f02FP66fv3w3CJ1730pCqC
bSgSm6dXtHqY4w8pfzsDn7W8zvqqRlUDWNB8fKvFoKZYWI2rylvbo/o0kJhGrgvC
GnTOJzQemw/xxDEk4Uvf+L7UlyrE/arU7pF4pN8s2F4Q21id97HFfHSzGDpDxnjD
SicZm4pQ/0DdkiRO/mLGnL3NxmDWnKaXGMudSJjKWKu9qepw7/adpU7A5wH5WIa/
AW37tnuzXWEzH2fL2hxTFj5EMAYSQnOAmwbWTv633yNipHMvqLEw8Eqt0N/UIa7i
SdYzwryTv3L0OgyQsazP2XgcgU6KjDlaHvCAbQOJe4KdyLV4rdqWx8833aB3vvPd
Kg/ntZ7UFhSjshZ9n6/DcrS9ivfH//2q4IQdMYMcjL+8tOkYHAGc2dkx/qb4X0bH
FpQN2inXkfcB3AyL2N8abPsXvQlsyzIQB7Arx3uCgEGgvopTpb4bHvACkH+f4hEF
aHYgnzVFglmzjyq5MI6YQNUP9ltOrg9WIOEsfsa62nzz9u+Kpdf57z3KvExg0uss
afjcWLWAlHmQGZFKpsKoopc/r0e9S2Gx06kpOFXyjgQb9q/n/GtDzwUqidChoubN
JT8B8jiD/yTZyUeIx1Gc/7p4hMSolg8a8rchrisXcvQssNdSf7zG/EbCRxJPFTMW
RhNuoj7ndLb1FTpeRSL8ZrtbDlIlcMzb7cXFfKWkHf5r49nWfPAnhhfR8Rfcqn6D
t+gckw1X1pNkQjLKu8Ju0XTSSoUIxbHo4pB1/0cyBFzS0sqBuhT+1rKTKgYng+MG
Wtl69yOP0pJssQvhgvbEqaact4+JEJsxgTY7VMAEC9aee5+smnQpuapk16mPFgZ7
2DRCbbucQudw9TyXpEep+RX2e+Cfol0UdFFA30qbvi4HmvNvyoThnUogYr2Flsvx
QFgwX60BmOQb08AnR8V++tf/h6U5gtoxwq3HBGimJrGiHuxJuEukVpAjumWMk7A7
XVGhJSKW8gADuZ8O8briyspWfdompDf3SSMrSpl9XD7nM0Nk5X8sQQQJf3VJa9hH
3AoJn/fury/gACySYYMqXy40bbFHyn7FOETkiGwrN8KPxsM5HGdMZH9sx0wlUC+U
uj7NAW0SmnueU8Tyksl/FElWlsY1F0lrzqsA/Ih0daKka4orL4RApF1iGxoZvAX5
3DC8giUuJMl2QWVDJB3aA47XGRnYZYxprWLkVrCnLI/GN2FuurxY67MucAtQBdzE
MO04VEl4K0UFSkh6czvmbl7gV3VOdsnd+e3ewQI90e/Nl0aRf2IVuKkQxh7aymHC
xIZWDkqPLDfTOt4NwVxhIppJg/F5tt5ZujbfVIw/v9tmNStJN0FHXdBzhwsqa5YB
AlNNtn/4RZr6IRUwsWmrIo+wSwMzV8RiAnqPr4gTW4LWzOxVv2n9Sk1hszla2a8a
jxR3VP6NITRVumEDzmIAsBwHzBRd1Uzz7ULVwX7vhnz5cacjn0wuJ9rDtLSo0Ttv
mWHukAtXSYkZA3FJZYvpO1Z4oAvq9kFAvCQM6UKeiC/zIaZrc5YEAtrneqKG990E
ye+p0k/0iauQ5xaD2Ei3PIkF3KklOqvSg1OatEUhRRxs5a3JcBxFhkhxqz/9AwPT
+B+Nbbh0cbgnSzuO03AwelcC79zy/wgD93EL58Kva9hPyi2kZevTJf85BzIpVEa4
g6yw7gsoC7bI4yy49PSGk5HFqITZtTdlW6Lwd9/U3HoKCQhkaXlNVIX2+8riHU+I
fDQq6Xiji+z3cx2wxocx/skp4iHk/Bxsk97zoQdg7j5gkECCz4cW8PQ09ckkC9XC
aiDN3y+dklaptVA8Ra7k+aD7JKDlD2ZJWhPNoceGwmbe7Zdan73SAcfmOPex0X2E
NaTcL9ITDpiuscgyGPHgn+4fNayPGoCxC0wUVVlGbU51g/TnGGWxC9TiEgwh6pW5
jEf5YuagpfW/BBfXUG9A4MRWYzrgT7598ZFgvUXHwJ2nFDbsfu/PM48Ym4hALwy+
bcIbCxc6/19ehsWsp/nFTuE7mSzmurMExDJmey419OuQb/Dr+V2ZbKuTER8zWEw/
KuhIsGz0Z7H/cM9kdaKXCZZ35buPjX5tWtSNA3m/er4kLCemG1l9TNrwJVYa4lKe
OluvIkqDSGRnylXRdQf1F4q3an6MJnTt7OArboZ9kGWVXbTsQ2mU2DvVoQAj+vgp
6ww8LLKD5DrlbJVe9rpXSf7pe5gj3ZIdn+OpYXLWvUMf3KFDXrtcZLmjlDF663pS
p86RqVYsE4q4bEBHzt7IpxZH6ucIWdeyp5y8+kjpTvbjWghILGdCeE+mH0z2zfF3
AO5fHRGl8s1r82WWbFS6/7zOStZY33iR6JY8bm6w1IrTxG7vyjYgg57ipmgEgl71
gQ1UDge0RV6KaLVLq4X2A81OjL+rPr7B9tsX3hPFq7CLG2z/8Nc4TLeocOYcQfkZ
CMFWTFI79CqjOUV6ZAfSAl8MVQnRUAT6apGIgAPApBi6BXGqZAkbSsNtdnPvJDSx
4cghHVUJN1q2iYTDFd+p9y0IZKSzXUPp/oh/lI4TxyHquxgKGx0Wmdg2JWEqwf1N
0G2vBeG/CClxagpJSLaHaSimI68sihEJ5Dh/ECSLQOX3ehk92o3jHPKgGF3zke5K
jfXQSLDFkLeOerpjuOyk3X4XEGYnp4ULLuh1wqwTH8deHlmZmVIwqtm0roe5GHFL
xpF3DzGxyKPw7FcrfrzW7zpEsrrEpxE+LuMdaOwjNh91jorFmCVq8uUHvHYtNcmu
M9HKpxB/Nd8eFV4yoC9x2fwGQ3kJgJRw4gbcGqfvrQYbWy0C3LknQMFXtU24lbU2
7WsPQj12j7JE5gFR4YANKai/tyNp3kCbryp8Pr5305LnqeUJPGOmmyjamZzQUC19
th3aCr+82kMjDtqS2geJonOWxnp2bwbcSn/cAHl154TtW0YWlROHqWtjVVbq3GS3
zF4jyeQ1FlWn+MK4zJVyYSwENXxWtUCYHI/LNQ1rpT80vpBmNYPDMjokCNDmcc3r
9CF2IzP5zdVxmMUZTOcrh2Amqe4im2KT2+vLQsP6Bn7ymncrxgpKrPRRDVL+7mMJ
kJR3EOAF4HHZXfy2XOuxBR/xQzi5yJPG7CmFQHoegyL6seg3W6w4pxpO02x+gbvn
jdeuZG8QZN9K3+tsPfxA7Uq/Hjq4eg/DQqhqa4iV7EbLu1FBcvE0MXOop5CFmklz
uSJA6n0Yk8+RplYNCzdw8cTB1wMvZYWrWAegj5eu/p0UVeMb5jesg2Rc2Ye2Ckpt
hKkupyagQF912tixxatJGn5zfoZtSIkyOcfG6qi7BqHG9Gy2MzdwBzPgwI6OZWly
GwJ0Y6K7OxniwcaXwsuZBtLlgyLiIVBbYyeG/rGplTR2hCtYav1tG+XrCFneUIUY
+t74Gt6ofZYEQzFmx4r7KUZ/j8+nAZj6TbUXkKAvpVqARsAPHSReZaPYXqyqDibG
YeZN9J5LFBMPq1EI0ICchbwC/DIbcil0nhr/OgPAU2dtutp/o4CbZNA6Hl0hp2aX
snTPEqzDRKXnhbZ7tNXugKd6jHAfRQRKrdKU3jmKPtKaNDNrK3v5F1bgXqd4vLOc
vhFNroAhekBOB62aRmw84syQlHsU5yOA1J9xVRjautDhDCnzpnV0dxWB+awY63yl
msiQ/8NfrHzzH0t/kmfq1HJXCuO8zAgdHOfETLphzPWanl817daTpPbtE1/WfVZg
xgr4dNRqDpb+vZTdctdRekuTIx5d3j15vfDp/GrbPAC68q2ZT4yWf2TG0nKnRd9M
+RFoNhl86ArK5kbjxPZQ/6CEFhYoR/QdAONpMNbyW677jomcZm/lgLmjhrd/0xXB
jchfehxIQoBT9uul4Hm6RM1w3RlygEyKU1DWl98ccFxzIjdHfb36mRDlbh3/2Rw4
bR7u7cdiUFY+t9B2ZnL/Gkc/PBx5baCnIh1odMbB53UFWyw4jdT4FtxtRAFV4xNP
O95FehBds6T+AenbzBWolc8AccCWcQOKs+RPx4LN9CKpQUGw3ncJ25AqC4TFhWcA
KDrL3erWGpa+MWvLfdu3Ywz50z0AtXS7C85rcTlKRgNtMlXnsE5melokCC/fbAFv
+kpAQqg7nMXQ0sczL6mvoFFO4psV7JWGNRbmQ3iaqTDMBefK782qhrWB7Dm/6s2I
PruehVF/0xrFkKcnlocvJGdmwfRsc6QsIw6ajt6AHpmeEMFkzRuzZemvp6RkVgza
Mmos+wud+FVY2or24abrRyjXn9LqgASHVbdUUsbpwJFB/8kli7rD/VGNwdGSX9tR
c3fW4rr0V2mEilT05OofELQbMvEN/LSSg2KJcKgL0ZINi3GHEl5yE6qodS3km9gm
WKrm4GBbQu6g1uyvTfhW1AcvFzzqYOjnSlfLiEABzPnUFcD9u6pMfKCznKrkk1Vu
cmSkZ1g0O4CW6yI/qmoyh8OApssCCWGqwd73Hxq91hJtPGpoeEynzhXFTVXODvz6
6EFhHTaRq7T288dyh2vJFA7W4evDv3WH5ijdUjLUhgvstnpYf/hYP4aA3xTG1GLD
2Lk5dc7C7KhkJEhNQrHssRKrl+/YkWmMF7eD3wKW76unRZ7YMQUv/WNKTVysvjLi
RTilJ616GS08pRlSQcytdHe4VJZTiP9Pba6w/w//+y/oonl20UpxT3p2BcUONz4T
3HjmlaKK0U+StzLni9eA+45pEH6VdK10gnL2ekC/sV2aSyqxS/XkdjdNkbd8dhgg
KqEefMZaEbvI1b1O3t+yAkGwFfe40Kxpw9KA1ABGAPlhNr3ScsWmYpthb8HRs78J
1joTdYBRfKabFrnF6RpCv6X3CiJDDPNI9eNR0kfTqsNGLxI8cfECZezXQaVFrSb9
oGufH//hYIIvwwsAuQLfkF6W0SBx69yr6lpLTc5AAeMNWdwOLV3Q078nhSKxNvWL
jhvn6ypzhIhCamKcNGOxlUKr7YUsfDp/34TK7FZPncr1GpZ+VT0aphkhCVbaO17j
Y7TUXjdfPLCImTY7NDVgoJ3qyDVu4bOT7f3u0EBSZdnfj1LTU38jQEXzqXMGqxKj
jd+0CgTzURwdWrYo+UYH9rlMOsMC3N0au0CP5FG4hoBHkkgANTJ2OSBanRltXuyg
v6ZHfKSG/DA6UJpvYuZQoE2Y4kopzsglJtllD348plwte5I0nmIpXlWhVl9DurtL
aOM87EKqR06mhWHTU/KUiAjYFXpmzgrCCdWNc5mmXX4Nwb7dN8SGxQu9fNBQ5hqx
fd/0kfh9Uak5uwXLYg9DPvgIL4Z+Kw1ZNElspPy/1OvASR7LBW56yVqseGalaa2a
sWozZ5x8dovp+l7W5c8i+AiW+TUmYfUIvjsSb0r3ktfQoE8QCT1mwgiEcTbdQWHd
/XuxLwOTT3qeoRjrz3AMmb11WEegVu9jTH6T76mRawlfc0wMbmmvP9hSeH2m5Wov
2eZ9hdjpOwZ8m3EgzOMqGLukqEodJCkaKBLiubaQKXKdW2SdzOVOxMZuqfT+e8yz
EQC1mnUyD7O3DmCVotua7/SJA7JdL42bFCpMBCDWgIdOBTSOfG5aXhSyQYwQNQTP
52sviO4NlU8oi/K01yYZEN6l3H1tnwof5Db1HuuYHsx9gUQl8kZoOeCKGlosC+1Y
f+78n5CQJFBj4DIoi1qcjKdkURoQL6YOhSs58clDOtlAeQT+vRyelHeF+oGjzBqm
6weFVqHmWJolVUB8dghtG4OCyB7v6DVkyilmiwq+0NwZ+Kc3SQDgI/0YSHqZ3bwV
lkHSPqYXKzGo1FSLTtN8sF1KQ+NFRS+uAXTCx5pCZsccCyZRS0nB2vJjW+pCaYzD
ORXNSDJvB+NBfZHqxtf7PhzDl/cs0tExdh7pBG4zckcRB/42lyOl/RwZJXecxIkR
6oPIbSiOcTimXrrWyo7Z3Kw8fUUWrUa+Diqhq+ptBh5GfVwRGx1xq8z3/uWzBjiW
O3LkyB4gb8MpCk8d7kc4P2I4SSvQZ1+oYhRkvgrjUK1c/ntKIUarjc8Y4nLbbTaw
2kZLAoudPeHMi60/1j1HHp18sOnsV9v1HNf8vuSXc90nBjtqqCG/Nk4jc0qcLWsa
PSkcsccocfGg/tNyuP+BVeIjgekMNbCq/Ch42A8Ey+SnASeg+uQI/UiidEkaTbfA
Lhf1X1/hcW2vlHuqdUa6LSZdp7/+4NSi/gymWr/QhY0pgUuPEDecDgzDWUWiFw2J
lp42YoWi+eJhZxshLOkbvj0l9XXR7aKr+8OqynAHQh4sPxdhknMh/6sCWMoYnYH4
DsvWdC/qJoM1VGEaDsQy4VDxcpdH+oHxq82DQh0MSFYvXxfz2arV3A0tm764QN5B
625AeD4ziWwSse/2dGhA+tkYY4klBsd0gpSfoSQ6SDNGCA5dw1H8AuDQlGrOvivA
KgNID+asYxfY/OoI+x3sIAobpSqDRPtCiQ1HUlPzC21WQCSlQn5Q9FjPSPrRzo7e
5mjgOGmsMEmfL6bsoCtmNR6fIPciYssc/tkjyjH+CY5KsP60/ufWCri9ae4YtHxP
UsndxFX60IHRA3/Ujwm/Gh/Lwf60A2Nqtcw1oUsU4lA1kawebtwVy6atwQq2x6dD
1eeFx8qOXPSYgda6+v1i+OnP/G1QKGmP4JiSrukLMUhE50F+h+82T43JPnru45lB
aIiwjRBzDFsCMhTF5mYlwT4gezgOjoixdrZYVeAoS7cxrWp2LiC1PzbxU7NigT3Y
hijMsRF0KLKqdVGT4xt/RX14kPRlbS8cLzXSezwF+kqkNUlF45vJO1oZbScIrNux
goTeuGbTiOlCnfeSCzeJf5n0ZgJM3IcaHE2CRbVbNbAizf5WLZ4JjQs51OQ7eIdl
EHLNrRR50aTgpLbeIfwZ1T5QZEqntXQ5EklhIEO6Kg9tQNSwGqhzStRN2b3bsP6N
692e3IGwo1i1o442EsZzcUC4k453D5+ogR6y4JY6zfhVSntNC0a4MoMwsPfWQ55F
UJ6Jdqv+PbqOVZjjoQGJfLIG0q8dRXuDJ9c07WmJubO5nYbe+YbG4uRTbOCnfotQ
X9j62pjmxZcWNZcIHsyVqZw1Wn3p05uFLiNBbHoa7PoBRH3O8wWRIBKTGbe/A8VJ
FCEzkA8KgFW2rwYsCpL/sWhv1xWScCpFHOBrK2uPxvBPVZLSB1KcYzmDhJ57uDuB
HSStqKzYmqOJwev2ksJka5s1ob05iXf+1hnhwYm851hR7JlNkVJ4xpEFd7xcvcxM
nvsP6K8wMm0+R0YU+x3ygfI4WulxtPMiJ0NZKIifEG154HHZUYiuFs1mjlpluvkn
PU3C2v4dc9dnYZ2xhgggaAwxvWG1oY30bpz6yvZWsXWWKBdqLYMKRKiAMp2hcFBc
aa35q0PFcvj6aanR6ju0ggmNXdE4wrrvG3ngZvTDRQaJSGd6+MLtH07syLhCx68a
OAVmLxsBSkPBy36v+f4ixhq7zCj64Fici+CQVqKM4P+63pJ4rThE/x6bjVOsfxMU
2XBUaViM9H3+V9fGw+tpSGvKfZtJPoSltjXDW6n2UyqSHLjDHh/kFIuatTqi/Uga
Hdpfy5LfF7FrmMdj4QXzlRo4BxCdLRPHiaHSM61UKR8GwGVgdBxQJNlH8n4s6GEc
JOcpd4JGPDvn/MNj4VVWZkTs1i1kxv5W7zt23GEDMjB/TiEBfHOkiptkyfa4Mgwa
5Xl6Dz2McXdd1e3Bpz+SWnsmCp/mWmPxjFd63I+hKUqRj1v7giTgsF2p2nIZB77M
C19iNnHCFngNLtob0JCbMXdwEKNZXESeByBcLvQXD8BcrDAqjp3IYtQltQGMWKfx
QKL2gqgNWc2lpMkqHinQMOSrRhjcCKaMg2X1iuhT/cqTezI3DVmY0pyE8oCaTC1L
FRj5V8cQd3jXRmUK3nZWbkJwbeRI/YN71wsmnjSNLLQh5HU8o45cfrkzM4WwdtgI
3mCtHmIyPOXmZDi2cOpywKO+/oCYJ6Sjbim0Y3ZeeuzmwC7TSIPrgHqUsg9q0gJ/
WW+IHrS4VRPPzjRIzIMoGuK134OdacLDUjGNUEYxcjEb0D6N/4MYG5511hWW6tje
i9mRhhjoBb41TVCXXEyHem5b5I+chBE83vU41FJ1WXraK8ite1dWCDazfCDLiTIL
fAMFSCG1Q2KHE8g2z7mR0R30RTiEvP8ZZd7vDx9C374pm8qEfobcmPHbERORTRbK
AyBWhJ0WLsO2+I+07nh95w4O3XihgLTemc+ckAClygyKMALOAGRdhalae4cj6ucd
j3ek9vDXYwNkUnlrW/j2vKqMWTz0piUMdWVWEjDPthsc6jRpZjWH31KSMSW9Rqjy
KboiGGf2lXhltCQB4uYFZMDP93/jijnJVyeSHewDLB7AjwwXo6Mfg4p2Wk1pSaA3
YgAlseMQEq2knlk0LCphmR+OWxsyImTTS8AtHWBCKEsrg7ne43j7bXtrN5Mb4yJy
xN8OK4OEyN0tgv8zHpfLnLBAwo0U1V7e9rUQMrsrZOqbvlp4jMBB8DGJyMCFXwk6
A5fUXDfuwVhpjHYERcxU1RecY0ctEZ8CKIVtuuizPhbF6RJx5HHhNqNpMUqSyW/M
9RuGZnhgzosXNTAQueQt+6fqU+Ztn3HPiaVeOtzJlVq2Ks1Ij1Iy10bxbp4rTTca
4dg6nMRfMquSc5hejyqpRwVwVarBWuON+RnCQenaIwWYNhOTW/Xp9Il83P2pSxxg
mPmUcY1mZmo5wN8vZn+Z9olmR9dJUMSNVmYPdGYqvHPzjahMolR4qzC6NFbAocNh
/B3Dcn1FDhkZtVc7uEo1J44hMFIip1GxgBDU1j+GYqYTiyPmDo4tkmQoisY2f5Hg
FX23G2czXvk43SRMUTydbyP8vu7cim3z4+jU5aw0tBk8jFYr+kuQGk87ORgaBqEb
sNhoq2jrvZ3eHYr8VoAYpszmy5yEL4HTnSft25sdGcGa44xH6KNlS/GhlQtJ4UVV
whrFuXSmFhPXpR0XdjWdmaWle1a1cW5Q/CsKL31v7EDlRGwWQ8h2CpsoAC2Hogzt
aZSbkUCHaGhHIGT1Bm1ZBeTSYCRb6ZphTrC03HU8Kc0MG6URyzb0gDoKf976uDbp
89RyvwbScOwSKJ8xBV9lTEYsoYDPgkQW0zcTHdDHmlcGQMsugbacuas0zHFtIRDf
id0UssL04c8UAVCLyE7GMVsDFkSZZ53ZCaSV1HWv2dHB+xiQairkSam/smmu460Q
wsp/28o66N0//W/GPVSUHtZJnyt9sDfNMCET/x5L4jqyeWAQyAtzCKmRpGwudHuV
zr7JmFfph5FZC2v89KMTUrmtAI4jms31yKmLXdjK+yfo2wwB1h+1rnLSpXeHGsmK
9wbsodmgO4qN5Nm6qhljUdtdy3/ApELt9ABW1ahNE6CVT7rtyZeTGNvjS6ExdfeT
TXqfgMIWKEB0sLqW05GqGqejOe1HTGjAsi3lbsUd2W6+TvH2h7Rns65Smdc/c34W
+fqNxTUjeFD6mHoffLUGEMpCdlL5n/K/EqXvNPEY6Rg5bSFCsoytnX23QzcMTw1K
E2QiFuXtgMpRrFJDuLkXp5cO+7fTbbOM3f+hYSYl7iJ93aSqvKOS98k22kw+T1nv
/3izitxxBukQS9KXskHoOY79kcv61uVsDZ0o8MGNs5qLgqFQkmZMhvqdUj3aehAT
h72uNKtMmrcr0Tfvuh8EElz5ozdAptxaYXEZEb6bhVeV0eWdu9vZmOTVUm+w/aFY
UGsEfYDXAWALYie3dbFw4dCs7SFhb9YnrqNFsfJCC+nUclWbws8NLUNzBheqxCtb
VbwZ+MiUirvIm9dUn4vsR1dreJtGlEnEEYO6/kdOgCLTbo885T8kkQAryY1aIoRH
ethrQFN5zlkeRUCvQFW5ci743mDPRBUgBR5K9Bb2BgToYc1GET0L2sl9bBBRn0MT
bZEY3PafnTBBMJvcnjxssnR/jlMi0QWCLHlTWGZtPJ4yPFa95/cykmKoD//n043F
xEYEy99ocST9m2bgFx3Z3Lqx0MsBVotRKZBXJKZnDSyte+3FmA6WJiDkcAcc3/qa
BkaQQG1Xjq0cIBsFl7j7qzIEp/dpu6Aqi/2hli8qDoYvvg4yPyZRAVW5c6EkCLWp
btjSzRKKU9R5jLYpSeJVs4qhgTgaMTkpki3Np7dFvjurmAKaPbqErjJBVaGExtqB
BYUdpgbwjQnshyrCEcb4ih5M/9i6BXU4Wvy8iYWpprpjP6VpXqY5mtggRvG6Xijp
WdWN4jcec6tqEBfWeWWphepfQXbPf0mB3vnxthshj5+QldXtBd6RH74ivVhpBSUy
oZjR8fmiIfkXUDyS1NNL7kuk+ZTgWBH8aOejVO0Ws7WT8n80yHrF4gnIQedYecDx
DVpZtertFhm3vubfUmqCXhEKRnTOvlTBjk4A37grJzX5aTPTT/F3HipX3EPQUFrT
bKHpOKP3O4LKmu8xA27jNwU/0KbSJTyQmlUnDBRUKKqaCtwBzIfMJDu0P/5WtJHa
XouN0bzIWsDMz59HouBsqisjrmLMyiW4zjNgQpKH28knO7JrqTEiObEmkTH9TkV3
6/qUvNzksv10gLECv4Gd5m+OIAnzlLntgXd6niTT9d2k3QWJ4hytwO4zHJPaxdUA
9z18Qzwp7ROyAQI8JaC5uk512c1GJ9olWR9KKeOsXjfE+ZAsDSKsQRZSw55SFDMW
Bh07UQQ1YElrlF+OeHO5G1nxx3J8/TP2AdB6ksuSH8uuYCQaeuJ5LlOjyueUl/9G
9BmlDNrluaeXwMn+NY6Ik5FvMILtGvFm7mRLhPu+exDxNFHl2jC9Xqdzbs6I4ZJ4
0Avzf7TXzAv0B7XznTtgqKz2zAXORbLC57ghs7h61Oc1TkKwF9fGhgYRYhTP3nWb
smC2p9kIQvJCGizAYovUcbE0etRFu3jlWTnAhgE7BagfL7I9UA6+vbNXsZS6xxFW
M8JPAM7YTM6g20QcIRKPf2YxFaEx2/ZZtn4JiWd3YXsteySXNYRvKvieKTpUOap2
k8yu91YPPfcTErCYlIaS92YPYinuN44PqggguqQYIJ2kgwuVbJX6inCVQuG9eZQA
wcxcfxsC8vbwn/+oD8YegNotR2BYrp7YnMY/UMYBp/+wKHUPSg0o/SPdw1a7xghM
q2eZjdNR+8R0JXLjHi7aJKxpNuMVgetLams26XrKrGW9eWxT6o6AtlZeAbN2SO5A
PJrYETm/PGrBloAUllOX+2RsRyUgZ3RAyigVX3+Sg5Tpoj/NB50jHIgFDGGfUi0g
ND6yUi3NdwFHAyeG5IA1vatJHYf/nz/PvZhEGYrC+nfAe5z7WSW/FrhXyAS2Dcyu
rlDx+iGWsQvURIrmypOjfwwLlq/vFpsmcbRDhrpdTpPw7vLGtWRQ+NmxLdZcujj/
OY7HLG2oQnmE2SiVxiY1rzU98Ab8+81veQ2WacAspH5VpYmQ4A5+Z9suu1Szq74W
XnXsC4NtIAHowt5xusvEss8msGQEYoOuj1QNEnYpzArESaL9IQ13jMGBrfS2hMZM
+jMC7SQn1P0FeeaQySRxaYitxRLSnMAuOSs94P40viuc5qP4xxF2KcQDNcdkdqAD
n+IW3iH6HcWZmZtMzUDZHtWzu5A5lVjz9Zt4dtJB4DhZUmPGex51siuSuzIJV82j
zqE5vth8h4QtJtl482/KqscHlsT/Bk/MhPKIaE6vNrTLDZqz1u1pvyc5gUbvo2+/
YPcxx2a2JEstRr3pj6Cz3amXX0hot+KzWRmbvp8cN5z+ND+/KI/A/dKIU/EsGBYC
QaB9j70CE6C+vzLxPHiaTAVf4L1RxBXK2R3p3bRw7ksWN3ODeajIOoJk/5QTQ1N2
Cp8D70VPtkBBHqqduvWfVsQqiCTfLW89mxxwUANNULX367mzCq/1SyPIBMgnAljt
3GKqAFXsnIFYReRj1RRwmhO92dbVmrtZDBqY/dD/CGaTPsh9otgUIcJ5LlzMUh2a
VR4p3O5jVYym9tqvNLwHWky8DURYIPSEF1CTxlLSOzhH+pAMEvoKvJiCxgYHu6gv
XQTkyZulaQNMtdFpwGfx+v+mKB9lHgIhEG7gOKbz5pv4WoFgkkyoDiTFBy1S/B54
vrYizDb+hQ2vY8YQnaIETYbd3s4QArLLXooreZmZrRrLeGcMVK2G9peRmoqXc8yN
ciM+EaUvtJm4X8xwEdgBXnEN6GMK32TeSz0tZfMx7NPa5Ase93rkKrAXA0yVJwq/
to1v9c9bgAAAWPsXTvT7teO4GyNcHAVzoJmedVLFpF8Hxb+2U7IFuz0/fT/702/I
KZBOYyG/53uPJYPMsKp6Jp5iK/zYeIomQTLGr4SYl1wpCgaZ2mJrelzd2UTsgzQK
ERSVeGsN+xddVbdJMWdrwuGhMipTkdkA7QzD7DEXgHpUUv9G46QZKQDHIig6vSyw
SZc3VwkSGMpM3qjMM4ORXQ15eaVd+GNH/Np86BDYv4OPuax2DSUpXYagojg+5QZR
gPEPmYPVbQ0dZQNwHQ0MUIP5lBNH0z4/kVzNbzdGVpBBZ4iEXNRsVjO7rrPKMAYz
tG+Sg7505azNshp77nHlRHFQOGhzQIsC+VfGiFm4wZoyJpUsRAkbNkrv/exbqnTC
jgwYYFL88X5KIMtpr4h2vgTw1xYDmxK6K4SJS0PTazvRVIzf2gj9fY0qmjBWyCPV
F4ibOQTtrgbMiHb4XhOJD1B7ququ4NJP7rOiHLDwLykrtyOlEeSImbanXtnrwjrx
XT9wjjzvuzZAPCeriu/d9fXwQpMEKBRiEnkKerzI6F+fEj2l+M36QMby+yaWJCFx
Jz0jf/jSNYMgKJCO/ygryjCHhDPIYm5MKFNWNvNk0c+3zxf5Rru2XNk8Um/jAlEL
UB/eOL8NWHzCnzgaP6TfeiQFyjicsASO4PrrYSyk+BHYvlSKfmHFLHVGF2H0sv/U
v7HolQy+oQcohX82bOydx1SF5HKG/HeUPwLZuF2Hd4wOYgefb0OpJYvmuzZ96Uzu
TEA9X0llh18wjfdEuEsDT09blKWO3OO/DAHPR/AgRtMKN5eF5lteSg1o4zjP1j65
L1MfKzpJV/wsCluMiua+3S3kzK1vXpW++AVpNZazPNQEiF8mErn+o7pdaaiOfm5t
w1anSatFoSJISbNlBVBzeTdZhmlgyTIt2fRXXag7ZMULOUFAZDKjzIzu+e8NZnLB
QboOCfpBDWONrjG9P6HiloCmwRTKexNNzXJESj7lYKq9QuWE87UfGlnhaAj8M+pu
v19pqoU2O8TJ0QuEjJ6p2MqZpkXNuJDSQBm3lFUZcyUgSrhtc5I1GbpZwCXa9275
N1EJrqwXvyOyulsNm2du3A1LmVK3wjctnfAp3ODvafe/exLxUEPorT6bwXwei2oV
XC8PB/3ZJskCZ3EpTYk/rHo4A+6i4tXTOWvfZIHe64SMTkAwvoOF0E/fkj4nlzIh
bGLKepzxK8dJVOxbhM1NzlBvCeSmrhyLC1bGfIcmIkqsklHCwshHKm8BsQy7JYPZ
tD0Pd0734SEd1WN9ugOovozTjnm76yHkoHHpZw/twR1MFs748THzOLKm6cdX7iZ9
RupuqEH+VHYfLjM0gdhyk8fOifVVxoGlRrmTkyTYo+wev9NQ1YhSxv0uXUmi8mGe
iZVC2u+VvQyTJi+YhJd93ZHv2BnBql0cqmbSVIx68xagiptQ7dYEhmgy2Ms8zKwf
QAl3vrE0S4d1msMaU8ky++VPt2CO45fopuR36/oDLFKmTQpXM8nA0NA1EAdjRXwP
6+SagaY3Uo7cgny501TsdywAJIXs9RjJyg0HhtvSLRrE3aUgDI80GV+Q5j2gD7DG
2/5xv875Yi9g55HFl4ejgs1xnfKGu85lffU1Uqd7ACjsNDqfvWjRsEOchtEGotnk
mkiEUHmeUzwYclW9eexar1bApuu1fV3am+ArDh5YuRJwNxdTDUXrsFhAn1A/g+vc
3xMFK/V01vOQui6yq7YpPMB7Oqln3n3Yv/a0IothJ9W03+owiHXDXkWKG5aKqlfU
ITz9db/5sCBSCXIQS/sLsAgSPG/fUGOT4StbBUKGcSZHnQNnIqShKJmREjnQDcPv
+Qc1lv3QtKUteTuVGgvLpI2o2EO+HfKRW53YicmnqYTMuOCml+H4CFuSVZ2IKzhR
KmfHzXAelVyfMHmtHPhI/aDNiUeOGccNniWB9beLwikLhsmln4t1kWkGNwIqEOqF
8euCJpLFkyYicl6QduAJPzC+d7ApUpT0OpAkQpVF0qDVoM1ehIY1ETWZeL/qyKkw
Bzdowaeip/Z0w5wkMo+mpDW9oYOvUKnYLOooBy9JS1jnzcYRG8ZZLNFkOzPIptDy
fow6wAAvvMkcHNre7seK0c6jQuSUYtUEI8HbiAbAEEY9UPDmNZO64WbgkjFnlGdv
1RAn1Cdogyi0hNSXnaN8ivHlTxbkftAmhIqx8mFWm5qdwPdpdV2lXwj1BFl7HNHu
hiBan1No0dEnyYsMn5kZFekbuUgj3Dtav8C2KLZ9WVu65yUZnKfAG59fVm6fijj/
wGVc72fTSI3E1Rfn6Drnc6QMCYQBN6l9yyhnvFxV0MZ7liuhvBD3AweF7KQFHTAQ
xJoFnqz3kh9DxiqlsRZewxwG/DG5Sxxvi85vsz/jnWlEnyaONlODr5Hq+KjhMmcv
hjiA+cX5iamlSH9LPq3wqmbh44d0DGpyFFiKiZ1GhhXIRL2YK4Z3tEzXjKcU87NT
nU1JQRITVg0rEKhvn36rNXj9X51jonS0LBaiIHjw4p5Hzm2jOpcbH7ufE+oibKn7
BGVFo300B/FwK6k9y6Ge8goNX7FpHFPzLe+4JzoDJvVySX7XQPx+mjFpZlW60DjT
eg9/rckjf+ug3W/DtIVrTZq2cbSlu+7f1fD2cBtFxzQqG3d2A4Qv8fTI5cOQhOVK
ni2l53P/VERsZ01AUOrWl3DIrl4g+sotqibYBmUYMZ9p/T79L1k8czYKaUqWU7Kj

`pragma protect end_protected
