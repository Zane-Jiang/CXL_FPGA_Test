// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
0GHj6DlIX5Cw8u8dwiv2LK9sFGpGMG1sbEEPaLDKh1Xy1yWyqFlgzK8RbWkzQc7RRv4CfJEPb9Gl
Ni0QatpJA0hm9TEw5xxAjTK+XWWOph3MI/sfrZvLGLEbXasq8P91NpKEFbBCBZbByLZTuWFmrUAZ
vnfoE1Eo3n7VehL2Zrs43Obg/PwPGZhwOIfCgCMVCr564HX8SVPwoYLDSA+P0u9AL1khBSOy6LIK
1Pqec5cssTMqfDoA1N0lSfEKAFYN2pvYxGrIRw4O9+7MaCIgM7PFC3e9316iLkFnLUgOiEDDx7A9
NrzCik1hIhoz+b49k3lLAsC+2uy0/47IAebvMQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 30944)
VjFCoIhkiyc+yMxjuDArYnkkBdkllb3S5rhop2nZMSwSw+IcB8rvRo3emQNpA74cjjmvD/iRGoNE
ISM33ACZMs5qDbu7ZYuwgS5PsBnfEarkbXP13KA3ST19zzdAL9ZpqpJkxGaSwH86D73YbIN+VUIS
c8tEe9Zdtl8P7V07ciLX03JHDgEHXf9agjebLKEbbBxT6nZib7rerz77I23LlfwWx8w+nTsDXB/d
ufo3FNmY8Dx6M9Tn6zsHbkvCyWA46cORn0V+7a28TudB5FTvZ7QP6KAAqTzWPC0+++tV6NaGuKEY
7KgBrGJhvNG40JMgIskhtG6bulVSsoaPymHAFBP2QvU4LqQY5szIqXHGeNb+Qla2tA+1lT+iUsmV
zS/4o8IC2EuTPyfea8hXB0MXw/Ft4yQMnq2MWTlf8NBWmVYG6Tl++HII5zMZY6Unghkm8jNOQLah
c8rmd5zvN+yVUQAsJHqMwMDEQ86LcOAQdGBZj0HxhGzgsXj1V74zJyDdWg+9vheOGahVJCyxaQkW
ATvirOUEPI1YzAEB95RC5JdexLDRBvk0HRYKCpHMbgi1BbjUtrouJ1gVIiibTYLPJLOdRGT2ahsh
WIynSRSXXSaRiEI2/GOfDgrUWRmTsJPYao6pPRb2GvTz2M5iXh5ZQu6ol/gllUzA74bWabrvzLJF
k95lSSLCglsf4jM8WpHf51xjN7mOLa03fLh1l0f1pxMjfp4Xm5RC8wYI5sMzp3HGIu7cPaEpZzOo
WspGC7byXL2i0YkKZ91QH+aNG0DQYl1ikZiiOxOjfJRn2gCZvxkmoN5EuT1PA+wNgRwOCYIH4RpV
yINL1tjZBWK75ypD7BTzILS+vy/6Pu+XQs823BhdMSwfqoA/uwU6Xkx32rTfzUINEO7y+9hcEDI3
WdaFGWMusoDVoO9//UmJ2L/mZGGZGC4XpGWsYIF7lRxF37iSOCqfF1qh+FAMgnchJ61iYwZoue4j
C9H/7KqYF/xfAWcJwiCuLyUo+JhgzhDkr9r8mD3DpWwmJItn1/ay4w1ZnHKR7L/0l9D1hGDHyP4T
F2GF+rOjBE2+JVZ9qEAwVUJ0JIPf/bbSOiitDYAhhRST6NHPtykIS1bvf5JMHNWOb9HuukK0NB85
VfQpR5Z3ggv3rEgGf+VCIa4wP2T52ibFAvg+bs16z/owThxUF1gHWQlFF7nTCtoTXXUFpANHmHV4
IQO767aFJk9/GtpBVUixKc+4l5LyXQB1iBYyTUEGh+HhZDBK1aKmYLXd/bz3pzYRvbSkPRqXtLxx
BOF20BOhhqjvs2EpNneYCRN7GKT7uSZIGce4Ql1+/zqrQnA+MR8QHMkKBi7llniiXz3TUa1jht+Y
lg8CDwa7Qig6PFUkukm1QXRv1B+o4y9Y6LIRV6GbpFCRWMM+PcSX0tLuJe0+MfFqIoBX3Od9Yoni
rjbzJMX+jhvC1SjwfcDZVAGaqvnoOXSsmF27p6St41RyovsPs7aAg9irRJgv96MD0nF/P2S1I8bU
uLGyA4c66I1RSmK2N9qNsXkUfRX0B21HIW/SAisyk/DbjfodnaE+n2tOLAEYFdV1VqwGSM9GJpIN
50lN20BhoL502yB7+/lORGuw5gKjOWbKIoQ8jgeXoanzR0oKTvLoHhPpC90HXCfv6Olus6a5+XMG
5JQGgE+CRWd3DTgHk4Ii1C1mQGGFHTzxRFoxev3daj2JMCKpUszAY+kIk/dSF1Pg3m9oszIr2lWY
qdkXEBKvjD82ZW+VNaKNnX/4stUZwsSFLSr6eUpPsJ3NnBajmI69eIhsK397zB1lfMABxdM8jHI5
VZg+gTJczjnjvE5BgCGM9wJOIpf6gmqzAOgMfrHTZk8U+S8IvAae+klhf/MUnY4UFHYC28z4DQBF
cIkyVClDY9ZgXr/ymye24vdtt68lla/ummqG321+Fgrcfe1gYUOn01zMbUMTp13hZ09/1BGlGguZ
81FN5pTaWqTQkCHdjbQuOLLAwAilb9xnLJsP6ykpGX/gJurncHlDISI4f0lBYYn7WESY852FRotI
w1CKhfMjJqy7kpGQq2HtwbzW3dgYvSXHPaIlQJQEzO+J02/XETFPEe9Vv7hFQGRDrgtJCvuqf5Wo
S0QcbiNutB9aSNF2c9Z7dQhECVGGu+B5bVVwMDSeqe1FawOHPwTeiYyEzAoTq5B8ntu8Dx19VnQK
QXP2R3O308Y1ZlhOA6/7zN1gjk7PSRt1jOM166kfL9liAt79006PCbNuGTOySXSM68ME7nNjf4Pf
+v1l4hy66WQCmAvEiiI24z65ycWP86IF4QPFY+y1fWl2PF4WOcBikZiOq1bxAkGSga+zvRZtLkKv
uFw9YAUAkD7b1A76cR7173DtakcAW7UKxx9YSIYiSWnmmef4HarLERYfuFbXW82tCoWv+Eu5mXw1
LS9XTY6zkjmkkzXBtJTxPXF+hcW8595pkC5nuMbGGksVcA1lIuNZadw0JMoX1/4/t+1PIpVOJGd0
9hsnAVc20YxIZVnw5NIkDdvEJNr5pNpMkm3SjeXtdJ/q9WhdWq4rwq0Ce8N5kTEZiD+3WolD0G6R
KAW8FdCGTKKYEqWHvFNCi6GjEGtS5o2fY4kX2JyyHMtcdHCkd4kKsuhtRujycRQM7qabLZhQhT6+
BfXtuv9UQoiseG4I4WRDJUWQUALTNVGSWaE5KjfajoZixXZBeKORAdVwl8GI3Kr4oNKzMz4GrtMr
A67L/PgG4Ldl5Po93rHKwdZeCMosx3tzskSneuxuymowpDH7J0ACp6BwwAl41VYU4AEh9Vj3+/JC
cqCEcwzltyq94oEQYEYgh1RWIt/Dn9iwiaBfNBvaC4ntDDIzOTucvshNec175Zfhqb7+34odN8Ef
8k8Q4BgWFABz6teRR9AzJSXXVPygq5Nbvbnjf9+hWERdaa7D5zzgi60d2PYnFQq4y4WbbqRZmfz7
x4hxoGx7uy4wpE7uA4B06mSU9R3wq97YRZteZu2hHTam2e8g7E7fJkh5TuK+b/Xb5qbJ5GIfJTZs
7LioN6Qh18ZOKhHL+oeqh/ScLpRlnaa1LwhIy8v/MZ/GESk4YgVjOK1hrgAy5dnSzn2dBd7aH31k
H+0uS4tCws33XVfqRT6dAW4CC0y39NOBCdkEcgwp9VGuzYG9dMAeM8n61O7eziAYATmK/veEOmBx
jlvq6YCoQxwvUU37SCpQo9GHLKitCuQRf6htGOi7rvHyt3brB1cymfzJJOVZG3qfbmSTMl/w81QK
LZI8jbn7Y1d1H6w1CgnTgqKsas4j5lx0H78jpIg9hOmBu9UNUDljxMdZwhj+roSUhKGGzWkmrFe4
/wIsfMziEbdj31QHwbGxzfcHbR7R1CJduj8u2klGMAw9WmDMP1ESEnsECfiqRQnDzwTvObc4pDhr
9O4/uSTBnIthutGGevibo0loDxI5RhuT5urebZcvoozQF4BnBrbRxPD26gvRo5gBrfkXs60ftLJG
33CJ8+xhxePhBpRVkacIPwC9MJnPU7MY6hg4ZKITCntdRdlb1Aw9CkoLCbA1I+BGTjPRn8JW5zlA
MrcFQbsHih/2f5XBClvth+vM8/nysXbqW//ZoYG9t11HjA+qlWhV/b3f8Or/riG7MuBu3n4vOenG
42Kp/ZHiiZOGL3bcX/sMIDrBFxKuQnETKrlniamT+Yb2GyNazsDeJhkOrBmPNKJFV5Aa4PU97Pp+
PnZFpOWeJQo4vG5zpMNDAS/uLt1VM284vErgcj+lXDAlK9JS9ngfi/ZDH3Z5LHnIMfMDx+RZ4n5s
KaS2SBv78Ws7QMALtIR9EHlI6LJO4Agz95j9/sDF6hS0rBWXLokYjZbV9hvJaZ4fO6pp6bPySZIY
2QKp5DPXe81d5c9JjyAeDWYZMF6zsUjrntlO9+ZdH2gut8bYrfChkDS5RT8V20yHIqw/4OYWAk6f
1LZKjzSm5mBlGPw1iNSf6FLNHV5G0ox4mUfC96Kg4SrjMUFp+0IzyVOS9mXs4aG8OKkc4avbzv70
QQ6UZ8BT04LvvqCysMpbrW9U8RIAK22nEhPUADLDmef4iTYwf7GF50MzM+yL8cld0JLuvGuUYetH
rWs0IQPRywtMtljuwMfCwCffvd/+c65yxjiLNB6TVd4cd1oZJVZEM2IwxEp5zHNX9eaCK1z8BXYH
GriaKAmYX1A0v12PJHR1RSwLMkpSM9Ac+kL6zps6vEFSFLlOqnUYAZdJn16VxxgV0ia7vTP/3rq9
pB+oI5ok4F7XvX7oeXVdLkWOxStmNNazod0efYqx34KeU8Mu5n1ddODuQZULsUOPZlYgUcrf1WMV
cpvzG5Z2tvA+MMNyFxgqmz0Zsdlg5xA+ieM6zoDglvoRtcow4NYUm0lNFKWphtc9uZZ6rSD5ueOm
wk7n/gyOosHn9niU6+I+B3liGYKaZQDJ3jE4I9FTRH7/M+s1jOFWngVu2sHWpNciusZWq2hsk0jX
B2LTouqVYD1siZB+VPhk1e8+8rJ/HPilS/4qkS9JST3JStPfGFmeyX8WZeNPPoVwrdqZWL5bKYMV
uTbH/fbMulvcybHeacQNTUOBkIQ1/kfBsVKPAcABOWDTMTN4zH2BsqkBevuZViykRbZxyH8rfo1U
47s8CinGUvfgEYsHv+QyKSD02pgNiIOkxazddh4ZV2uHxhE0n0RRddRgNhFf6QHzqU89MUjDV1SB
4mx+1BP6Qz4my6Y92y9BSl3Jj24PcJJsFnekQNWEB613Txts7gZE6Y9oZ5f18KcBR1uC6j/yKFKr
ox473jVjGogZg4JLLrGdIhb9HLufgJO51339jacwCuKpOmIg7uf1M5/oTK8y5hm86QmjNRnyyIU6
moZ9V2e7qweMfddZYAz1oK89SycEfPV3zYcSSpgLdvQqg/wKh5ScnWR8/5XYQ199XC7NH5FB8qe0
Cb5+lM1PosMhGlI/dPi3wOfkiMVFsPDQdQ/ZF52NH+xkwGEK6hh5rQS4GIfg0TqpqLh3flBxY1xq
iSxr0eQE/RrZo+pHpgIDuC75bXcxlzN1ckJq5fe5SDV/o0/aVeluk/EGibddJZ54OlVN4ckCLRsF
xb8+jXS8laI7y3E7QKBSQbQHJrFl2ZhjJAyBXwjP0ai0vfcWN7FYZwRDoe2bGIS1+avKlhYIz+QF
0R4ZAiBKGcOYAkJEBqRr9c3R7B/Z3owdyqyePB1IZHGcai0d9FH9OK4MEPCSiqGSN0lixUP702NL
gfN4oszN8MTb4P0biIkSJTybm8xTny8Ma0vGLTXxm32Xb9XZnmw36FAF+qyDe7EyUCJ1ksKL++kZ
TiIAUUNlfGYiD3YymyYRw3Ce7Us5T8VjjYSXOz31Y0es0yOAx/qgGytt87ZDsKI/33IOBSI9QRqI
Rwi5qa1ALiYU0QLrBRQ35O1Llzj2jkI62Tq1DFt7+j/k853f6PKEyaMhZ965yQRDm/+d/JaIDB1N
DPtDRoReNOqP3OdiZBv8UQL095aJO1ztY0eFR4ynx2hYnjRkx8b32m2QW/Nq2FYMQjnHCpS5yGxA
wWVtcsYQ92TYh6oFTZUhLzThrcgRhrVODeFBpLSgGifcvIVGh3T5sR2le58sJ9jU6jm3+zfQjJsJ
9FLJs65zanQ9VXWezTG2E4MEiCMlVngwtkWuU+pUjU9X5nLorXcOlC73t8N/kxvky88SOLAQpD10
Se4POAZgOhIvEb2A/KC/bqhPSlgY6NervsYvjMkRbetbs5nNTDXOn/bVUZm90JAMJ77LjQY2Wadi
dDR0h26yQvI5CUtYl70hUNcpZSo104VlwSDZA7pvJwEHPwHj8kxhG+kywJGaEOc89Bjt/RUTfKrZ
AO/DdzDGC3LvWaCTvebsH4mkB3SOt22oAmPV+l2DHyl5//6VS0Vrs9AoFAzmZRZXvOVA3iAek4Kp
4mDX7DTNY0658K+kzk52vM2Dim3VGA6hwZinrLZhKtF7z4RwD2b2mPmmmXeBXHALz4yNIdUyAAUK
c5OpypziWlY9p+Rfnufq9hWmkKddHfD2yPItnoAu6qqzbKlsGF6BXzjHXfwx6qjKin7+dAoSjVTG
o116NAM+gLyduyEPVM9I9eeFxuvPiYrfrpas0npWoH/fJFC2c1XKx9wKeEVMDlDk8FGyHeV6ycsQ
HGqEb6PdPyV1Ygv5zWtqgaZfGVUay3ayw+LAbHXy7e85iMYDFqQUfd1WnDTm3d7QJ89Oku9SLWZH
ItkhKfGRYYC/cejhfHrFGOhAauo8DH+33DSeF6H3g7HrThHCjd4pVFo3wCAjU9/GoxjyDosFWw3a
hFtxVANuFm0tMkSDaEzZf85bfKN/g+mBwFivatXBJ3OLZzbe13rGq4g9vT3GrpBl5IRX9ihyRffw
Kog4cGE1NOeEwGjbNZdA/CNoFZaIDRhJXpI16Kg9bRcmd6TZy6q3XmfjWTLfbfGfjIhXOPS6wrD6
ZCFW1l0UKG0d/PbC2rnBl4MEzL9rX/Hm8KN/bC152pniTkHXHk0A+WW3LLXNsAk5p8YP9W75klw2
HbaLfsQaAQ0qvtwuj1QGRROL6lpXr1aWnzHAvNbkKtki70Xo7+fbXTCuiCbOa5tNwbc1RYleW1Nn
HJ2iexJQjJQG/bJPAz6Yfyv2cwO+sAzho6ec9AvYkRe4MbU1uq6EelN5r+oBryuHGnEGHp90eOFS
WL/fL1FNxyVVmZfoYLYGagFoTxT1frVjrCUaau634P6KEKJb2X1UUy13PTpEuYspGMXjtPEgFWf4
WJ09xJuTdsHGmCqhpttl6Alw06YSYgLukf3uWsIvf7yLxkOypJ0qfx0KysoJKoSgLCtktMRsPaCU
tpLGDUh9/GXiSSXcva4MjctFI7ctZN7cX5FDCMNczoHXJP35tgKO1yuVCrnr8pFI06L/k7YB1G1d
LQazD42oBS3qFNbKIn44A8+zbXbW9RdGIbBehzq3mhcZIEi42kndvtt2aVc5jw6QQJTBynLWZ96h
rpu1wwWalSmhNIRBMQ6sfCmWsEQWcOCPJgU5f06fm0jjzpADSutQeFpvAI973BYELUH7LONl2KkK
Q3jRlXIHnwLDKThfB67JV9d0KOyFlMZx9AI/lMgQZ65THvvRC/RhAvjgR2YQm6x0RGq0cXJOttw8
aM+zJeFWjMk1ip/NJnhhirGQWW/COThIf5iO4Dkd6w2/eTuKfSn5jNYsHGwuja4k9cm5xTGPkjR4
3NQUtzryyB8WDd3kTeMJwYlWzoJl+IlXrhcgawC8HKbZff1ZcxDrtLxCmag0stawtonT0ZaUxtlm
lxxGZ8RCsKP6eja9Ru1Ms6GuYjxcmABmEbBmTA3W5rMFTb7T9Tegn0oXNfzheRa7Z4V3OpLyVBdT
uBFXyvVDX3zRxCcjOnVmaekOEW2Fft6KvSfhV+BQurWB2HUCJyiZT8HiB/ECKSMFVfA+/yruhMeh
BrBUuPiewGYnRSBxstKoY+GlDeI0f/msUSZ+yqPgC6UwKO450uEBQ2nUHLUFrbwH5twS4BKfyIlK
Cg3cpsJbGNRAaYBjQlC51r1Z53BRvhz2LfLWCpezIVHFNi6LCfdY7NSZH4VUwJFNl+mC8Ak9Gcbs
IJBG7Ju4KP8SbkRILH0/C/etp0k3fumLcU4/bg9JQ7Vrkil7OXngSI8f6OyxbmUNbJ88cMxUxuLw
kOzpc5S57msWVcZqi0yXFB/9D8jUggMblR9haxJR1shWY9iXQefifBhwgS9lZyfkkS0f1UbiPbMM
8CaACRAvFBG9qakhMateg8jkbEFOLcQeTb7ANfi7tD9y/yNODiwThXimmIHKgpHO9FFks41jsr9+
bvYV6ayEBcvC1BJX9mF+jI+WJxLU4GRNXcQwaVi4PWzmFXJnAjEdggQTINv3r+j+Tl9NWGh6wUO5
z5W/39LNxvo6qAeGH9hFE3JZsBuy3Iv2d0x1rL5bUmzsqblB6bcEGJGowDa/bHaw6IQvIeQp/elh
hB3nX+xvNa/S5yzkcBU5wFB6GT1s+zjK/74+AVW+rWvO+sI3PW0B8gyyhxiicim/uNdAeABBO2uH
XMC4i+IVhqGhqXXR830JAM4pTLxWyoN63xPI7aUVOY0o+YkaZH7GDQaWsHY902fypDU2tLmDk4cm
dHF+i9wq8V4268LTzlOgxuJwCVEQpFnUNKxj+bM0E7yAKrui+QEh8HVGIdJtUoy688ImS85O8r/O
FoxaBUAztHdLtSqn1oaZ+HJtz7SJKWF9LUL+64voIqk43HbfXZBSC4R17uzl0y/s5htoCPZe45Gb
WIOXjieIwhCEGQfOZM5VDh4UIdVjFZ+zhETfHNzLD94cUfRRv6e01S4RUuEGxiRXQonJFt9adwHj
TeuSaDz9obcn7mP14gTLXSk/xf0/aLEZN1zeQ8BQBnLf0rNGoYde5ad0t6j7ae7Y9AFh+iuHFjdf
nvrFkBSfhPrTWw0hHF1fQBpgHP6YVOM2FwGivcJHASO3mLt3TRJ/OXBSLh3BBeYtwUbewDbQAuHR
4EhPzDGiIKM49j0Qne/RcrTKayWBimDNB7IQyU3zvWRYvZRB4ETOSYxqH0XAo1kz1rIlHa3Hw6jp
8RHHKlRVBJ/KmLxdjuJkdLGWVDscx9qaOsGtiveyFeyGdSf0g7uMPAxThidr2Rf23tWSSkuDpvSs
7zTelAHvlPl/JVgtGWy0ib5RjKBMgEb9he7axwo5J8pMjQxopmCPn8G1l4aCvBAirJ4inZ+GsiT3
q7kSVoS8yJGMNoM19ROmlQKJzdyKKq8OMaVyivhGat1Ghlv5YtzjnEtWlJG3/s5virR/GiRpym5C
zrwC6J08Ro5Cj5/C+DtMJ97umGPcWbPL4fbkwhS6+u5WEuMJ6XqvIYysiwdlg2BX0+BYzwexx5Bi
Llqz9sCs5v3attJngIKMAGQf884XkhmQZrvkORG1GwaFovJ6YV5G7Je2tP0sJbBhUkjm7rmlpM3g
+IXT1dWm8C5MLchyoOjJEJgzPKm+IFQl/jSJx4GwFpc2bTL4Rb4k27jTvDJtrAuEGaAV7ut41KOv
tJCidp7qWAL+tmINZSIKmUSJSm4RQZgJJ+WuKBIgml94CVsnsnnILI7kTlb3ndomgAghKxzG+82r
pRyTt7n0DmC0UUEZO6vtXZtNVwnarNsJXaHAJu35B0AuUZYui3NBIXuT30WmtzdjqKXXYD5pl12t
j8t4BYfAUskxtweLb4yCY/lTIbdxqOb2vrEyhEQ6EC+U97IhBMJh8f73SY0AHmxj8eCYfAS0ir6Y
05Ydh0F42qVb10qTuO2352htlMf9Pek4oe+p/aVSLksyOnSyo0D8MrKbroqm6OC5wF1urIynAS9E
7m0G0u4CEZ+Iys/W7LR1oh6dOGNpb7kHXqyRo2/o/Ei5446ABGv2/jxYohyHkuJ/HV9enFx994/N
0XmdxqzlkyNDehAg/nrvuxBPlwlhLdEOy6BH0khaZbebL+SgqrDT7IN6ywszymClGQYOdfZoHAav
TH0bZ115zxOhoJdKHlqrH2AF44kma9J0uZdFLc4RqxMGSA/1/xEZUYEB2J+w1oP3fMIs/NCpLR42
OgO5l1Y+H2fbnTCWvKUtUcqsj/5MtDFm1cno14jtB4C8wdG++dxYwhKSz1sFdTHmlJ7efN35DWnC
GCZuAh4j6HeV6ypPyJQwiLy7WzhtD3d0+X6szhQt8xwsnD4RmFCZzt4sjMSNtWaIu1WDKpJfUi1F
WeyCf88BKJTdZ8lVa12N8sH4WAtFNo2Mo3PgHyTDyq9rbkvN9kfdTyvli4ZJTMbAb99DIfwYm7LT
AjAnJGXuddcKGaEix89t0w2wSzRAaU5vF9N9tpNNVaWGVIHnZ1wOtD0Cvp7hl8SUvHnf5tzqtYsb
cPaQr9BSj19XxllKsmRG+e7GQTc6oGvkFiQkVjHbUa/Sw+XMC9GFZ+0hQOciK+pw+oRNqUNoh5+z
CZ0tfBIrq6+VAe+u91SvF8e4W5p3i7C7dPK8PtRbk50dOH+FQnFUaG1BGk4egzgae0SPMnXz78lb
RwLEnDTYQNb8z/wrSquumaaPGC59M9Wi170G5iv+pxg8CItNbYhxLMghz9UhKfWCw9EnTbQKvN0V
Z5oIgucalKtxuo9DCLTyT+uUep2rmxjGXgjcrypaL3hApUtokd49sjNBohQpjMzp13CldNFymjuu
MjPJ1eWHN3H8j/VKLWLqYqwfYL+IdCUZUSYU0snU0Zs57SyuGcJQ5szml/jeHVaisJnWW7I+mI5E
rq0L9jXAwEuVmUPdnGWO1CDLqalcLiEnyO8D7l6oYmq4fw1lqhe4Ybi9oMgTZyz4lczVt8zQUqrR
siO+fJuDznAizwJ6t1wO+hu7Q/jNaZr2ShlhQA1kFyZO46n3CuzfG7lbVVS8G/gT1BGmX+rLArdm
1SffMS4N7VS+wZuxPkBswKMzzU8tQ4Lr1CHkrT/MoqKGZlhqTw5eCzQlhO0T+2etxc/SqZbqySBU
ZjQxAk3BiDQ5CBhPH6O8ncssbzpndLFFmp7x2gop74AAjNSSfzAKPUA4XLKaSSGR0PpYZt9K/NQi
jyVr5HdEkGVcYXjFSX5szkRnd+oxV4uNNX9+yzN2vx6yvPDTr2nPNxbAI1NLURwPf7GHzoPnEdx8
Vj2dOETJYmjRNS3y3v+goNfl5QMWtW9KuvhU2R3TVUzpwZs83UrmQIfYIzgnd819Eu/x4yHnKCnW
zJ5MUqyI4syVRvA4eNomCV3/a9Fgc9E5Ky1Yp5AAAE9dTG9EmjO3Ebpsyqvjg9o6KKAqQk5GqQBX
HediqpouuniBJwYraTqI9CbaRDPLyMrHkMweLCgecleMYE2iPtyRtyVom407mdhW6hVhRr5AUDuH
fj6/7FXUgzoJdzCGBEqAW0oidnxDqUVDbn/+oRoA7QnMwIhj6WGuO67nd2hCYIYf+inm3/f1AIW1
N70Oj+QQLUPjDZACovx5GSKvXukgGVfZe2Q6F8jBKIIxf8EtX0bAmjngy7MDbBRnVMdDw5lunRh7
ujkodrnQyHIN/nC0qWKLx/aRFJbqkc2TcWuN6iq6OTLHnNjdxYfN4CEV0JNeG7vOsp8r1I5Gndnr
JNSkkf0+n54wEJqL5pwdHTaW5IXO+3geUNY5sHZly12lPEM2V5TX0lrXZO1aKwFGREnlNkh5oj6y
KonqamVn7fklPoXspJ6IoiRx2A9R4bnmWsyEVskUEO6IYPzRqwT9oHv4jw5QLhcOeKAMN+LH6Z61
B0OjY8QYB4WBLE8o6jDBUEpg6s8OEcRmJP/xj+RAtVeIpjGdcniy6aifghxJPJ/+aE/jgFkUGDUY
wGpqdC7VXi1LvGjy8Eg2ohj1bYjCUm7q6UF2OBJFD4pVWmwkAlyhCAZfeRcwDcKPOT/2T8WrYFHN
cTq8F2dnRqkz4dNi2BOcZ5DwcNfe7bPtx75X91P38XTmWwayVISDLza6KVYYcLO1jPl7PkBkUUXm
mM9AXe/ZsXdCp1If6xg2tqo2mbueuROu+TeGxUB7Mxwv5Gkc1SMNLbKkUtFOYHef1GGTXk3mTaM6
vSzZa8oCkOrR1kH18De9O5Dx2n9Uz8FQugptSinDwlvdN1OG6FfFhsBgVd/LlchUltmXCI33aTsU
BIkXgTctqM0NyDpKHtGYF+U3bcK5PS8KQRAxe6VmKRF/5T6LKZEkMTXVQyWvz5rcidN7Dk0Q4vzB
2v0slqEy+aOGFLthwkHt9IS4IDyntIfl0LiTROquBdXjFvwcfMrf0SHn3rgzmPip7e5T23alVUCA
cocgdXwFLq0J9sCx7fHoti4DaGzzN1JADpcHSCwBM/uSMb9DC1AILok1TvPN69wtPybUFNGWjVH4
wi4EDeQNyjzLzdTHy2F3qreyy9svpeC6kXZkyTexLXg34T5jSS6YljXkKT9D1W9OxYpOXNfzgGVC
gGlMMVQLakFmDoXipF2/gW+q9YvEq4EIvRRGaSAGjlQGbDU16Cz/r1UbwD9yUVmyI1sUjs5lkws/
5odBhs+UCfhuZjr4xOjxxV8hJGlg+m3D6AgXkv4TSP3JbrijK7TeA60BNsVJ2dginvT9KRyqEzrS
qjledmzzjUSZamRPusxe82f/0N490H6PJBEdTlg3/VmLF4VkslsJtT+BXiCZUGuPgIVi7J9fxQjb
z3nIm8YyJvNJdWbw3jsIk5+5oaR0oYzuud2VuWx8OS7PaVhjWNnmpT6SzcBhk/VgGuIBZ2ooLn9d
WT1+qQgrRyJfzHa0TtQ//LkwxB2WCN3OEbd6pMorc+H4S31QkgUyJDD1gz6WKiBX7GvKTCyfm+gC
2EJHrOO3vXiuCs4dG8jSx/XYr/R+YL4Jr8C83t9CwNZaoJgi4IFgnagtZp8slqe+jGUvlhX6vBlW
sZ3e8EyQUzTXr/VCdFVUTILAAUdFY0DRhSCe9tcZb9+/XpEQl67Zx31Oz1+7LobZn7ep7cPQ3PFw
/QZiSEIIkZ8TABf1qMyROWwUwcxX9iGeIJLETYJbIS5Kjo3fCieqMhcNg9gGqGXtFZNvDRwp5s0B
5PK+bHzh3TjSKZ789w3rIxcGu/HF8np1fbHAZWbhR4rJzaaHSSLEziucg/hOT+4yMdSP0VHRQ4/u
YMSAmI3r8HRlkvOHSi+VCxMjnZqhKOKChtsd9YKHUxp/Sfz+q8JAvEC/RNaXLS9pIarJhzG+hR6H
y5mK22foXoPviPprAyEyTlNlIy0QZh36zOEkMO5kzSrb1ZinGwE20fhO99UfBYHj3U0Yavy/AdT0
Ss175xQD9QbYsZLUuBUByIp6cCYh4wMrwlaZcb0skgOry+WQPIotNYvYxAzMK3r+4Ky73tUcwDnG
uokP5jWUOobsN44NS00KjGQqvgTAEMiY81jTumYFe4Jt7L/NVlbTrjDexPevOlv0+ceyry4dvl+v
4wqrn2oqrSh9QT4DoKGdC8JwKfPBJpdSu06Re9Leb2Ca9FWJy6cP4/W7WbJ3MjjCxm1UavWKRNST
qd5dk6j2V++Zz9TzjpAcrJqO72c2Cn6VJjYpRvDfjEdVH0ciuTqo90v4sabjnEEZdKKVvk+Zkbno
iYZLSldBmS8F7Skm0K9erl7fuBWu8gLWblNWwV5TBYm42yxSW0ZaEjtZl9W1a+1DUWIdMjJRK2T5
boI46d71AXljC7gvvsRnbyA9GLtN67AqFE/1Z+/9zWhf9cbphwAJS8GmjvgU0HX0DtzEXTnJOmI3
4fEhB0YXgko2MZgPgzyWEc22EB7eFNdpvw4yImST8JOw/0PWDeF/eYp5n5LZ9XA3a8pmO7wtlw3y
F9YGwCN/kr7vcUYnQ0jaWnOOUqEqrqkHSjf94tQf4pSsfx7IoZQR7Pb3JvrboNZHQy+YiLhUyimm
ABubRwB3ZFYUk8/CQhPeq5D8VJ0SU/gc9KnOzN0FTlgRihUTMAmUb7EpjV0m/+tuMXKaWYrfghgN
tNg/s7yTuhUGg0jAbmcgpvJmC7kNXB+JpPRfGzLzPBpl2/zgednZ8+sZVMJ2ZAIaWV3OQEPlLHSJ
ibbFsw5JjU0QH7/inRFyGfZeshY68XEOsxzWuffu2fbUjQI0Ur6Wj893ej8joBAXLcrt7kHJXl5b
8fvW1laje1kiDM7wmL1EfOJU2ZvBsGAOiq/sdFYEg1k/XsSRtgkOiu73OW/Jg62XaNBausjznuyw
VM9P5CT+ig9J+uyVVAdgEwcPx4EhMBG3FA/dVoYRuATGicQuE8zbhjCCvujzIYPuejqONsFZ+Fgv
bZOj9xS1zw8vwZDxKKvq61wuMJu9LBhZ0sACTbg7YgzDvxoSAm/uqKDMyNC48QA6zydQ7geMPWrl
nKt2GKMe3b6YYLYIP8oGFIRBVawOe8hNW/CfHE5me1Pw5JP55KcrLgOA4/X6vNx4G4WOYU74gzoE
xbro2BsBhzyC2qFFtWgeFxOjriAy3Aw6h4VhHFTw+Kf4wDVNSHyZpvXz7+1Dc8lHWFIWe56gbrbv
bgThcroj1YxKywWxD4qAkBBEZr0w3n+2kZucZ2lQkuy5NBoHfMQIx1XFqMXj/zXCSuQkPeAJCHHs
TyWwLmRNPRnObCyBAvwzDpiV5bASzcJReiyK9NQ+b1+nRoFy27eulNN9dI7yxojxMzRk/8VJZ2lX
ASmBJIcGyM4QtyXadpkNja8VNuQhEmo6AHcuTiQlOi7NTXDNkb0wCMF7R9NgpsXF+DY4C8/n1VFq
cTZIa/hM/kcgeqlt+8f4jysirIOSv769PkvQB7trIBxlHIe1UnIB6V5dX7f+eOX2daWm83Z3NxAN
iRO0VInGCK2GLF37Rl/14JpNRrcAECPn4LeDpzPcN3tSG9I1LtPY6tQ8+Am6wzhejmx9zZzYpUvJ
8A78PQ320uUir2dI9I3f4vM/IBFqkjupVBlNqQ27MFeRBqJGQDOqOP+OiVCJAVkRV9B2G/c+F1iN
rIkBifPeSi6ZIawvhjhkP9zCp1wAJnmA6jmdM/u5bnGyGo5oPUUb8tW8LgQNC4BjoASVvM7hiuFL
Go3y8LQEOWOu2rJwnu455gRdjb9YPMEVpjDXnb4mb4dxIclXFexbVdsg1kfgs6JK1qX1536jQHpQ
bNwXJ63GHAtS4R7zOiaUPK/8+tCbLdBDOibQ+ozBV5YsUAAN1/5tNas1HBNJFcNH6vcIHDazxk8y
OZ1mgZqoA4LDX+c72W648R3BWOSR+vuxlemSyOCygOp6kYYlKKpF7HGTQ1j1Cbo699fJvRACtsvP
e5Lq9uyij/z7oU3f7Qhg1IfzkgzN1s1WYxCwgqQ5+K2jYX62eoUPCB67XiTUx5Hoy9c+HkDmbakF
2uhSWDN3avmj0Vl1YgqEp+Ofu8gO1Fjqj/URsjNuHKis4IbYfuONA0csiQ3xSxVGNzn/6EA1od/Z
UGzhaXcVNTd8N6j0K6IjICC5nZT1BEtHtFxIf907muw0MUS+8OhTiz8ClUggwYtC7hUo/KlNph7W
INHFYFHmXEEWe6sf7v3YKckBaWxJO7VcEyNBnZ0jjefyDJ8IxvtPSGBldY2CU62i9G9zkrkjoX3O
AmBGhsUFSdfFHA2hQPlETq4uV8Yj+huURMImUZ1ilkovS3uq73ucr7qWxLTKs13XnPiFycJavFOg
3cG0F0Svvz1pbttOZ29Qi/IcJswFUiuA6t8sh0UJk4TkPsVJmLNZIHqBWNPvsn83xw5gfD5seqxp
rUvHP79eRISqXlNK6xd1cbO8h1ohNnUxondnGVtIjMtkKVdCyv1qxn3aA0IdcNwtVKVU+CHnlwnE
o6nZ2BVdB4OLrKlDMy+qeR37dkgIZPxy48mcudc+yTOYHYsBJrCeNaHsEMpLMeJ1jaXpBRnwZVhp
cuzBwvzsESkSa1sGD6yUo8OhTPhErg1xFfjxDaSuZN+TI/XlfnwqTmZZyR9hMIf8CYartguRLhHg
csKvEf7ooPmUYV7yil90BiE8vhvuOQXIUYLQ9SnrBhojkB02INsCaGhTtlVpHB2PE6BdA0cYexut
3Ojz7EAz1+TKn3p7wSFPHSIKrQZYCW7vBzmvRUAoLHLctcBW+ROwqHfGac9h1IOGLTdR7zEsq3tV
kzVlPPTVx5o57NrcScj8YhFRg6bddvOfVzT8jb1dtC6xb0H2y4jMNNI/1sLGk4+SaZue3IgKBQH4
2YPYvzFp08ycdE4H8OC2I8vhvwOzz3W5v37xtLHuQQXAGQY8lXua06VctjEhN9Nr2Acsn9iF0Fv/
6l0wuW2rt9CrTPNM+8dVGOoyS72yKgTPAWyUwaNM6Jp8sv2/nwfd2bN1SSE1bmmp9IS0aFIYCc5v
xBLtIzIXjGgysmuPgxBvl8LWd8AWE7w0qFn6Gw4E/NvOAiNiUjFOwQoaQCsr0YpKeSdRM33GwBQ7
bf89lmXcud2Nr2wCQlJq7G1tGEndwqfFqYHqpwFzzzE5lyrgUiNHnrwSclxqVmQyGCnkO9Hi3dSp
L20Al5lXh8iIV/g28g24cBA3vDXTj+kpEQzLOyV9YUi2V1lrY4ARdPlt8BaXef7mC/dCw4BRnk6G
J+mQURri52gwCCE91om14gtpBvJCx7AhLbfhpgr73cnH6CfyqWaaEIkovUDDMG+WhgSUGtFmFUbs
dToTBQ7jVNVQrbr91QUn7pfspJjw7dJbTCJ0rbFMxdc7GytAwfDEn40Rq/OaeDtFecZyP1Ge7cJD
AKVxqMQe1YSEtwk2dS4zHr9OES040epm+679IQlpZUfOX/+0JLksjbydFRvj507hRnucrSeu9IGy
0UBbGI1rOKoiKLUs1z5bgsuqWxb1JrHhB6PF1eUlN6AqjFYV4LrfKCqCG95TILxXxWkt5l3j2/wJ
LXIzuTSs2mQTdWY55QQrE9lkswk9C54kFfrVQvTW5LNBCMydUOkTJhpaKANviY8QQELEC142O6f1
3WLfCI1ikoedQLyolLjswfyRbW4vx2pe2JDm6itw4//ho6X3oHiSbLu+SlEvIQhpEWRquMcVWWQi
rnGRAComwGy8ExG3n6HhckROM7ErMoDxnuln02tdPrtKzxRfgnT1tEri4gMP1+LmA8NX6Z6j2pvz
J6g8ZPLFssCXEI1jOqy5qUqkTpciEfF0ei8a2bR4uipAOhg7gnYU6NrWtHtWrUggxv4ZzNqtrk4e
5UX86r/xsizwaSOwIUrKHw/QVxibKjOY0PtIVaXWMqVUZ1N3gtJgVUBqaY1m5FrVJeRxJ//UQvLA
RLrjgSaXVNYT5vlxdwMJVdIZ5byIsOv/H5THYOyETs2Si/FrB9CdwdSS8pkZizJOxtdliTLfMIzc
OQn+9FkN4VYsF1Ml3Y6o6LRz0KqksOLIkNssYYgBNGPAXHCNqZvMRYJzItjYaupY5uPDxPRODMgf
YRAr9YMrYddhIrONnuKpdpwv/wUl9NYugY7S/ueUFETOG4nhmz1fpN/xAc0BFfTCQU7vPg5dBjKh
uUJbnk8uYSlvRGabQKqNqQ496Tn2aA6p3TlIykXRwYbh60gqc7oMgSA1PWDokuMSCDGidyVa41u4
WnKguPo4kDfBa7MjV7NdKj6Oqlr4m2Q/jIB0xYLsbJcrP0zmb0jxWWKXuxhkwSJ/rjQ/M5QMnGXp
Hda+yFcBdI063Jre1iwV3/npyyuiTEQLOqcSjArZ0DILO/EbmeNST+vU8eGiqcEA9zbFVuV/HsBW
iOVq6ZJC4QMTm3zvd1DsHDMpN5UrPR8IgK+/1hr+XjLBMKUXxt/+96OWY5KXD39PVzykTMXUuupx
0ksWCzo9ETdveR1B73ToqKRlNJsJ1q1OtYA9sr9dnCjlKMdnhCrRtyZVA507cQOAepbrWBsIZfbn
07rYA4wqyc2YLQtY1Vd0ACq5/OLNBMFkXLkFenZMhjz9btgtRlXSMXgnCjcq3KDMP/vHfg53EGVO
f8UxLYXxCmgi3PU2lOtgrFt1h3rMKggbYTeZISuTJEYuJk860boN22IRwlltiNCvEIYBGV18JS9f
xpM/YdqoZPlF+UUaxOYodiACXb9IbbIzT63NAkof+t2DXc3BC37/Wujgah98Fme/Qs+Hldukh8pU
cfCyYQznqW3kMlHB8KIbsOSIb/l6O8k6WkTVTQRT7LyA+wPaXY1fEFKuBGTAfNg3Ht0lPi0rN1ua
uqoyTVrOMLh10x5MC4RJwGCq4dxGMn5hxuk5dA4SOjM/Pn6r1i1k2LrLt4BZnPFs1lv6/A3FFrQ5
VBqsp9WCey07BPvb8s4xUdTdTm26C2p94KDcSU4PTNdXkcFHIY2JEGe+78xqGThm4yFqsnTICWVj
i51UMaBuDz6GhvFmugTwM6Y8/ddu5lVUQu+bZdRvHh8Og9hQarDJ9oVMygO6nVR7+BUqlJAyUqPX
P1PzHdVWnb1TBtNjo6URzTGu3ukaPhzZqdUl2JkdT5FvVfmGxIqncbHE0lmrrAjfpnG1ldu200tf
3CAnU1Ajdby3z7pHdNXgveNRp1DcOLGHzFS6wR8vPTSbV5rn2MkldeWwEjRbkt9lRxNNEjCLCgxp
04tf1FMQXWJHnPm1C18Cyl54hsgYO+w/ZGibu/S/gzX2fUg/3rU3u+wZdi94PWm9eTT0joHYe15f
M6RCB1FyN7XAQyC3oYumKZKFjxm3+Sjy4NptwyVfTXmCpW+w+TYT+ljYRGAMRcwOSEijSYAPoCWM
hBo1vT105xbDLK1x/j1qDT4tF2mgItXW99cfiSwzmE2upmUKvHyvEb0K7aJLdhmyBOtBjsBRXNpl
pEYd2bB1N5lTIKlRf7n1fnWm7FQXU0ehTZ9W7U5QymFTvLZ5Pk/5X0xAAaTPxaNoJ6ZVWigT8KGZ
1CDUixFd1EQYHUpyNV7/pyM9GxqOG1XYM0tZapl4JJ3lssjqTHl4Q0kFvx5r7/pdS172bzBj9Aqg
vvznkFy2EpggOI3Ljqx0wgWFKTe96ZFVNWrLDIks2lfSDV10ri7h+GlmfKVh7XauHXkISM0IKITm
zae1Hrxhgn5wbxVsEAhz/KxBjW1xScyrs3A/mEVi0NNfHxvzODX5kqvEX9mSNv3Ht9azsbgg8bdc
zTjw0+AlyDkKmGvXQIdQvsWM4ySqtK9K8CWHsGSD0IFe7vKRd/nDXsGUgbX67dFPx1uXdmMdLFI6
d6W1P8n0637YBq8BBUCeJyndNr3kYJuEIHrht8fdl6Hh/NGkyZQ1866Jij1ByFaZb0i9JesdhwqG
z9ZTVRu8uQ0OdtmO2fqSkahyX3LtrAX/UTSJUVckm21F0OJ6E07ZxKuyhmpWHTjf/XLVIPHEaIJT
QNHS5TpC25l0IdakmJ3bQvFRI5oc1gmHSPhEizT/DS+0yjs42sCiyMmynEIjRO3cYA7HE3DR0beI
yMLJ8252e/aAkI/pNgMKW5LEGuEfmxtOIAlNW5FHpc7MIM8SqQoih5dcgd3re6awmLrXiNNllVSs
gUQG+oNB9lD5so6oETBP87fKGh2kc9ABfufSnUlt8ES9wQZDXUrjrpcx5/hdexT0n/bfoH3BM7Pm
Gwrio0nSvgYUFsQiuPG3jpYIAGINJ4F9BZLoiOi/3wLh/KVDgeNTjLZE6yaKS2eSXGpNw+HfGOX1
gn1RZFWnUQJnMH8mO8OtaCk2kADqOqlRKUmR9js3NpbzJMa8YY/7pSl8q4LcBmecxMl7G58MQQZp
IgaadRiyof1ampk2V3ohPq3e8u629+JHUynfs+UvjuTcEyHkPmRlftd9A4KfwrBSQ/gayKNjeAh7
8dO74nHwBlRht8UbyrPKFdSpb2E0ve1rEldFN6exMC954oTiTx5J2o8EMgWeY75xvVBr4D/3sNdX
JeqlcjDs0nF4FGfQH+ul0EoPxrkrX5Zvs2I+S+vaHCPLHpvTWcxEx1XPzqRy4bMgA8Io4cwag4jm
BcFBTNpT6p25EQ+QVnqbYE1WV4H2O5aMR1IopSEdkg/uD2DaB3eYk8R6TO/O+I0hia+B/L3z+jXv
/oBNXgvHpWn7xqlzasrkAAkEDkbDw19WFkgMitZwhjI1BGkTjqNCcp4vkLY6YZQoI3jyJwLPNsp4
Pwj4U3nklnCD5Rx+10E65wLclAqbHIa4nmzjAreosQFhnZb9e3ttHE48uVV8KPViY9ShAMISjF/3
9otRtJNxBx3R0fasDbO0xxN8pvqujzg3kJeSDrQBSTfjsRSuss/Vm49n07VGoQhaRdXyhdwWIzN3
E6A/IQ3+nMoFzkzBegsJtnZkrW0/gkJZuQtJwT9EP+ec5kxjfkfLJu8Hj5L3084R7MAUpfoAPipg
yYCNyvPNJLwIKZdj52owRskUGIXN+pmuE41YwrZi6d0LWIFeeNwLUHWzJMEJuNt4phIZloQpT6EP
X7OMhZa7rGW7rVfMU7Jpu+Y/sxFQKVS6pRxayabDHNpk9VBCDYoH2zgFyiPiiqoG2b+EyzR7hW39
XQvnFk1bz4Ez5D62JzFEopLgu6KYMp8BAcswxAX11qLvMoyzKLa1C6ZWaP/aUKZMYBd3CzNZQ0+k
yV/3rbm9TOCQ9+N2/pxB/zmJTdjLcAeXuV9P1mpS9bgMyExGbQ7NXlRh+Y4RQb+AARwUr9h5y9eC
vdAX5v9s6JJ6khsKYOaGNq0uTCD/3jpn4qUaM10dbcO2I5bdZ/7pBsW6e9Nta0XAawtnuKqhqEE5
skqVoIzcqeidwk75qzwljLc2G5K/rIKCMduVW1VrkXeeTBtJkAsIROl+cIz4qI9Ol73aqv05XYbv
f0OaJeRZhquobxmhGjQY0wkjQ8eOJZsEme/BNicd//pwAHBcTqVBUo8Msyth3HiAEYLeKXyJhNtW
22nHeQEhFDVVCf/cogJENHtOhnKPxFEkqoW3n87M8XK3nHF52U+g9WKzbzGbBE7skP38XOHeuIcG
iUUWa5L1pj0SMOKbq4+ZsgJI3czOMO1CTykrsZRn1zIteeGZk0FFC3hlvtctH1vLq4d2afT26zHl
rH5gkDY5LiglsYly7WrHs0gBzQb6fvXMza3RnDq2ak2qhqCqePh0WzfxKXe0D+kAKg/YkX9GG650
b2TfMHeqcp91EqXT78bIOF0MDkWzAhRlVby1VzFRGpuHErCADi2TM/LRkKV+hC6rbH3g8wrbTLNa
JPLS5VfDhqKMKKH4OIEQAvuPuRJbGuDCM7uyDZZZaQHS9nqvPZNYWRaqQ4epnivJkpYQHO9ZCwnE
lNyl0kdbfITXigR6CNHhdiLF8ewbK6ngWhdusyJsk2lTTKVMD6fxvqEan+SKRUokKSXlG9peCigz
mwLJwTpfsya9qrddbvzTEsH6oehhjNd9NH+Z4KMSxqVnCExVgJ7SHg1EIWeW1egOBUDzAIF6LDSc
jHup1UjP4o8p0ac3Xn5EQXmNMXEYq69ve2/Npwugh0S7GhP93Sqx9RkooQyGbW6Rxsh9khhnaM0x
yeVNP22el6ZsizL3G9GbSHbbUmAL2+vKGzDwO7t18pdVKUm2hXgoqK6JxLSwWKRGMctmF60hJw+W
W9Zren6teh0/LubVLXm7cKpkgvMHl6CQU0NVH4EouvkIq+71M7ZeMk4sVv3bUSWPv6fHO9J5slCi
Y1sBKyTMRXEl6D0JpPFtwO8tjxgdRi4FnjtRiQgtqjuw00P3D81JuvJLkjrsVXh9yM5ZA2khmXBY
++q0xbM3H6BpRmaMG15YU0QXCVNYWCa+zP+sZ/3I/HvE7p07xTmpRIn5YE0WdffxUgQhZz4Tki15
ZjVlmJPPN4HEUCd3Ehsiu2KjimObkmKsV9suHirxaEqkq0fEtu2hyn3sWDW96K0YPOJS4DH5ubyu
4y1h6adN9h5W/CxB8bXntOSONRMEJ0+QAhs+AdAUbm6UDwTR2D0xR5fK11Ebhbgz03PvyWoyPcKX
JtN/QS8f4N4ufVS2T3kdynFiz6V1HNOISNjQeSFllhtGE4CU7Z3nqmu4FiKvI1KLnfkUQXf3EWVN
j1ZT62N8RIDbwkQTIOTC3jLJo12BfBLQAv9rZgZ2K9OVJS3+EtNSCm5D8uO7M/T20DUYVU1lY1O2
P3aQPYNCP+QGnc/v1rsOsUei1d2cqGiIEb9+hjDaBROy88OdraddzCCfj9wm8JX2WsUo5T8W5Ed5
ua7Jh8J73hdpul9Mea4Wgsu51FeEGCyLd3XraMopd70fq8C9EPUwqhve1NJuSJN0teqsqGEUJ8vl
U8C6OlKKCnp+RCW6CrSJBl8xjNYM3WlWtRJ4+t0cLs2o6rkfizoWn4YBT/xCeO4Oosu30CzW9qZZ
wMNuPpxSq5WM1jh2or2ZnMRo6a2c5aCA7EgXxz9XebAWjaxgzTKBy+KSl2z0SuPUGogmsV3C/kSg
iLtNsaOH9BzuzJo/TSFX2ePSGDsVZDf6JOgxJdbIiIeGXusst7BWofjmJ0u61RrHxgwEDGnGYbGl
fEdo24qtuVHCj0HQsk8Ga4pFVXSeDDvsiw3SNpplOT8cKLD3/GIapEdZ4U5FQSaZJ6HZuQ1csr9u
CO0pAmnNuOBd6DtQL9FfugyaS1jB9SCX+XYhqgUVzYBkAu6VAi9zb3JB9NUy8qnblAOapo9FK5qS
A4wgt+OPJqeSlh1e6JTSSFPyEdbCOdxgJSgZah3UMuVaQ5E+FvF5UnKp4Imhk/9A9ccbhvf7UYI9
rCS5EjVPm5Xq7aVfzKPzbvlGctDrwyDPJVrJF4h1scLLo3UC8N6KoPBsKPdNxn4kRtvBZgFxr7Ef
+d7sPRgBVVcB0a2Onzi3l7IjQSj4r37Xvb+L3wR4xJKWwlgJpQh8Kl4p9r5c4+9bsMnUvE+yorng
gej4oppSlL+gHfOFl3kSDogYs/orlzTkFmYmcZyssBNkuvqXRi/VqPjjYyf2WPrmR3qD8wyvHrit
O1CEzssHreyfAkuCJlQael28Ptstn5QqGKSJBak8Ya4jLPMr8jM2r/smmxawhpxEz8/e2zGs3Asj
gpo++xw0NmVKUbat835mgYTWRpYFnsq/s02KJQWFlCZE/erKQRieNzBo4GAkAC4KFxi4Q3m3Y3dt
QCduNRG4a2tkmOmn43pg0Oid1lcdHX/myy8QgJ4JX7x9kITYMrxsNAlfl16Jv1wgDZD2vkjoJSAL
rREEY1WEIzbcXws/rFcTHFCd9k6VM2ZuJEzG0RSYVBoJottWBmvX5jDrgG5A4NpYIaZ/kjHgPb4/
2XJhp0KLVMT3bNIb9s5JEAFFKp+BOE08QdD1zCFg6NGfCJXb05WgoPvV8aHfFYM3+8wFhh8h7ef4
dXnbO1hGrxunqhyX+m3+7s9rvZzbHa3JltdivwT1zqvb/HgjjmY0HW8Z55u5QkDH5Hz46lsiYJc/
FoSKgL6VeH0rHRjc9CTj71wnGheiV6YneZUBDN2F9zPJwh/9zx+JxxFXs3a3tc7+Mw0Tz3Y3xtrE
K8qEF8aQWp37AfyYKomBfSzaYB+krSDtqCzEw+BSkHnNCXtDtz2XmUhP/vzkS6HdqMznSgr6HwDN
09Gkul85BhqOMb9bCDE3THmcPzFL7X7mhe8JfM9SKoInAmPWa96Jvg5k5oRbX38Jp3sr69NzGAA1
vOJOTF+n9QYWEQ8/StNphyH5ga+F4ZSsetD3rhiIaJnSy7g/kxCEmXaCyimdApaaP8l0dGd0bvRb
H5ghzIvS0Mrmi5ZAZdxyZ7whq+5ni3m8KfaJ4YoU/HcwNZNDPeZR3RpopVVB9AdgNMopv/2H7qf7
P0QmuZPanWWHlxl/5KL0tvUgeuK3+Qi2N5A+/giZdCw07EHPPjFkiHLkK72hJzCtuj8gVIIiGDxj
119ZmrEW1t33QgTIBmn6lPoeXu+mIy2HJTNGw/7A1ovj0+eC+yv/bhDgZ22rcNj/JfvJgy2DecP4
6ahtk4rrks0k8Vxn4Pq46qxHmA95JvnjHl8nFTTkMbXu+txM1Yd2LUKAfuEdmaItIldEg7ribWWd
brABjMB/01qQu1bMusMEpW+N4RvWtw/aInOJ22DueA3l3prGpslMebGz1RA8BQTydBjlc4YEob+e
GPGH8u/crhC+Ey6XfmiBBoW7EhiOgyuLbnzhuhZFc1pSgkBF5CUUOP3nB6FSYYxcbd/V5xp4OEaj
bOoivzGFE1vFgVzHI33shYM41AayjdImDx9AcCMAMETnFxyaoRJG8EU26gcnxucYQbq73hIvykfa
6kHFSKRiNbMCFAvf5+bNMzA4ekmUCKa0escYyRIdaHHhHZNzyJVr0vN7Ng8t1pdRG1J/sWxFvBiy
QgGF7mTJvWXLMday4VTCYNp2+VzDhYZJzcSJ3ddbIL4kLwj8ksN5ddFBXeRIp99mTaZY/5KZxbXz
D0fOubx2p3lRhj9yif9jFmpzZy89wnV47YJUcbcM+E6STlB51aEcGaLcnv9PqepmGEvo5/R7DKId
Ev1AAtCaksMpPC5gPWvqWT4HZAAyXz309DetM4MXXF7sEpJ6EHO34YnR0L00ZjajuiLagkyToCSj
+Sg0c4H8etsG1BpjlOWB6+df57OC2HZNaXY9Hl3piO8lgMy+F1mRER7KvZy7gXg3GE5EaiCHEfxw
DU1p2CwiAru4BUKWZI2O06OF+aXiJmRMV4+53oTZst6+J3lLz8PfhJHVFz1MQxdJAkxknJVwFG2h
Fwj5XQx/jgTACFc/N5rkjuE6cT40qXjjqTzDhfJIMC5Abq5RFKRVY2jkQrHYshZqoYHPq+PXGcvf
t9HQq/beuIb9U6N1Etr13YMMku3LNmxEUIiENLF8IaIfV4cL/0ewQQV6YHPfrfWP5hED2aLTwvf3
lRWdfMnwuApLhiksdy5jD0AxUzhy1Kqo4j5oopZXVgFMDIsyIvi1chxaJ2dZ3cavArZdMSYj6ASA
qR9QrCh/ZAoPss0232WsIQqjtxd+04oXsXIexhzMJVBfylAzTTCNUSr6hXkKMWa+7UnF7Sk3NzMz
XXYvztH1GeXol0P/uj610kVp21VilQuWhEmmqoQ8/hFoENB3jZ8QwHf8f9ZNsBPDuO4MzPASzgGr
h0WkZUToq8F4ZgzV3A8uuf4HG/9K0QPcw+mCr+ZIsRkZ3rx++HUVdL3oqSmM5iGz29Ot4XJaEKqz
s5dpCixOq8ciRaOBK2t+DjxRMv4jJD/2mceDk8Fbjvgt6jkP79Gui8uqyHARCdo9eYucl7u/7AoE
sG9MeAwA8xKDkDqpi+irjI1wL5iWKS9FrWvBS0QK9WzdXvbY+S12XxH845D9ergjL745sPsS5Hje
e/QsxokRnTzlvE2eh718IcvCCbACTtgcwEtVPSZZa14ZYmUsVin2THxAVf+srwTl2UAF86kYKPzR
8uxHGhjHQoXk8FuWTtrtQNLEh6nTbtXuYzcmStojyGLNthRMisXQ+nAvIacA76zJQ0Kwkb3W/u0H
+ORJmAqvVVkP372QCDxOz1zAjUpvmXy2L6tZylw9kpP95WFZiFtAhfmbPQ+diKBaFf8vnAZVnN/4
48ndfFZPszHcG2Z1OVZm/+B3DMNRnmBLIzw5JqCz+neNuaYTSnPmxzuu5oq5PcWBbcO1FIbQqd/l
iZipCqW4TWjCpTOuk3+SVab9Fo238ZNOz4Q46vga4JeuFQf10XwjrUXbNhxOFYxsk1zdJCU0tW4b
xV23V6vAJsP762zQ20wSmob/CrLEOFsCJowudPT9igh2LZ9mDDhL0Agf6z5e2dRUsvbk/KY98r4J
u4U4vnlngJ8gMIlrt6S8abPGMZUK/xwJAV64UZn5B7dS6CSMlUqusV+MfPc3fxfEp+injdX5HyFk
dNDjjyyoY4IjpBSWs2Vlru5JXMyigTnB2FCl5A8zlM4HH4YRe/hz7AO5NjeqgNG+AqTSB44W6Wuo
fNuleq3Rap12VDYgIJ+Cfh5zI4vpOW5qa3TM3o0h8FCj34NapoyDTECHe70TUC0cwhswPE3yNimU
a/1dfFxopN1PbT7uIeujayk+on66asUGqcWKVXuOuD4154DIXrtWPKcOOm57EoNpLPJJFQYAitvG
q/B1uLbgxoMfMuJmy6m3m9K/4y3mypTY7xCOAi/Psh79JTnm5ECre4mezhqLaS0PNdm0JyE5CVHS
FS9B0U/wKPWlyCNFMLW8ckO7yYUTKV9A77DLfWwyfgEXqsiYyg7y0lLlcEfH7s0M9TizUBYRQQt0
5j1cOYgVsRMaccQUNO0pDkn79sQlzdWzcUYlWEROISSzYjdMmWYsnGYkbL9JGxZYEkQbN8YhQx2p
bC1dFCvtyaDqPhOwPAm2ljvCeHpjWnBC3fXnHtkw84iyCz7PZuY1VRO3Ra44o6iZOFtCxeUon3D1
oBYfdGAoWWVl9ZlQWC09CnPbRvElzTHyTS9GZju58XpQXFiVgFd2Wu8ZljJcCaAOaF8z1v1sLjvu
cYKPBMMd0+WZuNr/dmcq8xW4BnbgOoVWSUyzjjS7Loyea7ho1aMerz2h5fiirWiZxsaIzuGGC2MQ
MM8e1ELKbSucaIZJqJet9qj0D8R14dv/4sDllXyEalN2fl+ISk1L1qhDXyQnP1QkTC0lGZsCI3Oc
Qlmh1JExsfRa6lrXDJg3cE8o5qD1+CTySdFJW1baiAZrxktpW0SixEVn0Pi+mqHL2PcpsOy01N3U
a4H61H59eW1z3P24hFlY2ZE7587Xy/tFRLeffnB04+h10niy7tVCKNcJlfYZne0MLnCshPpaIZUe
/CwGLzL0kJcdPDUMjs2ct4nJalXQ55T1UPEyTyffEhYapsalENptgstM5D8EzmFMjmJHl4PQfGA7
449hUGD10vj/tzteLJULxP4+hnim+5P6Ye6Es7G51xNeXwwunkTV92LTTeet9QVTB2nU1O7/XXz8
kJgY+Y2/L/wWvolTKIJqOA1p/zFFHU0fyajTIAGcDPN5xXX6mRfLgj5Ppbpy6sK8WSDH7zxNRZdm
9h4mNdHp48EqT/qn6O1UxxLpYCiBMeU5V5CX29SU/cTXugyq/n/OC5sKOkWj72GtcdOpMS/YiKgs
6hac+4m+qh5sfB2d+7o2arccUl2ueiHy9/iyUmv//JZbny/iFFfnSwgSVMc7QccQe2jR/iP9z8wj
JDRunbbrFXX6Pg6s5j6LCxibb2eDz30647LtoOC1y4yC2GYPkOJRUStKPY+wJwoE+xWw9DT6QKBa
Wbk4cWpBSpIZwbu+8gSENo3J3ssIeD5tKX9jA/19GhuEGmLcKjdEO8TOe8Irpg3FeRIoiZv/bcjb
x1vNsRtJ9FAPCYrJhM2tmRy+4J+NlRxCW+tnx/njP9oIuRm+8IOB3dZ/Ap5cTPHkNGoCYgyIVN3m
5Z6HB1NzQndWLidnwOsgysZd8AEY7h3KtfVyntOxecBUUrcgx6JO5JipFIRZXRfchBP8+yQPNKfu
9idg+7eZp856NymwaojR/tdiDD3X2n+g/QJkMMrYg63iVlvayAw/W9cf+ztvF7oJiCGQYSABe0R7
2FR2L52HRljxcvmv9pUBCJSRNMyX2w8/V1XxHe6bkDhAZxTf1czuJsfkNGL+6M5fjrDnr2P20Dce
tab8vmP13/5Sqw7ewvR+bbf4OCTDKxz6aTLW0gPDpCqQYl+j27HjHLENyq7qtv3TAk+QOR5M1KfZ
Qg4GyvGTs687juC+DcI0C3FQ2xPlncU6F0m7YEpfPYWAfJ7sLvxqoU3evndQmrxTeNWFRrjmbC07
txOkRFr1fKVB+cWeDIFhuqhnSLwZPgomFtRKQje+Nv5Z41iEF8Ya8KTFVoXn9RTr3R/A/BL1B4FP
Ry/rBjOySQC2ECYyWYr+dMi3Ol8x6xOoJ8+qPhoAkJ9ksniXrdxJZ/tyV3D3z6RGiopqcWon9y09
DCkEpB2HE89gMx97smCFXQZVqrf/fuS2ciDY0GK4zY3bAO+Knq07wfE75mjnxV6L/35uaSsfVBjJ
4u+YM83ij5XgANHejuHTLwajFQaCC/MItUqoR3JpG7SETyZJKPL4O6M+Dk/5AcwwVNYvkwjD2sSx
wcIFu/Hi5MMK1S0KflgDBxeumBIRQqdoSQhTxC7q0SK4r2pVRACWxPFfxp4ExLitBd6LcF8YuKWY
A+OlGnUqqSn+kn9vDRrM8C1J9SMkaleSUmAYWk4gVB4N5jbKVdyRuC8MkNYyX6IlTymiy/4+1H1c
CaVRGh/XtBakXXqg9rGEpxN6s8UAvX8ATobu9BrWO77eZRiNREA6VzAtkDC36M209FQFtUO11iuP
1e3C1me/JWdKsOmUGV45ZeWuXiYitYuOIBq7ebFFjdpdqjX+gF3oQM8bsN6b5OYUQYEKaUm0Po1R
LftqdUrCwNZ3+QW8EDW4o9ohEQVP2eklqcl5V6Q2nVxOVJ+TnWRtlQn90WrzpFqNUquMTu49XzIe
CEI92DjBy/WX6TSja3hMKyEROT5yl2Xo/ewv1mh7hrhOqpCo7AwwR/EsK06hHXLhC/o/Zuz9hClx
Jbit9+Irj/nZ23/vBT8eYjbHoXD954jIDWwihvw3t6IC5fwX4Livfm9HTWNK5PPh3krNio9f+AzO
TyHrHbWiIWH4bNcrMPTUXskrMGElraO8zDUOyoIucp6pv2OyQmxU/nD5wvkmVQIx46cYk/bZkpG3
A8uOb42+9Ti5lqLWnpqJUEqqmQwwIiUfFUchJfC0LGpgbPgh7590j0zHeE7e7uqmQnikPfqQZ2d1
7P2ux3jAgoNkQyiV0BkYmRVWIMrltGQtxX0WkAWVI0Nz5QBLoQv5/t1ieKC0Z8dj9EWtB+tcA1aF
Z42dnpuLI7HwTZmZQczCzGT5kgQ4s4R8Mnk4qy18FKIp5ffLTCj2o9vkWSd993xVDVB3zCpt8axN
FRyVbOnCnJ49Eaba193W6xR+VoCHX8qJuVeWQyIOBKmxqCO0Ky/ulwJD32QI1alifYmMRn1Xa8Rb
xJacCUQsIKgdIeUEzsQy9Hi0YmRBA0vQA0lPZ00FYD9jFhj+J5ETXZYbLa9NF1dIZq8xrB5alpJ1
zkZoN9sOly1cJ4mGUht0XEK281seTmCm/hq7SR2fYdk05muGHscj+PtjYojIXjNvDDkrrLMfRq2/
d4YNb47sCECRNQo2qqD2o7gyjDCkitGKTIw/7chxD9kQ/8+lEeiTEioewvVur99aD6nWf7xv5e85
Cq8XazYnv5PblmuwJU087qW479SS08WRepgyHOEwBssOCHV/64tPutFvyocEdetNUOHVJDwbL990
y8uQeUwnVwleFkpOocvgl7NPFaZ2ARes4TEPBFqXzPa46v6OncjE+hX2JafG3/dNJqzfZDfKkr+F
kykBJvIt0Swo2U/3BJ6eZioq4/odUyzsIoa+Nfp0ElPyBLPrfjrlfvY39GWaJiFkLJV2j9Yc+/g7
LSLV6TaNo8e0KZVE5iuDbfg/rUaeBaMX+rAI5XLHLduc1cpapjiAD51v3LvoMnQaaQQjfCgjW1Pl
dshvAyCMVR6h5On1weQcgzFnp5bx+tsh3zBi5A6/MdusX3z9NXIpklABjkeCjOwVJ3l88a4MmgwR
GJ1piXPqWEYdxqdBU0nkUFynSWvBKdkaFnAsbP2yNedsicQIimECu0AVEBfBUpESBOcEBhuWUSiu
FZEg3WPawrK9+qsyWVtF9TRrnn5tkfKfJ+fy8TBDRnMsLZ27xd3QxN0zV13vd932YlLCVoMSC39c
IcNyHkTEkzmcjtxfxSqt18S18eH2bRINJ+alGjNczyG8aHEC9vlG6+rIk6v1zopvO2A2DWnjAg25
ti/tlLVHDYxK8cfIxgwYHj2LxvAJnk0ieDVf9B4toHkwueMnyieu62lLOSruHXQF4WVaHRXZxr3C
Nb/MLgSuxWcTaGw/2LuW6csoDGKiio0PiR1h8stEFGrT9xMBvaip2o0jaxOhC1hf4GNp/JqtaRxv
yL7TntWtclTIhF1rhefpC2wGqcmZKLa6TXbyYoX+N7O+uff+M83Yp613pGf9wb7NYNnab89xJ8G7
wKAQvKKEiKdUwUiYt+uMVKZGaJzk0q01NeylA/jeSzTvXTmOiriITaPjIw0xn706rnYddkK/w+cO
EzsMZQUkPvkYISIIDr/BuwIXmw2gkYfVRdSoJ9PlCx78vHCZXbU1YkL5cAMqfDUoqBlkPhaF72Sq
U1a/4+ir7U0i1nrwin+6Hz3DFnWienmjBFcLg1zR4s9AWlQZDDddFqJR30Ytah2GR7GSxkHUkGis
678rKBXiFQEsTl4Z0EDSUfeirUE5oeCeTwq2K6V7/Otg7av6qCMdRsEpavtR+6Tw/1p+gzslZt3d
gIY+ql5BWQECkVrRRXzzxAcY4O4NmCVlCZRNbkEOoKlDHY4sTbiGv5RPWrwPXIOlJnnciFgDfZgR
hjsu3btD9Md+6FfSIHIsWXgzzPVXSJ3pGoFsDjIW/YXcU0EVjxrKBOdkpoev632dHTXI7y6uFeOj
m/en0/tH9xQIRMhLk5XNILLow6D/HbjhqINUl0H3SfGVtn5NBcWOwvBp45Gj5N/MXALvRCCr26ea
pscPswNVJbmtlmymo/q8E04RseNn9wM1KWLMB6Nc6SIjItO0W1rpmZUPvryKszlBDL5E7B3ZLfRs
Jdv663zEKQtrdGER1oQy2HiAnZyVtuxBjeiaRVLezGUKB+/SFaFpUrZF/PL/SqkjlFqG5LFaSVZS
eAFjpiJMXTose6sY9HFKKblud+sq7cO84Z0u6sPR3/gYj4yiKInz2yU7GhD3u7N2qLkgQ/H6nhR4
mJ3UbSoNPhwtm7wOpr/pTdkwdKXzg5TBclev2FsDe0xXS9Qe2eDf9ALX+jnxZmSlvMilg69YbOIQ
Ju49OgEPVkm890Y/Yqhj9PYCiJIdDxY173qTN1cRaMMXF7Defv8Lpccj+s4HITTF+ZmylVQi9GY2
Lf+iHFjHTQEZooQk0UkxJXecwFekAM4u+pkR9xbcaH4XUnOiEpT/Hs0gyTX7rPO5QUJc22Q4O6z6
JNY8Iuf72ZRNie4pwKOla9LJfluuPcSYVKbKEDP2rRUWmzWrlwDr+W19z0nfWyWryd6ZBqMQxPvK
BXOvvZDuWimLd/HESw9M+wfMaqyCXgx86azJomSMkV5YbtSnereVHLU0DNtdzz4lK7VKxjynz8E7
1zg5fPR4VRaZdvfu/wal02HSVGtenQkFoTcuu+rNdnfTDit2SRg7muPaXoxF236X0uxyfxosERAs
TBvrx4a3yER2VP6pKluaiB0i9hNuJc6q5P7Zyl903rH61QWW4bMjHndOMsPXCYlYnG7n+yv3KKmR
hJsIpdsZTcm/mQnUBm8e8JRDh5eA2coxY/KGaLo2+wC1sbUTV7S5yLRD3qt9WBWf+EmbpkLCgWsH
TSkdaxUHt6bokzLZdbQ6QcSSqR4MJH/P3fH/79nmTZaZT7P4SNZsj2ygkvRezeST0v4RHv/Lc6Y8
xsOLdQBD6VYFCGKlf1wcnDaZ5hzcf/QnpAnC7Ca5MqJqJw71WBrdq2IgMgrPsiz3lH6v/3TNpmoM
jPFekWvwCold5dWJJLw8w5NhCwVBp1A+HQugZXoo/gyqxM8rcDMK2aYRqWMvbeAD+pebV3w1qVcM
nvxB1o4QYgmsDkpvGYdYLuqutmlBg83UDjh5GwesIOdyvumODMv8m5+hZh4+OIqTjVNiCNX/cj3y
IWnt+SSJXmnTeDAZVqoThtmvBjHGyaMq7o9/aOisEpP5meHgEnal21k3D/YqoDEm3CP+7R5OcFl2
Lq9V3jN26oRb4fUJzR+Zd6BjH2C2GzMqAtDaq6A1A7OfKDJhvuOl7ql/MrGgvRhdpazRI57ADWB/
QBfJeGt8G1NcPpPiXvxThtaQVk5MCRv7Lpetr86GVndTiQI8INoGVjERzbLOM4k5bIJeV7FtvvQJ
TCEomW8lhl8TNRyfZRcf98ElYxnE3PAwDoAlhY6C7DMBsWiJ+x98ijIVBXzdegfaH40eVJWHidKP
hlX7W/sDlmuZiKTudeRUFZBm+x9qmOXgcv1VBX5FfnPfLxpGwf0teinWEwTCV5zv2taWfjk+EJGc
y85yoWtJ+ouoshE1uzpwOfkhuSq8cyl6xlbhVZ11LZEDovZ8B0AOdpIP5o/VHjy4pmYvBOUg+npD
+QhX3hQx07bzJPPuUmH76mVeSUFKGpAtA209IEsDcuJgOqlJ1QsEe5GkYK3whlZbg3K/uTjQNmsG
ey73sWglE8TXhWFRohVQLkL5aF0tWgDspR4K/7L44zr3t0b+GXt1FCMo2uAc35LrqIHnayfsjRpY
Z0G/0oNaZiSs9aF8sOaUj4g5eOa+KPlvtEkq2uEiO9pSQFexytBnjtsXrxK4bFH1Ej8/dESXDEzx
WVSRpcTF9oQhAWSxovAifAg/Vpb3rKnZRV/YACPL5VxpxeWOWJDDEIbeLpS5UbLm3QIuE2Co//Ga
sgKZkWq841KJmTVmalWQSUW0MkRP+IUkjL/TPhsPLocQw1MPlDBZFidW7DaTUQoviYLY0YfoYGxr
q99PnG7DkQ1mJzKU89wq5bfdrMqXonsWc3w9/Xjik6BxhvJPh9Cc/fkUiUAVMn4kA2lLf9sMF74P
ndM5y5UQfsY+g8/m0ezw4zcPzYyQsD47l0Q1oNWM2vC4VRz2VaAV7ABZgEG4OtNfOhS4k2j3pw17
cNPqDRrbVS4b0Tm7XOdpGc9lIwh8iVBerIVHrzM7qEid3yNhOmNcPj/zZlQhwK3JUm1SbZsnhrv6
8hHZpU1uYegLSOr//GmzOObiWYAVsK2usy4aGTiqAadSvpIUmT3LxDOapuMmiYWsjRMQA7xnrYVd
4hPZBM7ZqFn0GD5QBNKnIvFovXwyWDbtl5AP8/f/xcCI7ch8EHxXwv+tY2talIlOvjoTiauhJJNu
RILoIzqt9C/kcJtoinxTPQaUaUXHATt26IdFJyfHEEBVqzcRGBszVQVGAmp4PHA/4urf9JsXTtyA
+ar+37ySfL1R2V3LndFaiMDagXs2m9m8W4OycvDen1mG+LZU42H/TnlqQXKPWZfSRecy5++7fj+h
HBTVgdm4eMiOmFDlDm7pnCOGgAzNzxZcYD4Z9ADAxlRQl1GcFxS5eFT6O1TRJTbRj1D6IHXX4zun
8o23wtSVyFmY9C9gBHEuIdBfqgBDpuWFbvfKELbtBlhXrA7njmcj82ti8yaOX6FfUq9dQ/zcVRxS
KCQ2SEjcp7yyMp8fC2/Hgzf60iFKEGAonjFGhHRJuNnMx8Ukje/CFKifzijDRS+TrZSWXKMEudR5
W3sAaod0A1Tgj9Dy3FO2YT59VWvrletxlz+ZPJVIzjDHL1KABq66p2OsDchSBUcpXPWbeKM8dw6n
bkiZi5skK5+TrkS+xyiexgkamPMg6FcsMYJi1KFNh5NiiSae8NcRAoXvqGjt4tIb4wIbfV4BjHi3
HiAh6MVmUv3L9VqqtPb8PrCLdtDB9s02MD9x4JosNHw/zL6wwFXH+Q4RTTPfp1+XR9A1QH+93q2C
Z+b9MWkWIh1wNq6SVcMbPW4zz0iAHMdZYvJTCpV4B8sJmFU0XL6+XXXZQB05dO4W8o6RCxWW1Q+M
RfiIIUFSGz84s+xJ6cP0lR4mLKvT+bRgdg2T9dumPqi9Nr/nxL4sCs/BD60LLoDcyQOXOTtcPgOR
FTGOAs5D0kWDQzqauWWLFg+ZnRxd7JLYQBYVrbiXYMnGC7QODRz9NA3M7TxNH9zAqAkRsbSZ4Gnd
z5SFHKnPe+kJG//PTGYHmCXo/DGgavHOIeGDpjt0YGegVqi0U9laQHM7Srd977rbg/ch3kAbUP8y
nVjZZLg9KqM3smlq4uZc4fRi0r4ispug8ZCMW+OTuVAtgKarENl8MguUt+oOYejBYFHS+jARTw6O
vUsLEGtNHFIFLxgIteKDiyNZkBm+2bU7wHUKZpXzSyiVba29uJ6rwm76NIhRMxX3aDFoYVvfZija
CLp82LX6t7LJacnsnstfRjTtemMbTftjZ9Yvt3wbGX+E5GiKtr7dKi6VJYeHwK6t6cdotJWIEpe6
ri1zdlFeHswWc/N4qCoSCLMkn4xt/Kato4TfFzNshZu3zfsMq4aFsXVyLoDAR3gmv5bhaKBmewRi
MigUCN9Yqp+PULd5xp9ATqU4vCmitatqWOWJbhnPp0duAkY62Wf1mpzvWEIhWO8GnIW+hSuIuJ+5
qfUyzta8jHAPhbzRRV3HOMa+NHmjm1JqM6CnEAABQuDtiuTPX4UUVhAaG5YssxDayQEI9KpkIWWY
+WszhLN4iyrZn3+Wteg0xl3CwGQ+T8X0IeN0KYIYWfQxv3bWWGQfA8wjrVQvY6LohTvouEw5PAOx
0TEBhR2zJxRRiLM6UFy2lydA2niSWjFCBtlUFRVk296VK3ETmuxhWiGeTteXa0kZEHUQXQPdNg7t
0IYJxUyQcOmJJl2qmT6VY+Ot3LyYGOZ6c3N9E8wi86cXgpLXEsIKxAFSiZ5TFN5UQ043L3QVtJoD
U876ycuIfWRyD1sLRoG7DeVlL6bm+SNU7KyIVjqdwfarNM8SIz9D+4Jfqn9jgSkcy0huvwRAS/HT
RtcpiQ4bVnBa8bpqC0mXlncMsk5I0XTU/W4or25MtrJ7qzvgueUq+Y93HGAayAIpqBxHIfGM2nOW
iW0jTnXp++9pjqsIKzp6+49afOLSESkmQbFg/Sotj0sP3u8tznpeaz2P+HmCjx/tFgV8Pk81FJ2K
wYIP/WIbz/d8ey/+ZvGStPIOYWXs+99Oj9AwjgCloWZiM1UYDr5SlPl+PJ0s1Bse/cBenKMv/DF6
lHTJdNk40vIDvKUq7tUJxDlyEo91VsSNeVkeLLyHzb5q6Bc7fUqYEA1mYtd64Ibo610PvAsB3/nK
l5RnquvGpL23y/pQigLw4eEfuM8JuvdiobyglkNltIL1pt3y23xOW00pzQ4kad6FYOt73hKNDdXf
PVNo7YMaK35N9EEXtXI9oOzL1XQcc6kafNucyLdN9HHllKVOGMqfZnLNcnVydupRMv92z80WboDj
AoxyP6v8muPbMnBBS4OhtBDtpGrJadDwda1yBDRG10xza3ut35zaLqF3gS7GUNUx33PvFkoJhZ1R
jUz7ulfoErX8Xb5/Spi+amLi1Dm8mNXcGsLuM2eEbj28Lp7XT6Wn1oaZUJ9lfVSJC1TKnm5oqlez
TNRKkcqw1NSkfTr6wrjebikHAf4k3EMESmUfby+qTrvy5fHXDKpNP87FM1AFQa+jsbgZQnpJ8Dyc
80FIDHRjyzkWeVKqaCDnqK8/a0nqrlPBgINCcyhzDSGI/xFGCVkZoC4IAaBY5XTc95Vz6QEjY+ee
vxeE7B2pIGQIpPnGlpOHs7AZa3S+Ib7h4FmI+zpWRQQgJNqHFZEbdrcr26cIBzym+FmkbLUqd4l5
MySOIedQ3hBg9ctQYLrnf9JIWu6cqRiOfvBtBk2DSUqrxop5JmYRfzMrqeBPxZRvKXgNmV+PsD8z
GMTLcvFyv0uBtJ6yReUlyXKcRdwRZpVgVIKfcrZ56ptmm3iqPCbt4xcwpLZBnR5iFzIixyaQ1yOj
fQAbGEpzLhiH+ygIcH7hG2A71brKwRNgNyvlmmcHuKIM2BQUrGi8uNFc+BwT8nUkL9A46VuhZI6j
SkFXkRH//bW4RyJm4xVfhVVS4JBlqfzxfEKaeyPJet04Gylt2Ma/UzIhyNB1i/5i81fYe5ojQiZu
0xjU2WARXv+eFjBViQnVcx47RcXjUSGOnlT4OYFIT2mSsg2auxxEPJ35HURgzCrY4CBWG2qi+5i7
aSGEqQ54obi/qQm8UUivvaLWzTA+m2K8lmMopFEfs8hbIumnwkn7fGhfdiQzmK9AWtxvqSMH62dT
Jc9x4QqSjBBUUBHrzcg7rMb9W7YTKUG28Uu21TQ4c5yNh203++uFThetuh5w+e8zhLa4xvGNc+FA
t53r8anda/WngCQyxUJYeGGO/ors0RPkqb2MyI9nuu9vicEo+CJM77f5vw0OBj+jQuyaYBsntjak
vS3iowy4WS2P7YMQH/3MlzS6Qc6wQ2MSe1tTHmQ55RE5B7b+w74OlkSdZNyzUiWDiEkLRohiZUux
Yh/e+nsADTu7m21C0wnbvya665XMrI4XVv8LIiKKjtY/CMAnVqZQLqcPnsVaFpjgZNAjCOXaODPE
juU01R6+aM81yyNyxwGjqwpLfkjKHFknm5qeXr2CCeOOn2aw0B76asnbV2ETGzQNTDAB8qnlZLp9
h94Nqpg/+uH/Ng/oQqR9euCchwrRE+S0b8ydZJpea5RxCG2xUM46avg5NSj4mWCSEYK05KnS3WtN
qo9uuoTbnfskZlw6XIbjqL70TZ9EMxLzrA+5WVQ0FADNjeApsZg60iEyXHdVRQhcFJbgN7lO+caT
kbBwcTl7mK7tf66BhXDMLqKA74pVwBDXnFVmh1vMAvGdIkN8omSfgl9rR4fpinA1noqEdP7JIJWi
WpkxanPI6rKbN+haLjxqSV9x4G6jWj/YzUiwY/qsXY4UbeGo7Ivm/QJ4UdA+1ajvVAloEHiApcT6
TZLAnIBJRuca2MvzEthjqm1ZJFWJpEQpX/3ONcMY08j28hkHtFiW4jEJvA3BetYJJoZXqdaR8sO+
J6d7vk6r0WNHmKBxqfqWJflpGqDckpODBkb/CcN8WhU8yw1fnL0wq244gKm8Bd6qQCUsRRICMfrR
8VPzMzHKnE+2+QtODTDFSsKmW4qjrtq712UhUGIc9d1BfIZy7i9Q7Jbd7DivpKqfNm4IafOAHoF0
xwZZutLqx7V4q2yd4ZnrR9RzBDKs0mTyNwDVb2dHrYdxiR094Fn7vuB3Hn6rxmOt2NvMfeuqWeNe
vjmHKOY3GIn1Q9Aeois/cFg0Z2UXgtzDxeMlwGO23O9UYq8uiNbvYMNACQ1TyolqWQe9Rfl6S3PH
jDZ3qm17AqhFyiIW5mKaQoeLTbHIvX40jnGWEwsFAZmDiTmYxT/ImORS3SvWLlfFEO/V209p8/F3
Ry01An/3oFxc57aZIbWU1wGaUcVNCrOJB7PRGlzRU+Ub8KmxQs030DZYdjH965fxNTCuwYy6GDJR
QPIS5c3TMd5noq0Ojcem5asq9KmKrk6tLGaL5xS14kXHjOajI67ROxls/hFPu8sQKRtb7qRFyPR/
8TP6hfoXOSJKWyaz6OKtRqN4mJ71W0zbmiqPpjN11POwWhfKG+eLexk+YfrvB613azzWll3oHIRA
JZRXxVAgwttv36YJXvluxlBXYTrhvNlWmi2MfBw44iN4W8xFWMbQ0NcsBL+zr6VMK+cJRgAlG54j
oXJOUwJ/TMvzqkjDT22YJt5ttNzbQ8WxlukmulKT/w+W3XePtetRPWhW/aDF8cxYympnUPlGAdqU
T7F4FC+D7A6C9SDEZdIrIoQe0wqb+dN3XO2fr7n4Z9li4Cf8ae7Ybrotmu1wtd8HZ4ca0C1jODQN
pDnwDhZWXEhdlGm8RtB+bgjzqRaYhUnjHy+rcKW1l8G2j9CqrSnoty/2GyMdojNFJmZe9nImvcw7
DMgsmbktfrom8zaPqmrdQuX4W6CbMFUErOL/e/q74ssxpU7/7SgvWzR0Kcgm0v86tk73Xy/K/uOZ
vtTzFlq189vuhxUcmXq4nq646CJ6KxU8HGrrBqtP7uRpJRjN7OUq8DSOVnQalY+tgFi4KOefmC66
bczfgtxGGAYpziTlYPmf6FD2Q8Lzfby66vKwNDRJ77jPipwcSqyszuWcUsPSL5OKRmNdtlsa9hHj
vzqXjS23YSKIlf7PZChHP6YWHyhfZH7fTJcbpj+mGhLiJJJ/44KuiAZTG8eN63k52eWydKtR33Nj
0lQn6blVfk1ekYyQK81Gec3BvI4l94dSN8lgT094tWbd4VSlUP2VMBHD922FsCo0cv3O0aBmOI9D
PNBcuOJmfez76vN9JKZJlH1sgDaLLkV+h1DV2tUwDuoHMygFqUHWRwYfLBG0kNs6VwXHzDe4ookA
2Z12MxNTZWyKm6kQzhpXL31xsqmmQMvlMDKuPr/u7lE2H/Qo3uthjrv+2UhO8hEpqsHal+vjNGCr
HYs1Cl+jdqMDPGTK/D8vcF9/usuSYj0ragW7CQPpWv09otPY0njTvLOScmk9EIkWYWYHhYzy23fW
OwBarOt9+UjBmvUJwpg7aJEu4GUr3D3Nk/kA8oSLd8xbbQafEx61KqUfq9K2RJA3zW4xfzbbYA4G
BGLwfA/Lmq6VFA+ePLxfaC47EU6Uh40Y4FDqpij9AQgflOg8fjOIz87xryt9TXUphJuPMimGRMa0
z+XSHpo3OWDWDnMT6orefZHyx4FWBYZB66cPtCu3ZXNIiK0ChIoqnhd3SbuwKv1N90tdZhv66AS8
zKc0iGE7szOztOzdNAeLvtUsf0exR3Q/3Gpqo/oFKVv6qI97muCNnDjyN2awavDRavoGFmjPuMM2
KT8VeG373eoITlKcE9wj9u3sLKFUmZ3WENczqjbKRrN9i1mfYWPB1wZjWiewbQnaUHbVmSMvr9zQ
24wqDPOqcxPc+zliT8bw4cyhcrvzwsWdoCd/C//1aTbvWbooheYCdhEAoNg0G3PT1hs5Vog8shQz
xNRejWiRoPVtbrW0GJKG0TAJrXg5tZBr9pwoIxXAEiKWPlpKUn846Rc3S+lg+ucuTpkfcYjVtJ1B
sDtRNMFhq8we7EQY4eurbS2WkppyyYbGVewStxyGQOg3oFOa7qxsJFFzZjXGopDle/9K9QzEY/nq
lzI2MmrJURySCS5sydvOG7tcbWEjJkR2FQabe4A4qkGIM972UwQq1L/poS2ZMggaYNgQiS7xhJWw
oGXmKjMjnlqbZyQjnEc8QE+uvVweJOmxGEuVFshPGrE85lFCzeH0Yz2JM+ZZfgZZBXTuBJeSNHkj
5CUdTXBZcLWxFu5pBoVmTCE8/ViGFU20HlkO05ZcvBYx1ibgfcT8pDvS8audk6wzrTirPRVJfY+y
poNQ2+VzO8XRbZJkvzPpm2+15vGyl6ZracKj++rB5ted55EaONIW8xunkNeEtK/KUTzDywKmbkBR
4Id6v7KsOgA5ASUwyaf6B1ANfsOTOrpsMUwBvQL9yF0jKt5VmBYGyqS0rmP6yh1c2gAVBDJJ/Lnw
rm3uvi0hC3s6YU5id2v6VVDH44H8d1UlqFpbmQeDXSLzXWx0WtypjL4djPkS8e97E/ERP1P9sgEl
eVtxuoi7ZS3Xk/e6uW6BNEP+Qc8YazRXL/ntDv0FEa/3um4JvGrAyD7FihDoveaNpmEEw3tQXb94
UKKsxtpvBquq8YCb8go9a1gQ8cqh1xDfREo9GUqbGwEEVkQN7iDfVJB09E+6tPNR/0cKPDMV7dH6
A6tBiLxO66wPP6HQrkGkrjo8DdS7XczUj80ur38wl+J5HiBrF6vCVaPgGuqH53/d+rlk1hg38dUn
ru6UnjVwSb7tc0bPc3pXDDGCbeZJOOA4PyHpl9WJ/64f4VkHr4kgaWeCxfR3vts79RuPLMviI/ni
MnuERqrj/0WaUXoihqaRrp4jt+se0mdUH2Rl8qFPjA9ZPFuolxBUYA5t0LKN1cYQyISNKAQ9zRWV
rCFyAdWkERQXeytXvuXE9nAv/+c2uedHtmVS8vsRML50WKg/OV9QeblR+jXyDbYnxCx/wuFdUx11
Z0KNS1jgSqhCmACYMhiH4Aseb9fRDMLhiEI7ok5qS/GIl4mId/qp6SHnmRuenIq5fM2lrxzU8qcV
ctKfJ/gwm2Z4RfjMBHrWJ9UjCr0V+rf6lBWSDkyfdVC3UEmbXvVxYYMcRg2yUqfCBzQ1TYdRrqnP
nEd3oN4WFs4/vzY8/DhwBf4PajpotzKUgI3bTsohFTK07XrtHID7+2DLYOgs7jXl+6Hk62IS/Wzp
fkCMkaOQPtMV87gBJ11iBbpDO/LJtrE9zzGLWcxO+YdysSZcqABOoNWUOy48NchOiObmzfvGk2Qi
0vR2JyxCr27PIDKdPix+l1QVf5NvYKSnJJ7TnZVMFVH5gC89+Kl+hVxRjBv+7zzPoQhg6vMIJ8k5
WAgpKk4s313A+YdIFBbWegx83hYcwYch7vJ0cMexz0XzWGuCZGSHpdQTNX0XBOUAJa09nCsSoa55
TG59VrX2Y4ZWwKpLC2r3UyOotCtD5Z1HUA40Qjw/r32X/s5BU7qQEjzGd1WHCa/53fLR07l36HDM
NGqGrs6modqnrZzaE3xBqpUTBrSeHxpbchMtYt94wXxOBzaUKFR/zR8o8+fnZx0U9RNnOY7ccHVP
qxoJjGR04XBUMIj37eGwe1KbK7Y3ztvVsQsQ0iviJCVao1sPJ3bd+5WXzfov0gTAWUz1yzR+1xux
2I0pPJk+xJyTazz+Uf2lHOjpTAGcHZrrTN8DiUdjRZTsLDCZ/QOjyGc3/tG3V1T7bctLex0zBPQU
iOvQYkvE7iP+GxClSHzFKIBWMVxNaGggi/znWwr+lpeNw2ejrtXy12vtmVF0exxIFDDSlbaobk4i
fU6T2NbA8RrEBtKYBKk723SntGZt+hLb5Sp6LYXKnih7dhbnjq0Ib7LiFxF2HhuOjtyLsC0lkHUD
pmdIW6bikWgz2r/IljfImcTAtrIeca//3E+Vk/1WJWZnyP00Yn39nMjp2fxmF0pZttmgpXVubDSX
tCfUTX7V0EjARmwoQoVgvciqzXo31kjLudC1aDtdcyfsApLwwOYMkETHH60L4aVBVgBQ4hCH1FBx
glfMswrGn/hI6l2VLW2e/+/yQRxHnyoJ8lROg3AdW+j/zdssVulZo3KnAu43AuZrcpMdD8LldP3M
+j3Eu+G2YaWqfLT66PsebPjzhXmdj1bvVSAM1xsFJSwW1Ku5rOzSCcqXQDVmtZ+gcnHFlxdIPOwl
ybSjbxMVxyg5Yzx9odrBsnOCVVfyEJng6QcqQBg1oS6h3kK7mLHu0J1h6HaI4GI8DDe3rJNWamIC
yCcUxOtlIUo390+rRrUWT5gAThDroCBLPlh6trVwR/+lyJCJu0sOY7QtHAhfMGWxj/Gr07HHwoW2
W8/a/VYRcNmoRcnzFD49kMoIF0rvdlV+asC2DAqcMjtzCTdlYuDj92Kj3+O17ReEVMiiVBqMBtlC
pxtByDcOY1WRhF+4yaE+OO/p0jvIkZxKv0pP2hQQANWIRCKZMo3amhpj6SgqT/CxRWBdY5TuM5bI
MYEXArhBDFOMwt9DpNNMqH7YTzgjt7BM1/JSKwzxeHFL9K48dBqHcBaKAA9uoGcXFmHxo7gdJrEF
begCthtozcECeQL/TOpbPz2JNcS+qZsMNX0uxgCYiC91oGpWoFje7BDyA9T+m+cIGeSnYxajmd0a
UgS/Vh+eGan6iJmT/Kd3k4Tk0iB+iwmzyur9RxT2Sc29R1t+CzcGKhM++qOh8Q4GKK3U+CGt6ukz
ibdkXuOKkFNFAq1vPjCHKU8VMP+Ph5LXx7fHw26a9phsQY3muSfzk+JFPxTTdcsG/ModwnEH4+Za
XLMNBpP0VwA5J41xPdQEsiNN7R4y4zmxwCj8LVTPdESyrYQrJ5NoC2PX18aDMe58fKRGedUwpFgs
SxGRao9umgvq2e7IdVndRpO/nbYziVmxvt7e8qvduO02YME/IXBv5BccjF3s4h6bJxXpKtdKeH7U
gmCwJ+kNks34HYWvfT29td6fEMzZIvI4pdeF2ywe14LHDE6jgehXytA503tLCSBGmxq4ApBcAR03
NX/019HRl27VxrR8kzH8+IeKFgPInLyRuGNb4RSKYUnYMffP8tCtvO/c8ag1A1kaOWcvy2fYOYy3
V1ZxuJd6txhOScbhfcrYccHdzJChbT6BsyPwurDAakpYJLFll8ERShqXFHqBlCjMQJM=
`pragma protect end_protected
