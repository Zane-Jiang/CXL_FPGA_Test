// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dZI/xZM5IO05dKLjEek73wrXP8j53WuxLSPHlg0Z7eSkpsH5TTbs5liY8Uhm
vJ/TrVH69/YTKo5VHggQ2LO6xZzQTCXdh4MRKYIpIhKY2O66w4+HA+s5loQf
bOv1/ma8pblAMibk25jo5KXxIvh9uw3kJjhMA6WO2qNwL1gByelosEvy0k/a
dQysxQlHKcso1s/MzyJubyQyDi7cmWspuqptIvRVLDJisIvHvBYl4dl654Qb
fLbFNk/XF0AbA9QMcboav4PsgqXFiVRwZfgrBlLaR8HZorNxXj1o7WaR+tIx
2frSaphQ/Dq+tJZtdIbGxtjc1mADJQl6GV4DYEMdPw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
olDyDw9cf4gLqZStEGh4pIQ6sJKZDB7+LuNF4fLyzDvU5SWvwS0UMUk7g3MA
H+DIAvHV7X70seValOmpZCqcFk+g/sGB3KLl4urt8k2CrEeEVKb65y1heodv
UtgVh81uXZTACzmPDTaOEfu3cyB2ZjQzCAVWEbhSRIECTzB0ZXyz9cRtxxD1
SOkDR69bmg4qGL3HDAENaj6gfgXwDJdRe4jT0NCf51ga42fPInNmfV6sewTz
hk5/zgt66sYj3p+d9w30uPgqbUt1mG7AvLJh74Bg5wDBQtlolOYCi58iUfzE
akUFEVAXxG+DQUX9mbW6XiIF6MGeYEBJQFqSkD3JZQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NWXjeRH/+XE+xN6cnALP6jksIoTmKnxNE7Pamx1oqt+NFNXuwvWfGA0ZvilN
X73hbYEhhmoHGKvQuL04hKIWkWIEr6FzoNR33ILIrn6THA/M93CWH+zfa2+6
ekVxu1POM7l1jQESsVYhDgKMyk49CrKeGbWp4OfKu5CufojT5G1t7yY5Wz1Y
pQ4HDnNcmXnM+WtRhMg7LDk6Yedtj6fAUpxTbHp2rLqMvjenzI8ktto16IM/
tSHpocGfSTcZ7vp8BAcRvCPX848xYs0xxzBtmSK/2GzaLO/jDQr90R9xpsRr
eo9Cny2puP7UvVqOIquM50tLtwqeadl7goXCHKRYug==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nKRd9wBHnuDsjcpiatE1MVkjskT3kKSQXzwiGmJ5F8vPrM+emEqp1WUCtEaG
VuJ/s3FbQ9PjD7icWEOsKEKPKktXjE/8Hb8PEFr0cZIF6/G9ITdRj1vW1zD3
Cls3M1C+/5Hmv2fMIxn9LcnKDPM0ld07WsHNs2G7+15MWl0eHAQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jMwVWmtAQ77Z1AfQ7BUtoXk6am7L8EG1uyh+8l6112SiboXq68apwOpm7k2R
smL2G2tX/VG/tlia6bP4H72vmfpAYBLOl2zzGY9Gzr2P0l3QxbiTBThTxINA
JT6b4FDtb27XXW9AZh8R89skS46hHswJ+EmOnw78+hLhIBsNL3Mz0pbArsEx
Jf3g+XWb6nNbQ8c01BMx892uFqS12aYntP7YdWCt5GwsBLEfzU+Lsmredsth
xEEnb7OsysmLH656zVEwndQK4m3ypiwnUeMxED11bSVlSG1/kREke/eGGFH2
VgTAVej8VYn5aTk8p5dMLnhGexzus5R2PIE9/3TxauxEYl7dmBojfpWtTWez
+17Bchau7OLO6izJic0xZhPe4OnrLjaKdWvSuo6jAQdNL00sSo+iIpN5f1uj
hI0nr/w7m1SGOPLVoTMga4xz3iIemEenuaVpCkErsVaDybAGcZFNhxhwKov5
1uyKs19Wu0C++PxlDkvRdy92ilZIYjuX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZOWjS4QxUk18Dtaol+DAPqwFkwD8Nvoe2I+HgzQ22FHcVnzkm11TIIy4QtT8
wm4pGIYJOji2ZcMMvnU+UyabnEilOYugKi0ljtoOCAM4zR6WtIzAA/QKkTz6
ppXdAAMat5XHI6aGA5F3Id0jj1gykgZUv9pcpWJtRmpLR9+d3RQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B9F4laPLibBmJntEdquXbi1hddbU2KobL53wbSm3lNZ39tSOPQbXR6eSvF6O
J2Qm/VwTrBBLn5JwoGxxLA758lDvwuLis+1r3V8GD6xuu+3IWtLXfPKmU4aV
HNpMJEf3Yytrn6OymiSMqoNiByzZYTjHL2BDRTBInm5JCMrBGzk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9024)
`pragma protect data_block
vU24RnRndUAYDE1o29srjCp5uKNsK/1yRGo0FC+0LJumDQRZpa3U242Z7XcE
Ozvt/ZRbwd2zJDfgkTVgmtB+W3BKx+l+21IKOtvfdhR8szaNlxM4DFJKTtW7
JH/kR91JrgBJpeEXvLmedNn2emHiURiH4an39PpNGtmr6j0Xc1AqX+0HoG4p
VnZooFlbV3D5yJfCg7Q2TMxUglj5RYKbXnMNXuGQxFHTtzLyZ3JeweDT5g5m
uLf/w9AU6s6zD5hyGFfrV/DPjvlGL1sOhwIjfTIunR3hVJaAgKeXbvCACPYa
S4av8/Mvk/xhD/XKXd0ddw7x2smAAhxbX22NwjVNMoCmpmdSyDmVUaeNSCRg
ZB10FE/yjL1m4Dv0/ePFbHNDT8BLyZjPB5ZLV50s+mAiRYhZjRVJv67OUjTD
Rx6ADxBE0mn2Ebag0bKDgEfSOYCaXqYuVIMBrhOuub9iUHHi3bcCklalzqiG
dl9W/ibuvzjAmKMmtS8r21+UmziN7B2pYKbSeH5UYVeOX8gvsKrb8ZkvvV3e
nnjjsrI5I7kj+6t97UMpEAEQkiTTS2hODQFXXSZ/87EpmiQsJL93TkvLU1eB
hCJPRuUEqsWB0IOY3U8A6Td29fZYF5JKLMS9aN3txGhdMIB90elaPgytsSkQ
9DuiH2ROFV4uMtyYCdG2FSFJo9KoHJ2BS5Wv++RM7N2y2XvpLwXwGiUFAYxp
zMj6uijDW/QXkPeGGgXSvogawR7rkYHVsCHXym5NzqGXtUrkGKwsrE5Fu6pu
DWHB3/sAKe05IhOMneLHL9Nsoo/1wvMxwhjMK8wpnty18cKISs+NJZXUSQ4m
PtOywskyDKkEsg2ZmrTZKZnfKGIwdPdqEI1Z6TBbCfeqpFSgcxFRbWroB4oJ
4f58WPuN/2uDhokfiLI8WjB2CJmtsmIl4mZMRJlV/1VPN30sJR0V22HRENou
GIOXkho6+rDkbEVUsyd9IuRVyqIzsfwghV5TcnwxODyW33hsQb/GiODsnEh9
S3Q6+nkE9ytOnpdYDaFwQBauUzxrkEIhM1RY0A1Xuar83XvPnj0b5bB+QuxW
wYKO3LOwvkuVHJafYPDd5Wp4SltlbvrWFQTD1X3n159R4kmVNRbfb/8nkjmr
TPrZpLg7m8ohP+fOY4cN6/ynCH8OeI1pCKtGkX8oE0bFLwK8glFRFw1tPJkI
bIMnWWe4zCMNWw4X2rIsYBiftQspTZW3peJzxb2eBzh0hF5dzt6qWwpjvBRx
ZOjrQlmjLCE16Xk9lytXxj01SDl8Zr5dJCezesZ3RL7PzFG/U6ODd0EvECmS
i5ZgQd5riHQ/zgJXinCLsL0gMks5sV73PHD1CMrAxbT+XahhGlzea5IdRP5F
gf5aRn0V1iDMPTYZFgHef7MCG0zMh92Yhf0qDdGhKvAgz2CvDufx0hMOvdo/
1Qdxv0Pf0bMm+KfBE6NnmQimb1ui7k675oFlyaAAGkjRkL8LwzJttXJXR9Wa
GRSxJ9LMPee3WZiSE3Sankl0CnzXNoDeGn/f++AXhVbyA+PgZFg/orIWy26s
N6MwDf3nf9VGqK2Zyd2RApZpyK5rm0oBxwQFPm7+I/9b+hfni0GVipefsFZi
1AUpHeNbPFZu+bWlFHWZBhLmmm40kJadju8lD2bJZt+4wU0jpBae9iCfeOPw
0qhdXrLoN+Fyy1yAH3/7a+3UEAo20DSBpKNnb0Cf7bNO+QbXqfjqPwyNn/wb
C6r8648SYeqF3RH+LjBJC3sEqeAdDLh3ebiZMNC/ckgqfyTdAoxJwZpwHxoS
hfZN1B29B2Oe/fAnK3WjDtLKt1Xlxn1cJeYgFeorKcMgEaVqjOgp+Q03gxQA
D27KgQHQ49QIS6284WBJ4go1XDIAziVrkWM2fU6Giz84wlc9YBUoRbqnNOuh
TzZ7bzMgRmThklaMMiL4kY2uUn8o0BnxQRtoPEYIUKfFjW7t/OOU5llI8BgP
QEa860JLdRpuGR8owng19H92j2CC7R0RIf1WxGesWZYJlwBVeEUKiK9iJv+R
JLXdTs7H5BTrTbEBefHrEP0gJi4eP/uzjEAjGD1CIepF7LBzZLmp/irnPjRM
lZivqcUIxFCphlzBt0h72uQ7HopQkwOk0N0eY8xSzdoUEFAD4Ae8rOI4j7TG
eZS9n/VeiNygfVqf2lK+gxTzlB4zb6445o613LFRL9B8nukQIwQcH8a2TFRv
qV8P4E2hCcr46IBoLTXXXOb6LrM+9qHL18I9Bb359Pl83H6diqF/d7SRj5t+
18pfzVebH+JWnAOSMoLuVScnyhO2nvswm7lJQcoYhBAhVVyZm/Xj6wdpVUfI
gArPlAH1Ui6i5RnDLgHqnMC8J3TGEcR3hdC7LSBUvhA+8DWBEqQ0ZAX1Jd+W
+xR11V6eN1YyUS19ccLqS6m1NUHDUrNOlZSF13OQpJX5fpcrs2rWk/086f0t
cCSyGMFOvRhx9JOk4Zl/+WeKpvtp6WpVVMj+AR/uUJl+rx4c6Lls12X8Et1l
AErkF2IDXTcfHdO7P5CG7yUWskhVHCSJh3NZKlZphlQyaMqq06+10dQBIx/z
axjLqjBCUeK5ZAgS7HbZ0oNopyOy3dbSxpzkO/cFLsdTh5I6pX0eg+1xVn4E
pIlgCVRAK7olZNEHIu3FaTRncQEQGWqGbg4jSDalLVFjDjdZINqOhRf9yQFK
FSqQo7LSEh58eJdHv1A4vL774YFSV0NzSAowCt5XjHg3S/CzcoljacKYvC7v
KGlnVE/Cqa8KDT1MAwAdJrNi2iZvF7+XNlIbwX8gAg6IF4YIulnXHb33jsfX
cuPdHefAjp5CrkqRyk+1rkNvIfO2QjClXaifChrvUa4HyTGXwMq1OrX3NNh0
C8JcZEglrrct3/JkynDHMsN1KmQ34Ukh4k2i5elXpG3slNFuZETzSgCtH56Y
3KyrIMAaBnjozuv0D7/9evNV8E55jgOjeow7A5WtKz56DTwwwBaIesJhvEcG
YCTZX5VC0CugFOGmzpzgfCnTwurRErWrc7zwsZz30whEn0egYKbScSIHcl/l
MbuRr583L7FEc0507flMqRFQC9rVQ0+tuh7LIjMtHnZOo6IltfCVVKKon+jn
QpsZ4a2flsPLUjNCgsnoLfHfWUr9ev2ypBMRglkZmT4C/lQxoCZeIJ9yPsli
dPpjQZ1Xu6wwehplqkyglboEsshCce+ORAKWSsdjJ0SDFMWU7FCGrk+oralG
SsxhJ92TwTC83UNHfYJZxMjz49R5aloJ3/dZZAL/rQwLL2VVN7TfL1GJ3lGl
orPufcGI+oKHKdV2s6efkLnalGSHOf8KA+OXp04dM8YIqbzyHLb3M3ynAgvC
cDak5kMvM4dDp7Q8PzOIjRxghWWqBwliZYhA6Few8D0Fc+qRRnPcl2WUXeu/
/cp/op2oLiAzPWkJDNe1CoZY194jwkiCaUXe24yvrcS4NzY3pPQy9P2pjUC0
cNxpX5EbVvojokotL/8NNl6V063bspUuAwFqsmbUToF6/LTEfK37kdweWHcL
XVqM5XiOah1fJx/pBvfPTdA4LEvLqCib+3XGJskFqkyWBiFfliZ0q2ho/aKG
WV8Zw+52eZLUFydej7NJo0CzHfemSZoci4MQizAI3cDtDi3mOsQMh3m2YY9w
9mvCDFC4z2eaiotf22xTefYdbqmZRivQa/7vINEQ86EwQ0mTDGjRy6Envd8B
T2eGVX4pLm8rrkkLGerHKqmnjlejZz4baf0pWgugp3ixN/3GBolLSpev5BUc
NFT78WZIL0W1WlxTnRZFI/MxAJ1vlMarJXy/2yugC4f1zmxJnufV1gXZttWw
SqHc3eCw5usW2SWr6+hhABbjiB4yfBJrqCAhMhx/JbNB2okGMpLwJg+moqij
9tP1zUjZX0XJFVO7T2xqvJz91D1WYfMhMJXkG0U1yuDIUR3PLa635mZ8peXS
qhRwWZhYmq9FLG2MMTCjEU9KIObhbguVV0XlThuJZUtRK251mmvKXnyhKJFX
cbUeSRll9U1vLz4L9glTQjhrsXOpwOjvy0gu6Yci8vs4DT99ES0W8Sk083su
ww0Th6q9fsCtM8vrhay/7aQqDa9PyJHKJsKb3hmXBOQNyF37TO9tNUyWIzrp
SLmZ2R5jhKGlnw1REWQ1GwASJ6ojueilMxkRDrNt8hcGJ44Zo/mPxo3ouyXM
XRy3y+fiBqZTYx63bHi8MQN748sewNx/QZsg3f+X97iZ7S55u6jwtfT6wT+K
dEUxy4zA1qgpqtI5rIwmo7Uee0c2ylnJufIwkYQ6WVMfGlfjalqBN+D01C/n
Tk8ZSwdOwP6Hnnx/DoQw7okOtGY8i5ow4KQ8Tz5jaJ23ojyl0Eo+wPMa98xB
VvU6rDTTFtTGXxUGM2eebffWSOm4007vjQ7jTuHE+5qr3xl9G//7L4uGz+JJ
1Dhw/fb0IkHnDO1Ibtj7JlkeOmbohkrohCIASDP/I1U+WslJnzKY9NMCzgC5
Sm3rVDYBDFWzNpt7IpZwLuUSYkI2W34FM3JWERxYYOxSro3DBIspaifdSgM5
fsgmwWCuZtEnlNgoVdjGqaQqRgl7AYPIcBdxbPyZiufYFCflxIWdCFdIyB5L
aENHtcZHlKiKA81FsTzrOTqbwbYZTH6xDlJm2gk+lGNvJOTidG3aL/4wh1oD
LUWxponvTUg+kJCiTmmcibzjc+T7SmLRKBMVh5yqvKfc9OnT8Z9DbqFehyUR
MbVY1bOD4ROKs3kxXkqAQWa+bAwc2axNa1QV0aTrpRCPDVTBg0XPic23xxN1
xmJkfKb1zINlsTeg4J/W/yIu78Z2ajE07vmEGu+mvCJdfnYMQrdnRZbJ+1Ts
G0ect1rB2iBOs/eXgLiYhhlMonP3i+bSou5cL1glC6p2BXqeFG6AVb3LoDdw
VNQVljUNhnWYUqu5dHXampb8FO9bwvPH5oMoA0YTUMvKlI+0y6meZYcskUNc
CMn/ew8hdhUV3F3xCGCsd+61kj0uMnjKlg138U3jinLuS7uMrrnrBQzT2DKL
azReAiP4eqpSzSpBhCrHFsePH36ld1GAa9jDbbEe2cW/s16NiqQ/03OohlcH
KADI7AGAYyb+e7kYvwWZgUTcOArqmn/mOEaLCyfURn48r8IJ4FK3njcSyVJT
A27g6V0ofDE6IE1SgpRaw1ap/igJWesxsqUU8iERoOTZS/bRUseRKXiAqfRr
orUzzHLCcPk0lU0aEKnRDXOlNRDJmFV8/A0C7O5HYdeOj4lT/x28mKkl14XH
FNl6bZUu8cV2Mpw43z0uorjwb3TmDGume+pRnCzOwuQu/w3vrS5ucRl4UdZr
xu+z9ko0fId4GAoVwScHaiGS+MLE4imjhRF3AoYg6W/RhvAXjWhnwcDjLcHA
w2RXMKFAqdj2ga2xonF8DlcGRlHF9cTKVIbrP34YZNjYDcIZEGve66LS0LRg
vccPmXdIb6E0LyT8jgOW7EhGKh9SjP1XpTAo++/uyZodw1kM6H3bYhXFtpxg
jA/W5t44IKIrzfAfWWExJUI0cg3DsxQNifdmwhriB8576MqIz0zOSAV/fZla
gkOSffcItrijskI+VHk88hNPB5jcThDdI9No7H7VlrjTu37GJl1TPoT9Pd62
R2mauCrvwr1a7ukMmOE28/6W61Nf4LYwuhfMzaNTQSlbKGHM0wkrPjqhyFHa
JXAYWyWbFGKfTynGAvE5JpfDarYvkOn3U6RqRp9lZnP/k8WOhVSMU1dkmm77
Jkq0pL3CMzr0aWOp0zqb7Pl1Pmi8HD1a8Px4/xXrdwLyoXcRCsJPhJ4qVdSj
0PWEIbN9CQNcfmnTIbYtDs6x/y0AXTb1Vs7FJAIrsQuGx3obF5x2h0FhMpfZ
XAjilUtgb9lXQaLb2Xr44B4T1KQsfyGnrjpP0rnE4HduS6W6GCaqMkDcgQDo
JvWmaqiKnP7TFEQpsb4X1JviLxCEjUB7eGmbUbQNFakK9KQ/dhfs3p7V50qr
+kDj1yk5NYJZYh9v2+6I7rfMHE1sZoCsmXyT5eDzzMpo6r3ClxAtqQlbxme4
r6iHN7RKUJ+ZqN9szl7bJbnm/pIuRFPSOR5ywuidC2Txt6VIZguE4J1Yhqpq
teKto70RfgBH/IxyxwvYdPfuay+TT3K7uqHeK6i+BK+jmYOw3mSCA2hy3X6e
gsNdkWpVjRgr+JBUVhe/MymGd0fpPm46AVRikCFAIT9d7oe3/yNBzETtN6oc
f8K2Up+R1r/baVR2yBGSAin52syGmM0fOmbk9crjv6LyS2w9BSdrQWN7Fvxv
dhqA5AhWdH+lZ6achd+jbMd6To8atJEEjGtb00nVRzQ8bKSncTAg1GM786gd
n4TSAxAOF7k969HJ489Lsa6l1tCzy39tTVwhAwSrh9O+ddd/zLu+DbIhmUa6
NzESEgV7EB9HjD5aEoPZjGSzeaHaOcYcNDSITkdVV/grhGHxEFN8JJTS1Wet
oZu2jyKElsek6nbsHsJQFKlp1NCprElFLxg5FVBRmtXqPZDYjjNHuIv5wPVU
sHeQc3TytaDcChHFBxy4bKZ0nWb/l5K9icYU7+lBxlcbx3DzJKUzsFSwdlM+
+GfkbpHvK8tBrMCKKEMKYs6vlLMNabrp4/Qz+Xf9Og+x7Vchac0bFhOy66Q2
sC3n5z7U/NkrIVc4qExcAih+Z/HjAy5XKPC09NIMpCCi+9wULAqntpkDFjV3
wCZD+40Fb7VWFIjSU8HqzedHSekiRiAwjdpCYHOrtuhv3KAvVhwN+NCSZj+W
j4+L1kF1g9WValktoXr3ldQ2ZekoHsWnF7vkjQu1v8dbeYo6/abmlBVxgQMB
Vpvd/RfLtXEU3NQ9ZTwTYeYj34dFdP7uiVg1UsJEVKhVe4iWAmE6CnzlKRy1
7T/J+CSNw/IakqWTTHWCJDeKxhGKiVEl+yjnC00y5CKVsoyY1arnsYYT5nNK
GnA8ScX9NCiquKWELjuvhMeT2tbwZJEO2P3rbrzd4CQwUFFd5DL8Vwaz2WrM
+4cEwxIkBeDAphBPpx18bigEMJyQxSkK0eoF/8Co0PAbJqgAQc7AWTY5lEbs
cdnBdQp3/AX52HSvjCY467SCrYDwcj+yu3NiZ149ryx4/TEm8lHG3Pmc7mfn
/KN+1XAX3/1sYU1qhcXpSx5zJzwdwoTw+hPhuaW8/sKg8UYIX4KlWVbZwRXI
M2EM5ni5t8x9LwfAE2cT0/G9QkysB3hhLvwkosXOwPMIHHYHOfocafIafTjI
T+k4JyIrOOhQiCpyDF+5NkXkwrlSw+SOxas0FbL8YAzocG63Ydp/svAgBgVO
sJFqP8xk5rBqmqBM4BQ6jtDuWLrUwZXDJudbAoyy99LUMvK3JRBk05CKl1zD
lo052L8TfldS1HT1VYXBwhiFFLBn/MvwqZYi4FmoLo7yaF9r/6o7if1ENTqS
MEMa/70aiR75p5A/tLRsH50JeKERzQvcfO+8N43zYcDgVj4ofwUZMo1F5Qrv
KLcpGxDgsI1RU0DkPoNiq0jmvDE3ZBUKymoGlzD515WP5wMni+7bdt2oIk5A
H/MlgvI1AyuIFqFqLWDwDl74MpDa1fThHoKCLI6ru2iD9l3gKrFtnkx9KKdx
JuXdluLOFxx/g+6Nhn/l7Gi2WS+zEPCrf9Is+G/QMPyNs+rOYmT3B/dNpw6O
ZegyV2o3cuvwAlTYU28EKMsJ7Wlu0dGBBSnGy9BrPyG70/iV1evjQ8y2v77M
o8Pxsy0fu41aGNPQdaIX9eQyo6IsC5Ghm3BLENTpgQx842264vfeUy4I7+xP
nXDo8ROEpnf85pF0KlrHTwmTwyOnTmXZB8njjlps9RXEafLnlhBk7amXo3jy
mlelXVnf/nPR2YJBMBzcfuLNx9zwDuXSrxmewn0Qt6EIVCMOSz2x4n5trVA+
/i69vpkIgXqhsotl8kJC4Ehxh/fHaX3rK67waLnQudhcWeBomCcxfnuGm3DL
UlnUsSAwv1G3BV7CO/QotzMOYi2eLuXWzH2Ot6rm3VQY6aqlCYJzOHGA+jJg
ZekHfyztis7J/PsBJWkLYxyLngISFSIDTJnfR6zPKDyc2F2BXzCopZ46r5eS
9a3bGnpcOtxTLynaLHtdiMa/pMRIaStYiPkzMxzkTZIGxmrEIzzLE1XEXVZM
hE67B4lnmbyUHz6ti062cs1SplD0GOKnZbHyhYMGqrhDb+7sPC66uWgYScM5
avl0wOr2ju+FNta78qgCBZpQy7YldT5AaTO+w8p/mpPFngWIUiwrGwfY2aE4
b1jMrzvUHKKSF/E3WGQVQvP1zYRg6rHrbbD+xQb7gDpoYrQNqpiDjl6stIvZ
e/y3BDNhPeJL/dZDbEQmEyA6ts59OVxnZgd500ldNegqw51lhd5PIIHY8ydk
R4d8m26RDBpqHXgZZuWbLjEEHUlxLOlehxQCXX16ZZs7umsRQnUsSdJuwPCu
ybu3dkizoGL6/yGfl53KH38DNAesJF+2Ym7E2ep36T5MNrk+C8i+TaBFbPvr
ne1TwHB7yVeuVNP1z4/FV4+Z934uVBKLs9mY9zNbSrTiYw3Nqxn4qbO17NTm
yT/CGgH8eu2BLz5gMrZWmd4+AoCNu7In9rKTedEarXInYpqQV8F2S6pbHq22
bb9uWwNHaCv+g/yGA+8ry94v45H7QGWYnVSkXdjIflvcFCivd7bzJTCPBtlZ
FJgHqJC82Lay/CVl9aKDL1eW6dkaaXkoO+bFM8rQW45QkWqqxxDYlqP7Wr6O
Cwwf1rwmkxekIDd5c1V+GAKNKvLsexikacyd7UkJrJEWC1Egx/gN5WxBMhUF
oqgaLA0d6i+5bTLy15gDwEXWdcfK4VxYP16A5wztM6yiu9T7avfqagArvqqN
YB4pBA//Ysv2sccjouUenASWx4I9vzLKICh8mnuhA6D74V+6WgP9YtasIqYd
Z5q4XVWF2PCYa7G2KDj/e5fnPI5hxVdLk7xCw2ld7lusOoewEO89PfNfxx78
qk/RwmQ0rVwrpn2BjokOqE5InP5detNOlAg5cf4rM4xt6UoL2h6yTZtp6RPw
LTLdPYYJkY16AlWaXOFyIIyTkeolyuiON0is1sJqjJSPSykdcAzBr+tCXQLk
pqkcZ0vGvOZ+muKhvufOylJxueRIdFzbHVxi96ufyqLmZ1e/NuUi770VfKOc
H6Z+3IKSu/HsQPOe4K0FvH8uMuyGZhI11NF4v4iWQ1MljNn0odmzMUkfEL6Q
mV57NZYNM0X2We9Rhp7G8oEm8ZWWO2mgoygx9rOQgDbsUyDNgt5JC3OifVZC
idM717NFuDMYfI6Xjxt7t71y+gyGlp0Fnr8RnhtIMj46c9OYPzSeCbCnQfHO
2c0tWBmGF7Ew7xiaXHF1Skn4biujMil/kBPBodHHwinQLE0OjdFcz+sLAyZK
fj4LmXXq+VLrI8RCu9KpKkL1HPaX6ajJZbLYRoX9LT4dFp4cDKWEbj1PQlpS
oubUyU+MvvotqEJ9ml5gklzBVNy77x2IepwvLqX2mEbWVql64i2lgaxmZF/z
WkriQx1lVrcgL/cd4rAPWwxnr1G7qw+Pmh8yloP6TiP5jtlIvzXr9EGo7HqN
z5DmZl0/iHXhcpRqy9tjcDxXyTqGYO9J7mhT71S9GEv7/sSTdKc+PSQ8d8xB
Phn9/bMY8u8f2Sr6wFkcwVXEujHek2qMeJo6cffW1A1Iq4h9TiCXxFbP0cPL
uBbGVXnQrAAPz1rvDsvzilx96SOXyQIR5SsfSqwuZNHGVtGYMuCWBIb3GLAo
HZ33rRC4x0nXuoeNif7mDpcS5kKUrwOPb7oZ+9N0BhawFEppTTh04gG2kSE/
ToyfwvK6HlitGDiO+PB4HS3LICy9btRhjaEsP9/hqboSsnOq/qPKkXcIoC+U
+NbCXhuMY+yf1rClLR1vf3EkbcFhCwvTfaTJOTb9HdQ6oRUICt136jL3E+rV
kKWcaIoJMBRLixhVtFDuGhHMvDiYIgjpV0VeC96BwWrcpjTuXsGgYqhqzW3K
/6sfc16YvWSydVx/DSvH77uUWpl8pwtcFYSDv7fPrI0k8L6sWYj8sbN0VbsF
4DymsU6SqFVB2xuet5/MIouxAt21WFUrnWvwpePFMXYVI+LjaNvxX+NKRffA
11BffCLzu+jaCIwfq6AC1wsJSuLmxDyqYs93CwPqX7w97a2UwsW8HrUXpoV0
ncs9JAHXCmJvCIcriDQR4am/8fov7mFZeoY/Sd3glNmJ8t+9cEw5snv8POsg
irac7D6GbyK7S/34y1WPOQMrvKtWrs16B8mZafYOSHD/Zh3H+c/ZyMNNo+dS
8rzyyzKMyypjwCCK6CylbpAxK/BbUQ6UlshRfxmNFCNnZeJZAsjbHQd5clVS
Csld0S8i2sq6SL30pYcMhNbE2Sq5uxjasF4UYIQzR64I/41OfdDPWwriiIew
kGudIWaFqEWSKuSIDm6S2Oy6JuHpGyGJcj4b7qmGSVWU0lmTALcL6Fm3rtht
1IEYtpjW5IM/PRmS1EXTdPJur6vb5oJ39Vmu/FZ5QIip/3onmYl8W2bbSldV
vWgPiXuJsKKSvoARSurW0I+cJwva581epqz2HPZst2/vLRRbDdNG22ZjuNQd
HTtSS5tv9orgcxfZqw5AuhCLhZCD4u8F06VNYjUBwPaS+4qx1E2Pt7xvbYJh
LFY5unBkbasN1BuaAyFWaHpKwmxOxAiPfh0MepD3rfJnpEk3QvZsQTYae2xk
Ztt7zPvBbcWTp7P7PWgD3eG+/MvUYjm6l5hvS6miLU1Gqt8aqvfc804CCVdy
pCWRoLK+RoEcChZjLTuh+UXp1ts8RvJRAatZey71xFaGV8ZzQ8jEqvNvGrCh
HQFrhuPXTf/b6VrJroTVinBZYSuMV/WsSc6PJNgVnpyPDutRGO8WD2Pzdgpj
Bb0y57dOoMXFgQEpfEZpibP56prqHcGY1AhSqGIw+VRryixbukPofdI4Fzpf
kzqM19BFXr80TQC1dpX2eUdgQ1RwgSPx/r3TI7+m11ZNXlI1iIlVe/7uNW5Z
FbJQk0zEgHppA0Md9+XgyUqbT7iGEuq8+kXshkOq2Ne9kQUVreigL0pWR16F
nGPmyIqxGnTZwGw5YZ5/iLrFXH5qz3fOdDAoMaYXwKO1GNEztAQmbtLQeiJp
7bJWp4wrkkwHyUpsxNfwQBvTYlSUZJdguGxum7KaU/pwGiMOU1JaynnxZ7Q4
jFQp3Rl3LFqmqkt5FnyhCJLMblvvxD3D3SqIdi3SKTamJ9Bnqjh/68bpeIbW
aIjv4nG1n1IpckfVUK3oM9/knpUMlzEZZ+K97Snmbh4laVipr4pWI8pWOFle
HwDZ+VZdWVtA0I9VYWp6S8zcaHB7v/HanmLXtOPxcTXJwoSPdRQ+pegx9ruq
QlcGOcPDKUMdYtOXlm46TRohvQXrdoanjBoXiwKKt1PC1L2x4jJDrKUg0EUb
GnaA4bGbobMMS/OLhqINkHAKuSN7TDekn9i4Deuho/mbg+Tr7My2eqqB0Rd/
6HBJtzA5jjjE3GtyUvdLmsFP1jEKNZ2H5fCfv+oQ0doX6C+ln/pbZPLmvJvX
JOWK0IvJSKdwxwRA5UmVMXxnSx6L1+HngQxsd83pGOSzNZsXa4fVZ7wOOgfo
mEts3y5w257tVmmRLiq3TTs1Anuc3w6lKdDtx8WI+O39nHok7/sZeyunqPSX
fszxg8V6OtCR713R0VPQFagDHnnTWcl0c4/n6kiQAEDtgBZ4cIfjmu281+7m
MZTEVCjGy6flSdinCFRt5h7wyz1ENez3goNRFv+M+r5d0OkYwApiU/fgjUMk
pYXnYvaMdYeY4jp1flrz3JKd7R+MN5EkAP6UByPlZvMRbkENBr9jQU660Im8
TKv4Tx8d4yxOie+r2omjPNeTpWgJPCnKRi+RwGF17U1eoPKw5ZSmF9k4ELY4
3HGlXlwWCdif4FeU+NW49fFXBBgEXTnEknHB6HV15aJTho8xhjQOzLqFaEBg
uFIZmx3687dFPu++usvoj4xyAfoBmxBw

`pragma protect end_protected
