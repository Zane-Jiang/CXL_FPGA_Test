// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
rq/5B8y4KVHpIKqV2QUzaSFGGpHu0+m+Ke2SliwZL2rwTVy6MDdWg7ki++LADu58
6/E+8MjSbSJG2Ljkfi4XNiDYTZjiuvlp7/4VeiIegS9M4ECACUpf0pplvjntZHXo
pyN3QLM7YYzVrlOP16OEldBD/xwXo0GM0oeoXYQhuTQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 74400 )
`pragma protect data_block
j19yd2fvJ3d922Sv4r8/5YEZiXNUqC6aZyEQXuP8faBIBzIT85FkRj/MI+176ffG
RQdyqdmnCRDNUvDt8CZOMcbFoeKJwIJoP5+OZ9kZufs8N2FDsRVhIXAKyPryrkZM
HNhZ4p3u8pTNDi+DXy+5scWvAy9JmVnQLf5QzZu9yov3rvbKaj3FLM06MIov4yl1
ONfMbnHsHgyWmwj7Q+Aj3j7DvxNP6V2nBS+sN28RRECXvEhKZfIQOKd4vVln5KXn
eQG2hXJxmWXarKVutdNREoNW3kLonMwiLDbPtmq3OzmehvkQwDEj2/iM1JVIXu5k
9P02W6V1LVjzW7otL3u5ntbjWct2SeCMffVQ/wR8xWHoAaCINAipU8nXAu7FhvDH
LCcYFk7b7BkfJa6TeihbOGMZtlpZhgsapBvDOJLQQLAM4uhUPbHXQpaz0Xq2RN41
KABkg0S1uxfEamQ+Ijq68yky3X/mXZIsSRZWdl6CPXdO/Eev+MX/t1Pwy2+ItbSu
n5fzJbV5XP3/d98oPfhQLXSDpOdFmK+b7YOtQzkXiQvRk1W66SqWUFK3btIm5MuB
LlT3hU3QWGStDO40QgPTR7vC2AG7F2NfBzwGnlbpSr6uxPrG9fnPxW45BLkU76Dm
ojV14Y8w91bd2aQQLG78cJXJtlX4UAzIgBccVOwPBYsGRmMnbXvAyLzc+2Rr4Gpl
0zUIuqwn5Cvq8Wvb5Onif3Ky0usYddHhvx/gXcHRM4sQP+Fwzv5EsgwL7WiD8w8D
wUGmr2ZTmKJbz8M/jyDggRXEwFXDcSOtDO0HclPyGsrr90p5wQLufr9UQ4jwY0Po
nR+W0bRp8BSGHq+XPxR+9ThYj/ze9moR8NkOU2roW0ZZhJpISqkbsSQvUdYOMwhz
1z7r3AxHSf4MMOCJVubTdhWhnScYbdAI4/E3FRBl7EkCreo6vgp/rhWLsbsxeDHu
6X72rg8ZArrLSC9Ci1k3fOTRe/PtB0nxysxmj0/ML10nLad2JnKn7ZfZi8+C8h7k
Dl+aBfzFPROXWPJTJ+DUCNj9gk68K1CELQhwxXE54ydUjEERpdZe5BpuXA1BtNmU
JhooGf8Ul52qUIMZYlsMDccE2SGGPdtGdMDujRQKm2/SSJUkyIDhMLMFDleSTjPF
A1ZGAYGHI9FmhWUp0YQko+rjnz+YlmLE310eF7B0R5C/iQdnkq4tAsEE2brqlWrn
SWNMuOY7+kjC73LasTzPUSsbJVBCc8MfABzWcNtPst8xBsDca+M4k/3gQVQLobdG
OddohUPQhqHsI0osPhfHZGBV0PD8qf9FBcVaai3ip7xS2skBKXH8S/z3ubdV1Xc4
j6rThPe6f78bDvYfhe/P0Hk8ugtB8Xr17+a+goyrd0Psx/7g0BNlxkD1M/Ubm6tn
aUbHOsgYMEwzWYfEIcCK6yy7ph3guDGQUjFj6TkVyYHIj9Lp3XP1/JNHO1n2v01G
m4dIvKcAMPP2lur9uF+tmSJcDRA05w8YPqdFc606p85jLxVPmc0IzwQ55BOROZr4
XAMOQWz07yxlLpHBWic+6S+7IWGGFz7j5M1MQnsEdWZX9TNNR98W+avR589QuaDu
WnPuBQg7bh9PcAmFldrPbaC9Ct8vhz0EHVqBRpUOUGn+JmLD/cFmyitZ9UVmTM5w
aXVdydTJ8NNHYbIxhATPnjbj6nHck5wUPfeSk2E3tq6xIqqeDGNNeRNzTHkElYbz
QoJWtanqeAq4QsR6iL5RZpns1yrObMVPMdljEE+DWK5ZhcLgEe5zOMKCTiEyRkKW
Vc5fj4PJ1Db1BlXmIdZu3ohCEIzk+s18GJIrJc8GzENBP9AfqKMa0BCQ33W+tomX
2q27io/PZguNPcQj2kDs2TCf6gMvKKp5zeh8AL1FUkTsV4F+XQk385n33N4lcgAN
8wbsDEEpFRhklMgDPohFSjZaGdCZXAHuY96kplitEOGo0+agFSxHCj1TBTu1LJdM
VtNe+FXmNhb0QHduBNTpmwxITExrJGKcAPXgbq/Kzoi5AmHbvvrVuK9KgLpXhS3N
sDPuKggnRZ/v7LbHvmkYcHmZo++vRN5pbeTQmeEiEHMsLbeF0IqfxxjQovyfmxnf
PhKjNVu8LEslRDbEmJ680clkbJ3AtdHVdSwSKhkfVyUedhok+MPXqEX/wM4UTMyO
tloJTxHWM37ddNp0SPU2gmgSQFr575vQ3bDI4MJCy1E/1SjWfUVzHDYfP/K5FO+B
A4if7gZI21ddi1bmw/73C6gp0FNyQDXMX69tGTDkDahbzMyImkE+EgFY1qNgI03i
JYEjsybtoWu2KfW5oFj8hBMlJiotvBYrbGrt3yP52TGr6rRwiQAqCNYxP5mZh5r4
l/yKDW36mEbctdppZjaX2+YYsLu3GLlnebFPHZiH8+SnfrSMe8zKljuUEozi38Y1
Vick17yKvD2IoYgQiIXmGI7fmNJxCI0YUsB0ka9FfcXDqd8nTo9e5V35i2NQuQNW
aA6+ijTFNB5pVlnvFjKQStaMM9WwVseoJlGCpYylrgszYQdqkVj9GU/ljaIYeHWj
jkEAVWakAJNJeiRqx49cmHwLdKjO2UKOEWMm4K8TxO2bSLogarsWyHrIpz5AhwjN
MkBEykMxBio5+HBFoyadVM065d67s5txuKWMkkdiRbsdAfHd+MCdS4PEvTqv1EpB
/+t6sVMlnyTLvkEKoUqEa2aBhHuJheshIwjYrT6LhEHGE1UWXLO4uF3+RLArixi+
g3pI0RRiKzge+JZ8yDtGxrdwSRvwFzJSBYWl38SmOdYoVy1aIsElvtwdP4mte+9Q
OOzQUOZnbl3BJ2CZsU+r/S7FFWoPB2y68079FOt6IdaIKVyRyeGifZzJ/bcMeMON
jEgU09s1ukqnx0jP6pj0mCKVm99E0xT5jt1C0VHHOxOnybsB65ElzJPKnhXfroM3
caIa9L6u/yIVmFfcDnZkxaQyI7IvkCWYWNwili2nMfDutcJ/9sVJpOM0QlRJB0Ce
AtnLetteQdlRVJlBsBLBqlvTTvQ+Vev9hTvVGdsCGQ5N46piS5J8/2h9XMF1k4EF
pNI8ySAjdnxqDvfbe/TEtUdkKvhvTtKnr15bpjzhOX/KrRzNGdy1Om+n81L9DYNQ
kyB44VhXcmLnUteUQ6APiF/9wOcjbJBc6jCDOxj8hVKUNq1BMyTQ+oMndmALH3FX
rNJGGL39el/W+7g3tRQ9t6OyWA4oo8GTEf6xVkWxYN40zn0oV1bpP6OQclTdAjme
RfvAPtRYu1+X6g5DPxk1Usf9sp2pDxczCNDNsWUlgrzyDMTN0Aa9IV1hzJm5JM7+
w7fqULOMD98AlOPocPKLrZIjeZESSXYsMYMV80pCRo1UurMjr/f9MLqx5I39W0Aa
SS0NAcEhc3AsRlzxtMYZlUoDuAYCghyi5blHrnAidK6AZjmNvXyLL01bE5+IhG8G
kzdbLtZjKzFyx0Mvam3pozN+20HidtktvH4CatnCgc32KJ9epttcIuR644WYjgqM
68pjl6pVIzHD81994kv4CA0yjal4v1KdC0c6/tgOaZOitVSEXy7qlsItUhGhMdQ0
RwPPklmQxO4QHnlDrFnSu21flrO34na6ckVWAnHwUOcSYe4EiXX4OINZmbxIRMrm
xgc4mEaGFxmFWetuRZcNSSGmB8Lbm1tmLRvIhryqHz/Wq6kwB2egc50Hr2fkGpMC
TmuCs5QAQogTU3DUGLaTwTiN3eNmxQdhtBOfzEgvHeVkxoGJiZ4awkSwENHY/xwi
ENYqeA2J18Rpwn2LVxptzAFPr49SEtPvovrmh30YB5TvF/u2CKWmtMW1DngIB4BJ
otz0WyIGdFitWYAZG3bxsl4vZOL6DNr0DFXm8umOS6ccyrysT6elgt+kqD4PvnIr
mZpBLeonTS5Gmqw5KOmeW5GJG6kG02PAou7s+p2dZrLBg4qgvb0/Nx2UKhnyP6Xf
K8aI9RUjlyY2QCVh0dmy2GwwV1INKBF8qyQxd7TBF77H57GBSCEEN6UovIuAR9rt
yo97RNzDFriN6fN7IGjvJOJBKL8rRm3n9TSSfD6DyY4GcXopGW0lLf79LFqY367s
BBtVq6yor+3rDNe/qtP6FlqeRQd9oWizhjzdr41q2AlH0z5ZijkMCGgjfgVJYpBA
uhfjjTDApGyt27xPt1kPVXQ8It+ENzrE/Ib4SDkyzYhCnAYJxSeB6f5iIRJR+434
sW+NaSCQScjVKcqB1ltHTDb0tO9RnO8Bs9CWwpav/RkqC4u+RaN7a7VaZCmBg98C
sLqjIsdty3wS0UlU6+qK0VqhigI8FyGYq0bW1FiqtWZv7wN+bjUBj+Xnkor6NYhG
jSf5tCRpM42+L6BQxA+wcAatzZPOc++IyPpsLUmdUqt0Qae3rQXAJqeaOaI4+dJd
49sJeBq2cA52IelALXIuqwGvP2D4OnPvqzp0ecLGxwrSs2W/o/HoBTSgKAgRca0o
HFeYWDyAAYpWFlx+MoRFPMX1PLjKajKVfEwwo1LJHzvD7KtiQtwb1KtRkKUHm3tk
3GHGOLAleqUxMHZldYqdDbM2/C+KnTJsVXn/zV2uKSU3Euvs52lP79QhX4QJcC3+
2TPpt8WE7fBs70G3pf5szY02OGWTsD0jTyCC65z184DlTrbWb5CL0TdlfilbuLjo
2GUwXZSUgAOOWmBWn3o7AlxMx3lcxGlXmO2pcaLeZ0OH2/DE0xiGbBz+7IH7517G
h7wevSAOInDqyYF3FTfeoCuwgfHxZEjSgvrn8k54+r3RR/AAdzcF1onJyfAgg6wy
tOC7obTNfUr6kzeuqVJvgp3inMLmB0iKEg9o+pLjjCi7hb+ebH5A4Pyg4WJQikHP
bWG950fwczv7sWKFKbQ/K3fDnQrPnLI/z4ZX+5l/Vhfr1+X2sOG91QdLSFsxc0ew
xsVfvCdeMLxID3qQ7d9cth4tNBRlDvskepfup1D17BT8Jqq589uaJJ+c9QrQPoJD
+XiPX267X464XB4RLonDdPVTMbpBURtWYSjA61+fyyN54m1sNX8KdDav0YeIkkJm
Y+2iXLPGaijXISeG1+U9Uvl1uar1HLsQVKhh04RPdClDe2QtSV9PW5roxk/cjbxD
RvNFOe7k7yFdSDPTFP2mZeWKCbH/ENPclJeuwH3e6fm2MnGH/Fl9skHVxOv9V+rb
IdRHLnRXB+t8CmHf0T3pcJbkXzivYep4RjX4jUGwujSstW8byXPqLfBj1CFzpREF
A3/V7iRJ9oA20OrCRCYdGMepFYY8ZvqWG0ehbwpIlCDzBXMQwlLq5yIr35+Rs333
MbhvZjX44RIlDLJbceEVe7Apkx7HfSlrTi+v93NoQFfZw0Uh/eZEkDXzrPxTcGY6
cDj6kDdfPVnMmgo3TsRVJ8E1Y+QnttpXvSHTuSAyUpQ/hdzdpg6sZBxRp42ynrD0
zKNa/K+fa3ypAf1mMFG6fBgyMEPca9VPC6wLvHerVqQKGcTDDe7OrdZv7zOHyhRH
i3Ho3jjLs3o9B59ermkbmMsceJJjvKTAkqd7vRfyykpzFz/Rc2LOj+MGv4xuxj4r
WGILtLXCIpCQPMcAwUlKK3apDEVQNEzGb8UucyVsI3H+RywbAr7ksQmFp1CqhQfD
QJX+OUP8X42OTWIjz9Gxpvs3eAK0Nze7Oh2ddr8asyuQ4naCY2UALMrVcXlFf18X
VDV7tNEFe6wx8WiPNlsosNWGJJtlp27ZWS/2Rjh0Qcmd0QbR+EwEZuVOLSgg65Ks
Vn2WLOPhh7dgaxnhGORKLNeRs6zq6TLXM0MBNcF2ghjKd/AHKHhUznST5OaiKpZ7
6SdB+2qNeSUYSLjGTFZDlgu9Vjtg+q94DdalJlOC6osLDuW1EUjTobsX7CuNwKpJ
XrydcMqxQCguW/Z14Bs4r1f1dOFXsxFTigYOVgVd81TPMCZY0HZYf55qZKktcq5V
cORkEoMFz66b9znyRIEOsPIj/uBYDCbA6cyVf9Me/o7Hd5b/A4TQVFlFknY5Fonn
sNKCGRu5cxUANahgsHK1mSZcc58xejKmLQU/k5PYjbCacaeZaX05AbsHwhkRYbQv
s/+RatXqPCdzCbVfHWxYyZOdVBqtm3HIUHZ3HfW/69tlKWE5NeVCV1q7nx2mv4uS
w4F+rxhHJ98bIFYAl1CRJxxCgB/QF0HoeaxiR/+p9NMkPLThFRwwzd4y7P45s2ee
nRuvQwEQsxavgejQthmWMj8iZOuABOi6QwNhp/NWCjtrsVNn2tBkkglvPRPAX6TT
0/wBVhl1MMKjc0HAS2ePjIkxP8wSVcXeGY7dVAy41sOdAchqe+gCdfBJ68t8B52g
HBCkCnt38Upd1yogsuOjmU8qP9B+cDb4fjUKMTdB4qUFv/mG/wltqMhETKRo2zOn
WmJzTwYcxALO9Nt+4gDsg/JaZ3GesQ/Fj7wYBkOgA4xZzYfUVy+AxcoVQN9p+iEP
hGy/a5mdR1bR00502z6+l60v/3t3RG7E8d2KzvRPopJHIEC7KHlQJWQx4wPtBKys
X6xmBA6+/0Q/5VSw2BUpBufzWtXs1SYhxOocegTrw6Jb6hK2KDx8xseYSlMcFipO
MT2XGTO5pv7t77ZoeMOLfjMFHfQXtGN4jXyyli85YreAGLTQM1jqsTYsg9OnRlTL
jnEih7pQpzjPGdCsnrlNorPyGQcXaZZ0CEniZj4bJ5FcaEpqLdSMytMgg/0nHMQp
UaGxb+a6j0k0HIefatzpl5qJ1x/gXeQ5AnfblkMiVOlUcGBgsdPh8p6rrKTPnHyS
P4nyueYjngzN7Xb7S/65mXRKHQ7rLNpwG7+9ECBlk5GsCVr8nExLbXc/rU9IFHZE
PDkofDkAKanrK7hBZYZ2Eh0e2vQH/rvKuZsO67DbrXn4Bg24GOFsRqHMUenQwi6p
rnKffUBBoB0clV/zNYrPJuqifxxgSHJ8o53OM39170WJNJLtRJAhz7wP66yRMnOX
faDfy5+Dl7MK+ZBujKbH8Y183NpaInZ4BSwS4Rp+X4daliVrCGTI71ewHH6etWw9
uWBfjk/K9vMsXGRY4mJo4AgKiorqMNTJClhjOEzcuf/cWte1uOqY6N4mu0NMFXn/
+jL0P98GhwD5anTD+57Z93DWAQRwsD5YWy1TWZYzw2nOwqIW9p6pMF+pUjfvqDCs
J6qUjMrQJkzTaakBB2tmpPvz6cPZ4Xf2ccAXRZ0npqZNENCArbqVwpNHj/bkgHfV
EsNj1SvAxLI2Bfs3CRmYNJ5VRx+wgjVGrXoGXaBe0C3cvVr6CwTPzdskT2349Hzo
Kdz5hkihzkwkdSYvpcAqAfs6I5CjwfXYPV36WnYsaZt73oPm4PNKtRMGhazHNcbl
GVaG0Rstm+Abi3+9mlSHDO64AddxCI+ycLRC0hfrRDZaIrkQJVNot33ql2DqCDGF
9LKoDgDJeNB3zAVdByuM8cvoN6ZhFeZE7X9rFbrem6m2lNciFYM1tbgKUWZxht83
uUBd6adIvZkCJ+1U+Zg94+oPZ9rCBQbQlJATR1drBikQk6Xg8DdLdatE95k5bsMz
gCVuOGQ3odT9mOGejUGrzPFKvE9/Myc6MDdvs6J/VsFlVJnaMJJxzOlFdsuxx06t
mjXd/FKj2buMb6Wh0bAUgzePJrgpOHyBvvYkrHrXoDCpuHpQ1xb80eH1C6cE/8zz
nOW/IIdW1SSGJ34hiUCZrZ/OcJmvA4vNEThV++YH0nx2JJP4mJcn3HObcpH0fGbr
Y0ZJZQslZPrLRXG9oKt/rkSwDE17BM/T0uareN0YnU4djmZ5jTApsa1mpBSEBHLM
AKC7tYfsheHUBECW2hIsXX99HPjfhhoXXPerX6gLpZvy3Z5vPFCk+JCpkRSdXl73
79aCESrv5WoAvadB/pET3iJQwSHkxIkqJRAhnZlCoz9GRosuhz/Ptil1foJcsEBf
dn1+qefW34lH/bep0lOOWeJkRx7RPewX5yNrUMaeQJhW31Myeg4etwn8FTbowaFk
WIfk8LwRcJiP7ZNfHb1OSkk7YFN/IIlaPyQCZ7Hno9e4UJnHJ+Hsrc2Qr5Ou3i5z
siSG7k/Vx+PRRNd/VSEOUkJt0jJTm3TIWIULRKyFlstjIxvte6Ecb+lyn8tHfHaA
hyoUrxTnG+FJqnNBUx1zc7L0qkmnVzGQtbXnsNLl0XM0nUPsssXtpV8DhdOH6biz
oqE1tvIf20e2/QHMzwRMsxYrNZo3E0Xiltg7DxuQXuf6sMZXPBK7R4hSHNzYhX1Q
OOJM7Mn4zy5TqA9oY2nWC1nhrT2AhOpVZBF1pK3by8esswso0wu2g3Ay+kx7e2p1
mAKK1APtvJ//J6TXIL0I5Ga3MNA7zpTW5Muc0Au0UgKDgp53jh9KbhvbdCK/ynth
KR20rQlwKVW0PN/5gddY7VkVFsJTUb0LaEfo0bhoyjg9iRHJgcF3yNUJCK0Qlhm1
ThLy4BxL1ySFNGNpKjZMi/FyDeulYwsuxnC4KSwv2QukYG8D476whid/o0Z6UAd1
m82EQKgC0NZv5k1BsJzJ9n2YsqYBm6t/xzJSGGZIiCBgu7wFO8zBKS59/ZuvQUlF
m2FJHxvDLybJa1FRFiawmpYykpEzO7M3WPP7f4ifyI+B4uh9wXYXsDtwVhX5tf3G
1kx9sHe6Q+WUmQB7g7Cwp9RBaEt8Cn5fTCB2JB7pZHe9S/ibDA1reh1M+LEIrL+m
iQsNO0Z7OAWvP7eR/Zf1EJ+EZvzjzd+cCQ8vjzUwDxXdhMGfpYXbIr2WBhjr/Wlk
FbAniU+FFgsPNLD5a/xwmU4OuGskYGnWMI4UrYBwXBoxA8KqwzSJSTU0CmfC2L/6
sE2yMPen/C1y6kA2v+V2XtXBAg0WAxTf4KIaXYCsmoMecub87YgiBjbLlDGhdArv
z8tzJpAXQAKSZ+K31Dl8tJNp3xrQYQa5AWx0eRf80qwLDy1IJp/29hw/C6N2DbDS
8D0Em381Xj3t/atIfyFgK0EmrLVwvGo9pVxk0QM9NW2nnOulFN/52n6JoRxvEgWk
CqGzNsjvuD9WcSlO8qPBn0sIKuk3FLN04csKRq22wM0IRYOs+t58D23exdLHkXrD
xRKvoeYn4v17b2DNIxTvwpVLMikZ6o72rEs8aYsL20MwQNwZPait10qFroZzUzk6
Ny0MIpijrxc+x/B1jDiIffwO/J9GbiWuLxDJcSnEs+vr+8I++8zbdWpIzQ38p3SL
nY8q1Mh0Hlrv9ybrVoYT2SGQFm5qOlXarxWRijWTX/Zc4VSZ3UXDu3MFzBVTYQqs
XXAlSwBN7A++mI10V8FbsqOBA5h72QGycF8oemrTnMclmjQAddWE+kjZkb5YydiW
DkTxA418426XH6nu+3B83ATRAEJtjSf08Q2xdMrwvC3M29bfszOXZAMue/OSUELd
uD27/uZMu1w6dS0vuJNEHN6/xu49zIX8LWRMALaiCg7LWwyYbxS0zx7ljATj56m0
M9BmbXHVo6NRL9ko6VYwaWdkrcqdy1i91LbJApwlKKFXg2Bl+OBxJuG5HFEEfyBf
TPiLKkNGeQ7YwLQ6WEXpa54b83Hr2hbsFRaCE8PV0JYbjS4PHfQhBfXgRZ1xnBPa
hTaXwlHwRABI0AzHpBNLwqNp+GccVRck07w5EyHdmxGzTGS+yDEiATUn9hxrpx4x
Qu3WOqA2e5Qy/nulrZw31N6+kcpSxj1XgNLkhS+bjngaJB2ThqDDXe7k2fy70LhC
rwgFrfQaAbFAku2P6L42htBNGI6sPg6sVl3f0zWex7HwGoQVfj0e24Rfc/swXLlq
KqiayRE6Q3hiuOGnQpAeO1ZrJcZjqgEHO3V20HGEfq5IeTJVBfwpRI5h+zJtI5Rh
ln/wT48L39/nuuoAP9fuQENzKIOABq3lCJEqxba1H6c9YevHh+yrei0WQSORhdZq
BhcuSt8s9Zjo7/3+Wm+PIBqpSXgDvzbEkCIEsVviDvkJLlttBAyi0xdJNGrTZlkY
rPUzQ377NBe7pGnHH7T+E15WaGPuaWr9cQ7i92fv5E5peQZCMfbSqbE77GhsW3FV
78OwW4QffFYFar0uoLu6iWK2SYdsrqOecyNEZWbYeR03CfziymaZhevGp35cFCRV
/IZ/1o1tPeBJm5lRdQ9HZM1bw53NOs5SVTng07JOBbZ1/eZlU6rNLr0j1L40kXfo
ZolFJNC7FSs6/WHGQ5IUokG1L5j4V0Sd90tmLfmAkNbptUbeNZ9RliRjHd/ZZ15y
CLgTIOzJmBp7pMzjKxo+SVqRjcSSfmtRnxgYt1cOjj16CUbikMkkxyOyFbl48c3J
hRmTvUskNEzfPjUQsr+C+hDKHRVHdPTIcxNUuOh9kMC7hgpw7pimxAYXYz4wiCup
HRFMF0brUAV0imO+0D0AQFbgi+52tI0CI18xCy+AtX0eaRbWcxEjNyU3gYn+gkIC
NqhPiq4mEUiCShELCI/t5rvBRbssx9pNjxt0pwV5jR83ZmeelE4cGS6Z18/7TnwI
Ne4CG9AKgs+++cRv5ueQ9c74rL4BhmYXwb+xrx8KYbMfirlvkJiyCn3OUU/zVecj
vpcz4fOxalzA0G8FbfiA5Lr+J0K+W04EHOTj+/H25Z74YKsOKUFcDf4w0KnINNhk
FplSRSxKtRz6T37hEBRa36norv0v27d7x5ldlbu4GhweX6IOVyT09kkEfpsSqIaB
wXWGRaU3LDRIiNH6s2syTZyjn0579U+FK+iWMq93JZ+BSR26mprWcah0H8wKwDN3
qoixjmSe8XK3rcgwjPcngPw34AUR/+2mDGMr0scuvlFunV8c5i9N4dypUJ84CZIN
u68LXSRM6ebqk/gLk1w5xpGHGU6HIe95HdYKgEHYWPbUkOBUjXldsqq++bw0tCCy
LSXIAYCadNUtLDeSGf+kNzMxyxkZF65Yiuh1WPIIYCDbKb2WviLeA0MEIRg+5kCz
o4XUUPwO/O4bXpmXR0lw1U7S6Xr9Wuc1Y6s5GCZ+ITRY9irLrsvhKCs0c4+Kh460
CVkRPRNwc+awQIb12xguZjGqeuV86qsMiTOfWGC8CFAgRJQ+09ffJPBFYDE87Gmk
goFbyC8dXWfgXKv08mwhcTT6Zi0M4lSYGPwcsJUj9P/EZBNNvwU42E4uGQfAyswR
i7kied3bQKpJ8wu8NaHysIEgAY5AQZA5FhWqkXdqlYOWb3kXxtA7b7bUW0JKZGiV
DUIsyDmDUCSWCNf2yfj9yVWHY8RUUTdx4K8Sp5wn9fiiQFLx7k68T0D/55coEAux
T5rKpHhsJqUeUDFjXh6ikcf8RsHkGWFP488pGgL/Ww2ESTaoRhK/7l7oZ7CCRsSG
Cy0IM5bLwadMQEGinBvr/g+7VZFZKDGdAzLKpioy4ZJCZE2wzvsF/dm/FC7mTf5r
3h6X/eNHs4EnrqMZg7JFymPDydVfGYwEraCdKXQV6WyH6UJRmHY1n763oTgrduom
6yMAYQRpWTsLNtKkeQzozCo9jw/XU3Q6Fxp2Nk93NbQmdiNO1URWeNt4O7B6jrhT
zaGp7/rs0EiI66OFBF5A8NLSniFfcMZPvTtS34RKDu4feh1hb/DgrNQZ3pXdca7C
JYeD1FDWN/WVYTHCOVfoSZciXnqkR1J04ooqtabIe56IlKHgdzJo1n7s62PcDxli
KnRhrUm+51szZHiXe9f6QvQgsPsb1FpJ8bcroCVykuDiHUe6EaEbB4R/O3gBsd2j
NxfKe5FqXVG6JBXyhViKFQxvJlLssNEfW0yB9ytX6JwZwRl3LG37bpM70OqNNVEM
FhqXMMHLrJkbH4LqPUKI/wFh3q0qBMvJWKiNLWZ+N3brrxL6QkdPvv57QQhDYdof
V+a7Hifoo84+aUtStBXkhFmeKTQcYH2ViC4HqmLiL7fMfRMyxIFSHGMSu0uY/g82
bPb89L+ZxmI4N2vqUDbW5n/MxSn+gPo678ay6ZI9/rZliOYANkR5fpU8C2JPFYIn
/9Z+UwOqvyQFT3vxV2axHt6FKlW++fwTdNNF3MnfoZiQHq/8d2tzWvp4WGVg0k5C
ubufFpb/GlKBMrXeQRfq94V3ipl3eUkez88+u0saoJMhtq2+Xe1M2v+ab9GjiHj0
qr3XyJtLcmVEn82bSxF17oJSM3PuoLxh/4wl7PBygpYciRbNaT+mhw5iSEQi5srC
Tp9VLmYPLmgXlkooq1DJAe+Wj5MuHj/mh7lFjIMouy5rTCtLIQnLp1+wUxM3o8EJ
/yuh7riovgsR/DClueEte1kj/ytNOqAYedMXZL9wRJr1IoImVSEh/PHO3uNK6b9D
/Gopfe+J019e9bAXivnIeoFmYSIhQa5oogYIexuKt47LjJdMSg6k93ZlrH4hqRfy
qceNmHnmMA2H83cQYSCX9r74WVbuGGajQbHhhr+F3ONZrhE3e+YoI6Pl+tF6xzEp
eI1Sh6Arsp4rq2ZV6vJQir5txQGHf28tV/JoTnybUzVTAN2LnfBfObYFi564SunU
1yOHL1xLsgwh+ySfKyiSaYc6ngQyBUGftikzN6HCYj162tVPyTxdt5XPzy1Ul1/o
jmL4y2KXjBtbEpSMQKMmxJVv4ELuX3OMU8NPuEkbNfSIqOFNbZKs23rU5lvbFY6a
k8Eh5DwyfCwTjUQ8g4Jj1Kx86ErIEcC0IRnCgyenwGRf8Dvv1S/JVsmNfEYrYEQO
p6zIra4jTX1GoVapD/uC4eREY7Op9/qaEbq/teRaLnvmqyoeQq7g182VSxkC09H+
9Bm+xWMGbaNIYTfk5Bn6cpjv3V06UZOqf3m3E1jHVcO4yofeUhTYLXfaz+0s4IA2
JYgcP+OtUnIhdHJ16VXDYEc3PebfK/DC18z83mByJGE86jQatt6kibpUY6P3UALC
C2dCh+0gVq5TWThTW5rk5hcYUZAWQ8MuSJK0KLrDGPbArvMywaG8XyxYJVxYi/37
a7f7PQ+vUzebDk76zVs2fCwbFmjaTP4My7phsaA2GjbkLeYK0Y8HjDTbzSe+XMDP
7lKd1gGDvxn5VAa/bU35/yaWYMTI4jxJ0IqWn+5qaXRQg25SdfHiQ8H2gKQUtbTi
1MShuM8wwTqkuZZLldV7lyVqDFXxJTQDhdznED3/yglp6ZTOnfWAekuW9xQCGhR2
PaqCHJXs5SNBLIQeU/H47AAviEx/Qezo7kuo3L0f61wpu7fTqUGQ13fpxNB/8tKW
/QGB+8b03n0CGkDS/QJycWcxNMX1XDZxlEO43pbeizTy+x5gH2v27YtCqnsQ+B18
HXCYVovh+wYARJsKct4RIQvIU6iRe4whzUYwrC5Ji1hRjOy4QH0o5806qK7TE8pa
P6jBhaboo4X/3Igfu24ewCTfqZtlaIjocR90T/jT+fEA02cqH27Jz83TnCEF23+K
kBdpF1eZBHI5AEnaJ6ILkYNt1ooXvr1svz2rN3Pi5iU5yAojCyjSCPnWWpd4Wgva
JymhsAxAjMrmiq1t+pRTY7MVGPtkpI6EWnAnrPOSphlRXnyqMBmVLUYrfTYjcKyY
1VaIMmUlECIBfcy6NtMaMu4x6TTi19/Vke4cAU1VN++giZqaJfnsra+i840Kk9Mq
s0VPyygs7RQ2GOU7VFaOaNHeoo/AJtdSjXNRdTQrOt7U7Z1CkXRnEr7Z2lyAm7t6
lhKyGX6cfTSOnFS4FFh8ad58WaZ/mjZYOm5Cve58H3WaPVuSxnJSvza6+8wv7iHv
YGNfV24yVrMdRxPGl3Cj+xHUw3nWWQKjG/wUOzNPwWN3kFZLvjujF8JJP7yMRCJP
tHCKB6iJceZmeglfdjYUhDL3XZ0xTD37xM8zu8KRVzkulKAkmpD2ReGcrLPKngG8
phZgYSURch9WKp6Zl/ZUq89JsehrGM8QAl5uWtQqQApz+tlVBXz+3voJxIUkqIoL
U1TE4a9p/dr8dEXYfVKuxv7vj5vemXWcYzKbbttQvAiJMDnjsJLdnzKz+C17weNU
+SwxbEwgSN5SXQUhVHfCWmTrsTPZjRaMQEiBHQofUTNMMzpXHQI+4xfFxR+MgIwY
npc6SIN1pyLuxFWbNbNpGtQt5Xdaci+hoLaexEHqHadF9/9ieDKMd1KDD5EDPlkP
pCBFQdE+4PFGmPbcODSFnZydCrjw7GqgwTSvcHLz6HuRXkdA8mj6OLAzbaP4I0M3
wC/+N6+qE24iZvzmxnraWSzaIV7jMLu+3TQYhe8HOxw319XdcQ3ES5UqdLUvhsSw
HyA8Mll7hj9ts/S9wRXxIRLj/JB26HijEcxV9f1KJAlLzKg+PNQDSeZd8Z3UAgdL
EqI9Y9yLY/mA9awxsGl92/IZm4JqUhRI8f3a3mdOJtvSsXbyUGR8Z2iH8s2wrG3y
LVeHLKFQUvi6fZjzUoMtiw5q2TPPbof99gsqo6e3+ALHDeSXciC0nbF/8ET1GjK8
d08qd320J0lyGthWGbCI1tQiUv65iVRpYTYVgu7R1eBKefiRVsp5jA3YFr27WpAi
5zuxphYZCQzjmy+rWAV9ZIi/dhiZm5bvWvSyv+vP1daQKQpQxpZUSbriwRz8K7Bf
fkU6d4HPVbrvujX69iPbIvdChCrYSr+VFRUboxgXSRHJblGvT9hWbk5Qeia+w/lH
3l68RLHmPtU+sO1f2HOTDM4mrW2Mk+XAXPZ/AaqDaoG6jI+0Vd6Q8BF1JuhNOhqA
6ngW19NwaXpmk5Y+vqEGAWa99s0cgPgSYdGlyvP9M46GDi/4vsn4YtLrNtMPQEuM
B/NY9NcZkJuZnJFG0Jg09LM6ZctVx/+DnTxkzJHsomQw9vYQT/p4rRIogN56xMYq
3lZR00hYq3JqKctrcf2M8oZEN5eixZg+Hk6gLNoUdKTWge/LxJR11nkIF+Tj1Cdf
wEkmffVe4cWK2ZVMANPpnq7Wz3CxbQivk57U7ttIUnlkNe/lwslVH6MiyAz2MV6T
KwmwYNT0A0U1t2Bo3aq5IQqdKutVGqCabP8kDdHLem+ZAuAfkDa5sbooIhj+c5o7
rWHp+EHG1feYPWmII1WNOCeoXe1BL7SIUOvNrKsXC3nnlFHAgsJlMYpVJSW2BhnW
5e39hTz/NAciU+bppE00tD+wtZDY9ONJAXNVejKY3CKON+S7ClhnIbRntAuLISfJ
GVoOf68TjlzBmf5apnW/G72lLB53YH6LUN6iceRl0xJZTutinNp0RayqnIpPdGGE
3inZt98M9t+RsDt3JLUn7+D/S3/KvSlnz8aoV8hxtaXZ8hwQZz5fDToZn1JHmYfm
eeS5grSRGe0wVgmr6PH8tdXhNwK+axGJfRB7AI/P6eX9VHkBfIlPZEfiGtD2IavN
SC4xv4jur/Y7mz2vfXAVhYtlatBOPSoH2s+pbs4b0Rscjlh1KaZERuu5Fz2AL99Z
Le+TRXJHTDkStads2hU7BFbMQyKjYOxnW3AeOjtt9m1DfUfUh/lMDlH+Uw8ZkW8S
oEmUE+HN/I3ecrFAWX5gwQuhADaprT/hZmTu0a248TzrE8Pq6o+QrwEU84i4g+/u
uyOXBfnlRL2KFs2xrEa34CzABvHiSF67aT0UDFJl8mcidxedF1AFszTwHKLKD8or
pdP6K32xfbVjKJUzxK9bR7QGX6zF8iVVmXYuQ4+6ERTTaFkDvy5g3SZX//vKCxQo
JU4RKCyZnf/ccnt9/ntVeq5RiiZ4HPPrNk97peD17OikpY2t1kjoTJHS0LC6AZg1
7R4ehVaix+MYlkXxQbg572etbE6QvVm5RJgkRgvZsPaN/4E52FuOHtjnuKnbYVUT
VZ3IqLsDpMkmMkRH7mb5leoymMgCc6sJXx7fAIpNbDW4QjBG4UtPxDwsbo+l2JOF
VDUYyw5gLP8AO9qbt3p9A9RjAaZeDzPLvPdHU9eaEMSvRM9Zko8ZJJI+vpA0MNW2
oXsdwBWQUuAjcoW/25mgnGWYGNiciFHLGDpZ3YhAVUHaNniG+WjSxQY65Om/sY7V
rA2vXuf3pmB04VGpq5YW7VVKFppbOrdotDTKYortLfnmzcNAJhrIGk0GsTkN9+Bl
CAnO7wGEHUR/HbL4znaDuDbDe1ijdq9OW9HuDTCCVnGiY6ETT2yQDsUe7qSOFVl6
ciqTPC+J4wUa54VEB01poNKphyFAaj+iBSSp5/8F8B8RfP0uJn7qGumUjJqmEsG3
hTCSINcyivk/OzgUzqiyPmX2LW9bLYW4wKHzTpso2Y8+xCmt39Sf2SHSdHgA9vXd
0X2CgcBQC/3os3k+utTJkKseAqtzLgXKhLSfGw13E2Spi4rqDPFEQlPzmiCaB7Y2
JfXjIM/ltpgfd/X8fG9Nz7+HQZHhKXFBFn+Etg/BzQQ0XvQeRem0fyYSQVozvwDE
8T8MKs2XI/UCpX0Zt54pCC7oo/aZ/OL/bJit+pMElgh2EnMFOPDyC064ca8+Rd05
bM88vT2hzzv1m+Ja2DRtQmCobP4Y53058GlpWFXQBT2OHI08TsU1CvmVfv7iAdK5
somQA+scPlwV/NUbF80fv1Ov+ctgu5cNUW1j9EDMA2tRgGWtUMs/817PgWIavTyV
wRNL4QOxTQg06It/7rtv9ItHNwT3j4tsl1eskcRaOl64YhLawlBr+MKFoWvbUA/l
/SlcGwkrJNo61Em2FxAUdxco+Qrude+OMEYALWC2w1432h+ns4QuxVhHhXZ0lBxX
pHIYHSIwYnS0fCWCl+CxaI2nHQw7ALNP5x2UlkXqjswP1MsPWF0yD8dH0DPd21DN
IJDyl/LwAsImzPzu3r8Fv0dF0ogsXlAWsSwhZAVwsm03s2PjydwFkglBzXcZIPaM
eVtdSJAorC8KCP2wmL2j+RDG3QfWmwScQHH1aEBmzoOnFS4xq2G+5JsQARwyI6U+
ICvs7DkU9MR0BsA4ocHhR2lgukB4l85ywJkQ7l0BLmCoCwuZd83gS/EWy0KRX0Zh
N+zST9e0g0n8Gnr+zwUGJSyGEMaawsuRnoNmY6KbHsH6g5kbi41yfL0U8HLUqgmG
4JSwYbq76HxolGDLZsBDRaOZbgDKRfHNiukbiBSbarFQH6Z5IxcPoyaqPfpYNRxt
5uRJtduvz8CW1G+evTIRdWNbpSpRYXnRh5swqShGwZQ9iPC0LdGkhWt+843qImer
OMitIRcgNAmEjKdr+0GkKZfqXH1CWWyWmKvN8e05cxFeGMFRVV/FZiftoVv9KSvo
NmUqBSKqOXaXARKRryIO69P3ZrsXu1u3vjJkj/c8dLGNvpTuspOrzLvA0+5vSRES
svIu0ap4vXwPnxM0fsSKBZba/vFQrJdarzJa640yTapB/rHh9zv/ZgHi3ZAYPTlF
wXs4qej9/OKoPTLnMDnbambyJcKwTvt9JFVb8yn7j7yMt6oxlLLRaC7HzYxXGR0V
YC83CkXRqKf9fBP9St8cQ4SEugwyBaXUVieOW0Lzi3AUSF0J7j3gK626qAexBpir
/Ct5N4N54w7/rcE0eTFhjPYkGGTzS9797wLvzpPSbi4VznVgx+QxMJ/PCBe1rUS0
/lguOJ9na/TnjdP+GclFu/BwFIShf1+un0Bil72Q22xh9jhVw307Me3FYml/0i4O
EqJzf2GUpfWJ8jyE28WWyijCNaWzKDV8ebNl6eQP0oPdjoM0tAKceYdhn9Ox1VFz
f+blLuBV+c+dK00dj1x0k0O6i7UQn+ebKLR91WgqDTQq9725akRym5oGRSxI+MS8
nklBzdufJIg1tEwzYol3TYzQKN+HSsYirFQ5laf2EpLSvK738vqRkP9ar0/R2zEK
TR7R0ecIKnqMOElofqooWdhSsCURhQj/vxK4geXqmthPN5ThuzRkFLJ8+LL+9PTB
bL7e1qYVk8n9FRL5Uv/T6bEbJWK8jsp1OGi7GJaA1D9jOUc7LEhTNIzYQAmlpWQu
zpBQ7tjy3Gp1i5rUCOxy1qKyut3etItU/YdRnn08xChRNTi44YxI2lnqA7s+rSON
8RB5BOQ3WrEdBzW6u3ucZDgeIGb3/KF+yBkaWWVdg/4PIkKCOarfxLHipN+/DGqw
D+6vqOG1JiTud76Pm5mdqGirLmefEuZSdLayMV0ySnuy9tbMoe8ATdGheHHkgqsM
sREcpTyM7AvFg3bh/I2x3S7sqso8YN72oWp6LdrdQxTwsJ0Bj5ztIT0fWmSGLLG6
yOnqFgttogiR8XK3ESy8B0+w6LGo96I/bWqPZSHYSFxIyK8PlIJ0LxCaX6VcfhY7
E/Vlv2pLUamllRNM3pNW+RMP6WJ5yZDryHG7ib0YzLy4mczA+f3ahMHpHeoDIo+a
OcIjbu9ymPfccCfSMDO49Vre29Co2ALS9PjbQ1N9wrv7G1nOseRjE4utlzO9jNQA
QBiz/WMaueN27f5IkO0cM8Wkp2AN5iOllyeHNC47Vkszo351USRCAOlW86Rogx6l
WyuXMhHcQncc7qDBjjR9p3jGRin+jgGbJrHcUtzzAEJk+z0WsQ90ipyM+2IYAp0o
sZTcQSRvPSa85DecR4Z8mLuUv9b5kMlE20hHFUKlDEQJ1ckVs2QgLyErRahXWyTo
qINMASO+GhMUFxsq3o607b5nx5JzBqFVoAL9GRicqMOsA+0hq2ik40UsGgrt2N2R
qsjuCY95ZonajtHeGEdTcV+oiubs0ByVK6uYtWOjvf+ackbk5Ph5mpmrDw4usn4U
baSxZHZzzAyZlSC7NN67kBphP7wfE6zo7LvgRRvXj5AcpvQ7Sx2Q4I86G1Z12UyY
d4/QlFrIRlEOIBP6enMAAXQN1p+jlNFVI8CCmGK+nXFcjSE6A5FT/mR6vT6woDap
ksZS0zPpYDPsRAzan5gXtkp3E03x8hLkZu8+NfY9DiOZP8ar7nSmJlUp7PFACYtJ
gUni4ZtvS2D/YxC2qY0siiQh2Kh/D6+mzQcYrw+/bY08jyPRMikZ8sgLJ9jrfcHD
bKVPDnaclMM/cW63LWKYc2UyLjpS9GpnSmKCEagm6zYnMUtQOYhNJh+QKoPQbE+p
5JroQlb/x+fgp8CmYFuGlCpiYr2jmxI3ejvZnMNqyY3dExaPlSdnRzerkxL1NuWu
KEX8AmkLvRQFddKS1qpG5JuAVYgqN5njVBys2b/8QGSErKqdC4DTQ0auWkNF5Rje
zMpOwupXuZY8VawFQtnNY+bNvjINGT+Kpe7ExtieMH7RPd2tmLxL9lCLMOq2WQta
HhZOfWcItg41OOFID8/TKPgxlK/CQnolm1TgfrraPCADFrpdf800WxhchYhxoH2+
S2D6Z0FKtveM6VaGpeLBxUCF4p80gWbVrAu/NRduqW3AqTStlNQxTX7IuHGfCefD
DzVpXImg/UQ1ZQbWpMWk2xYxtP7ldgIcX7SFi/UWJCJunrJnAkqMoY5yphLH9IFd
3xwtIoQE0X9AYTkO8kdWL+ctI6u8rQ8xMZKU+aJZ7U2f9EUqFqtWL1lJS3kC50JR
iJoJPdLFQnCl9jIxmS3PvQq36q0BxkO7obA89GSHEqTUaKJxdTmlPLoAdbLVA+94
FmHHleEcWRNIMKiWyzB6XyTAmdEAvOo0cvuBlprDt8MvG9DaNY8VCrhanrLPWQ+0
/As0NPVUWoRpxQubFOIHl26ucKa6RJ1ySScdCdFiKNxPpv3o6mg6zEW+hTNaipRX
K/jH265pIZy7w+ARQGtejiUixH7468QOyb5RDEZ7hQV751EDk8U6n5pBTz+azYpW
xVdOfuSLOoXKROxj31xyVv97ymIXyVTf/Esux3J52OgO7+tWX8hDGgjxmeWzt3ni
4snkiTY9nlbQNs0XBy0jNhuBWp5aQFPQkrw6eZqNHQHFD8ct44jHwFtpBcX9fodM
+RmwHUiV7N89yXStubniPmGHXxsAwZCiiVlarCQP/9+9eSeCZdCZ/vo1/J3m0qya
h1ImUUgnFf7PhO/DlLB9zkb8IneS79zKVHzU8TkgqKGz0toWyBro7K4oF+CIqfYl
2ITrI63e/QogTkF/598PYHWIgnXG80xkGs8UnZ97zUJ9Vz5JA5sHOA3tLO8b5GO9
NveJ7+vUko0VbBH4eRvOSJyTn6H+fuOmm/FjUveM4FbFLJD9f/NgS3DrXMS2E30a
80xLnneycmPDs6pV6m3wYcrbKUpcpCo+3Pv4VfNIYviECEoXmttzPl7uhgEW7BXc
OC9en++Na9Qz3121B+uKtyh9VeaoIhMs/FsuDa0bgWgAna9HgJ+LStlk5VJcfkZe
xoLkDERwu9Kkt/W1yptkZ2eovbshvr1D0vCE8Dr5Mm9mNRdGWv+sHXnJnMG8qKBY
9D9klNQtBce5JpKiDTImQLZCcPClHlcZYmQgTHZwyESpkUsvDVtjuHcBcYN+yAWj
KZTuV6465frh0bmKSd9l9FZOJbBtPzso4ebeIooXBAAMHiqJUNG8a4v5f8vFtnsX
2tj3J6I8+BwZZXPG1Bv6cyucY2/cRR8SLp7IEpH2o/lQQwR5jze2S9MjPBvL7UXV
akY7JXFyFHhnpZ6PsgGxTA9WTsEHcv0HB8wBAC8EerG5u1EsXehGhDjmFvZ9p8XY
i7OdGZUcc3ylbv0EQ1btyBsWZkFBwVlokY7wI6xV5HxLmCKqAvy3H6Eqcq6fJB43
+lW8ZzPzsZalzv8R1zznNJJjtGVAJROe6XY60yENC61dFHfKhBF3agO5/6eK3LgK
+SkTs4yq8aqcMIbblV7GDs92Qu5gDa/dZJaQF4j6MmRW0x3wcnREpwrxNOwaX0Q/
+1qy1jfdm75Dzub6/Z7F4ZtBrWFlcDQBAATT3DGboe3aMgQ2Ium/rrasT3MMFd93
tTizBlEj60FqkGcJS2Z9uh2CUkcSQeU5nofn+33ReTYBQzWdnzFCp+lIR4OSvN6o
cboznafSbVkngMhBUb3YcoamQ8RLzKB6Pz39afnhZyzyBEnmwfVrsaz4KI/C3YrN
irBTp85TFMW/FKr/5y7969vWZNmhuBvzAU4nCWhNTM3RydFlCKxpCxcBCB4djEYa
SY37QAvblv9HBuM1zc5IjI9td9diBxRCZRmWLAV9T5hZXXZawAoTS8nEMFGDc0AM
/jgweXOX1NpXfFSeyxjBtcASvj0EvbfX84cPJtdfWRs6gtlY8aEdGsab/jFTW9Ba
DfMLP3bmjpYb+26SXweiC14ERvHScbJDtHjZO9xFWOWAOIZwiAYMeObRM5P94EUZ
/6VDQaHJmwpNcrO3G7LkTaOL5DYIUNldqL0zFfIPiJQldtpwiN3sD7hsH/FMD73q
EmOzKqU9omqFCwVzkjfKOn+b86FPgb88ySF3hRMsCheikaQSIEOSjOKI0vMI2+OI
RYt+XikPp5pw/1Q41c6MHe58bL5eod0g6kHwpGounJO+xG148upEwkPHBAIgahgz
uZBkIchPX0YxjpI3bTlQI0nSzMuIuFyImQDijhiDQJOKYZtsGdvUuOrJJbg98OJN
Hbc3VHqxYgomMPbJ9kSPJJAcQycUlasKgBxpmDRjffAHybq/oqSFyHDwoUvFYjVS
h/sZGPgOdbc4Clr9EJcsSUnjNMGKZx3Qb1thQK7UOzgJvpLmjUIXprQqPRtrqq0F
Rt/wOzKV6KIOSi5GNdgEbd68/ja4ZLueGWqdQJFMA9HOtBsHC5ijUvHRAnd5sqMt
TV3ga4fTSm/LhzGnDD2AC4A5w9lpVTLe42xt1CT+JUlH1ly0/rW5sLBgsjFSE949
bFUe1uQPOCXiY7XAaEe/YKCBZrMaUO+FiAhsfjGemRjAL1XhEie4iEeewJPJJE1E
qiErfuenVnqOFkD4PkBgTczsHoMbyK5svm8E+nLn32z1ecPUonqr1HKP3v8dWLcb
W2IP0umVDQamKBv7957BQX7NGcehloSI0VDyv86ctbOaFLJe46i2qHdlamt2MHTV
MG+RcdZcCEqSGuOfU3Ckb+unCXG+vEb3s5U7LOwypfZmAQl8zX6gSmk7fGJnz9RI
9o15OIPpKrMXp5YT6v8jf377MIPBRpo11+antLgfVxkjWbgSbBEJca9bIh63x9/J
LwhbiVgm2slg5M0/KpqZaPik3mZxUU/W07E7YCw7Jn75xPjdmUMZmctrxm5O22La
LoTZJlnhnbA729isr5xyJg7Iv2qNoE4O9E87r5Dgom72FdWjAAwZwMRXMGdG3g3V
azijovwkP4wabW9oL1PYmblFraYrV+6jSysqicZMy7TPF/DvkU7+fEXlHY+BksTK
dLfzBDr2SoPXjHOjknB+Lw2opIdzz5sSDhq8VJdBUr9FRs/SblHqD6BZzVgRvLXG
L96fNgvq7IJ2xzKJ67B8JFq42/LKH9sEjsqwlgzGHWfIh2Fx+on6FKoidnXGdctg
uKgRA1UePC157V09f0/twkaL9U8ZlJ72Vt2Z6N6JyYgcLm+ijAiQnA66PCFdu0Jf
HL+fDrvlK4T16eQeoyatz7nUi8IZi1RpHpzZCuS6/obRElxPTg+sfYWb513ffNEp
ny7sKEo0VHZ1RI6GIZr8w9LBMl3Ve5p9btRcc4HF6b3QH934lpdirWJTocOU6kjm
fdu8miDLlwE0yG6vrCBMTv85la7C6V6TnrsBktK2VlUIlaBne9RDgqLp8tzGvAaY
7x4N5N5lmHQft3sylGHe5sOsY5xCzRKZLO8YjzUOpVcHqmkRkm5xCwvxMfcH0rfM
WkS8itgum/G1uuBblnnA4PnQDS+am2yDp1wv2btV/wRbVsq0S/og+pVNEQxXe24S
d23V5ch1a7Dhgisq9jhk/9iWMVcaSD4KHdj30tcHpV79zgcSSl9nk7LH/gbm6ZIr
YWmGBT5T4mm1eHhFoCqsV/VHKJRmT0/sP8Yi/IQJurgmEOifHA43dQ/U2h9HXyn0
HkW4yCw3qajmGp1FTQAP09TZONpPoVTtA/3MU71YTO60jCaxgGEax27FLMDR5RPX
Tb8EzRK8pYzRojYfXoI6QbFCh1Zqoa7nK5uIFuQpYi7UobnS6C1ivAImi78vAW+z
f2pWSHguUaXEa9mAnOaVE77JPkRUsavonvQ36bJwJNu3F9sd3eFNyMwCQsFaIqnH
FraHFU96AsOQu9AsVZT/4+z2JezMpZ7EsDXmoQZ95schb3TaDYuslIq2Jqit4zsH
nM6tfZm6qykQqf4lK3dTJoZA1mujuuC651LHZLlmE2suc8p1c2kqaUZFbYxYuhhz
6W+aI4AA3sMf6IkdYVfzkvhSH8M8qQIDDJ7mMXjxBfjhWNMMXINBkUA/NfTcKWVj
cNe3bUG0z1hmkcMmiqFQQMRLS+JlV/F6bFM9nDIIw8QqTZmTEzL4d9jaUPo72n7x
B6n62sPjITwQRU/Sd68+KEriLWXUEpCBFroz4GdA2jTddR1j2BG1PuhwhwJOTZKi
e5AUSI8mxXdFxLDhmPXCmgJ3yv3M/GUeeoKq92rsgy8kp5/E54M+kjeFlfBPC/qc
HixXwmp0ImfhYYRJWRz4aNUSw9tW9C/qLu6j5kEwmZPj0+6sRwBGcuAnc2MQ3qSu
MIKLwDGo6FMUhMUW556NWJ/5pkd11azL4qPtroGjTOeqm/BIwlkpAtBsHL0khyCm
xy/1Maoe/zBvpMFGQ9WkMqt/+GsR3PgvsAObFlzBB6FjuthZS8d9fID8TKwi5A8K
8b6gIa99Aur8nKqT7OAZNiFfAvZGES8u3nYrfrubhKPbpWIfP64snkZvB0/N+tuF
1aYl5G9jLHRsJqF8H8j8YEWtv8tLTB7los/F4u5ZdG+G+VxL2SiNYkO5MVguXr5b
yVeJi/Ghr0m+24PvPisflauBgFDm+D0AdW7fzW+g+iKxp+szkLnn8QFknc5KFeYo
WvuVQBrOxeeF8f4U71wC7xL5gmeJcFE99hn6Swu7N8l2rvP4ZnPQbfvgxB99tX16
TAGA1cKGFUEGqkOp/QCESRR+pESKBEnjE7CJx9CgbTiAXqu75+8Mteya4kLH+9Uh
d2UodhT06wyIEUynf8C1S5NEFTKmsG1NW3GBB6+eE2yzKQX4/fYzp2DD51nagiVE
FzCLqMS/K6rLUw8fSSNNcAaJIqMhuvxVXBbANQVSvCx1bYO8+TMytePqEPfqjMbQ
irQD7HRglmmydpbh8mAzV9OLN2C7PX0Kt/ZvxGwxiAq0wg520EuZIYT6Hbb01JR1
on3pMLUX1/AJjD+l6rM+cHBaORNfTuNkqU52jXB77IargllcxlPyZlK1wq0wQrBK
k8HcBOaEby9Rrz+xIU085As/dUE4o67NpHpxr/VGHIB9XBNM5G3wzKp8FFUpUG5o
gJoPENi+Wjeu4x8HgDQeejHBEHvlIxn+H2T4uzcp13cq+OIxK91HoDy6/q+hXoYz
i3EqpRIWL++eoXIFSB+Y09SD52bHelf1crAn2HlrcEQkFy/08rhMMlxwVKm8Jpxi
Uo+vNtURR2Hg+wvFa63XYWjSjHIcYSNAPj8zmzk/IfCyAs5qg+0ZR/mygWvJ2ymS
j6XaGtwlRuzZ5TNC84LCypsnhurWXCe9BYaFY+B92MCI1yEghdVVjn5LnGj1yPBk
EsDyWkBNDqbUZZgjqYQB4G8wnTC4WY/j3TMiPgQEmlwx3wTP8deeVac+8SsmaFXe
73zolgkT3OM4YqCkq7AM0i7vsGQl6wLw8ncTOBquYssE7bN2ZtOSow4KmsV5FPBb
phFnA6HyLlATUcPQbLRMuieLmWg9MfUu3uG07sc9bS5YjhhiypTAhMlVk3elt+MC
T+uQSKFtjOEQc+PkJdmV/OZcw2vvocGdCXDIkLc5buQvZVq3nZz4GugiUbnAmLU5
cFyuNwobu5KN7z7HtBspygh+/TwW9gRgdry0VjJ1Dt4aVWrieKLOTNmLvEri01bs
UrQYB9XcQbyYdJTFmMBEEg5iOSWOPa3NIKNqFbCZVTNc9oO2Lu7/N+E3xmhoEP6N
7mpc/HdYEK5eafmRshuy+K72Qs5FE8i1ty4j14O6Vhjz6PBo5d5DbOQSjWOrtTpX
rwSapxNzdKfnioGdOn2lI8JnllV5JW3PIPsvQUCgpsCriQa1+oidIFc5jME4+/TX
CTuHyczgFtJoeCIKg6TQsdohbpNA6/qFIyFCED06utKVxUG7b+8pe07X0KcIcDj2
m9VFHe2Z0OxOG67ygckW8rwVJ2hhmUWTVCYyEIm3PAixpo2tfhfYy8JEh+YCGRVr
1RHbp5zGuWQ1SvamyPAqUvF88t/uyQW0DHXNLES6EKIJNVCElZwldb/a4YAwp+XM
TEVHCdMcDFsLw/q14khJQAVNNvu8mDutwcNQCFIOQKIZYKLCpg1z6pr7o5RqpLt1
XtGmgxhEK41MKEZwqoWyE/gCWxGCB9uBxx1l2er9qhABrNXEi4HPz3pUs+unCf8k
Zs/HVxOZXP7vQkAakDx8qoyV95a8ql2AsGgev8Wdb/w/Asuf+8T3Ix9SHPjQ0kIw
tzPF4+tZBptl4PCxSPQQ1rEI5sSW0+vk+8ohcngGEUpT0xrTm1ULJecCHFOaD7mj
GTlLkqocETAKDTLGt6PUknkNb9D1+AbV6iSsYIj9IPwY5tQgz7nG3Tq/oj9d95Iy
DuzBRoZ7lTRZVxu2qwCajKzQRlv/hftuSwWS/hkfhF05JjPnUA1S6qVfflyfmcp8
Zuu++eGnsJlmfy3lk1MebpHXTkWpF/nOVc3mx9Jq0VlrEgf6x47R9yjOqS2gFzKc
IoOcdu0gH7yv8OBjvF0jH5WTIQaTRecZvredDaM2PX/lXYMthfJNt8e7Y1Jmm/A5
HGKv8H5n0Wdr4VcgT/hQ2iSSwQEZNIStSOsa+bh88Z3H+PLlGMaG1PHyupLRUUBd
NF5qHfAiC30pemSudOpocTZpEmlsrk+FspYdeDno+yeo2mvqNWBdvoWXEmAMHJxV
rCuTHLR3LoEtPdGGywQaRbPmz+7moUxfOk4Uq4+aeMv2REe+2g0fPTDRJgzj9fnv
2qPMCE/F6nhmOD6nfrHx0eHC3eRPZYbH11GU7nXCkNSgd5BOhtU+CQHW0b0hr0lz
LFaW6Fn55fl7GDEkhjRY8y+eP1rKPvHAHKvDabx17IgEyJ45V/aQXOHnbMitMr1g
88oiDxW/TYSHrWb7HI9JNMn8/V88LRN1L6YanAvLXH4OZVO6tU8SsY+RW4O9s2ts
fW38ZVls6HQr5cAX22FK9u68KFNFsgc5KK6INJLFYVzWWws0UX2gf6qkuVTCdm2h
soglDAsjIC6yWh3IiDuIzIpwYKHIitKui3kqROV2UwOmCDf9Mtpq7zzMPOFji5+Z
jrOSPd4gYL1NbZp04bfgSBDI4U6jWfXN78BS9WLvtUJnPf1MRzk1B3thDn8eX0Er
xXq36i0HTneoppS+EgD+cw4ChKNP5SEtm4G5frMQHv3Fec40SnAcOEQBIj2Ve1G3
V7rFsAcG6YBcuOnAPeXkmGanq8leo1dYCnXO9sKoaYXhoMqi+Fw5O9s2lkFgl95s
36w6ao9sHJzLoFFbT4MgaDQJDcF6Q7wYEoD+H2Eaa3TLxUlY6XK2a1XINZ+ANBzq
+QG9RGH+6D8UdVIQ1KTOok5VuLgwKnFuWsD9ZCsJztAJljsEz1XGqAtMwwm6Hcnx
CjStRMTG2Kt1hW6Srqqq7zLHYYc3AvuFX4+VfGzcRms9cmAVaF1tSs+zDPD4/iFQ
Ts/yQ+TiIOgrF8SAiRsNBh6mtSK2nOldk98kDuvOH0FhDmIskpEgT32EveI7rokU
glqFhARdsxddR7kioioMws5cbV13NwZY3KgiUJKZv9ccLWK+Hwo3x3OW1+5BH9ly
7WjK6+TneNaVptfNtEx9aafi9UYclwKrb2NQdKbp/OPg0XzGCUkU5G/4i9MLZCZP
vdAHKnXQBXP1nh1sfsIqbX9LGZyPrnmmYIYZm1XHhAmiyGIR0L2k+rZKNEfcDsb1
VLm8+ICmnAl/HzgsPqSMqfJmGo8Uh1W7ZuZ8kCfyM3oJfUXi+0oL4vXHRSQwtCVn
17WyVynjNyLMPqQg6H3HfVKGqC4eqCVw4x+PiP4prJdi5iWdxBwN5CPL8aDDA9JG
/OiZzg24es4bsIeQQCfeoV3e2XL24m3ikMVXs/EWzvPAjJ7xjBWyGgUnx/jjgWiM
Xs6poyk+E/asoCHgQnLWVKl+TzWAdcimXB31CC7hiE7qnUAqp9TnyNGQj4X2s4xA
rNokzk+JLWeX610z894KRpPJU3lfeaqk4wB3jLDrMocupijKhmdAlabdmG0uC3cD
bKtZuwZyROurLE8VABa2pKLMBhuz1z6BLdiXWUAXFG8X/J0QfTjU8FFGFICgUCnc
dC/DBT/lnY+510NL29Razw6TAGVn4BvWwKVncr61DWHHkX7qxJ9vINB6YxC5l8ci
wFiGZLcG0DErQLnZmoFWOsVftdMa+oW3lUsSUl67IDY4g9MU8bcLbb/F5FnfZiDy
vSs+/RnP9nMUZ+YYZ0Mr2+LtLHwU8LzP6m6sQerONtwsOwsKdae6iU2ZlOPPV2aF
Z1NGZXBUtceJ3N9SM4qJheSKGkcPv3xQZAcFv2LWTOn6D/0XHh8I1Ip8RJhHjsPI
aM4epAIbdMXcL0kCacunYqdU51Qul9pID4Bc10JW+uPYWMi7AqtRwdbDkem5pbtd
JPLsPBmU8OVDSrNcLbZ7GbrpAEWOKHIwKQuhzhQrEbYtXimtZlZiU3Xnnmmq6fDw
gc99XVVjiywv9rdO3d9/9S9rVJ+cWvaGBUE8kFDowWtN2PxpEXif4xa/wsGe0UtF
YX3sMVSs5fNdrd6DS20F1GtLfOSNkpnmagE2bYTXM57K5Le5Bwi54FOnDuaPs6WA
Z9ty1y3CWcj5EwYR5Vk8iIWh84iCpoA2H7GDcXoLdcuU531JLQ06ZFbSo4jVImv3
9i6TxxB7GZaa6m9F1XoMST5Qr2BK6NejLmqIIYWAxzj7tDcOCizlVZsRBAgyE28l
ergPMqo0lZwLDMk1boUnw6vcs+vCDYKJhsCiTmJ97fUBMgCMgHW8ekOwn6ihb4il
EQX7lMDqAFMoKc9TV81Ke9nZ+kfypkumSGRHKvKhIcY+smF4w49564PX4NMwu5nd
f7FxG5Qua5BQVGSc+GHoiaahEBKLibr8C11DV7BPkEmwW+H/7Wfy1+yBiMRuk5rx
bo/17JBZEXxH1efr3bbEOsMINWgqTFC5sIoZsd0kdKq5WBKvJ8pQHczrcenrMDyC
yTOnG4fWgEOqqoaiHZjABINv41z3sxB0kLm405MoUEbPDHkjQNoh9/Awttx2/VCk
+VMKsBR8fSHWg98DqX7lYk8XUufRtKyq0FXj0LU+F3wX0O4YLP+jhCzfqmAUUsx+
8+vX8Otat2dZu2jaNGJ3mssVYqIRoSLOvD/aCBPwH0JEyRvY24Ugi2qfllIVLbpv
3HRsNUBpynf7T8LGaK7nQJoKY2VFdDb4dWDhiWL/OFbfopKum/rR8qNTTbBdTt7h
ly65AFEQ36yGPnJbvqn0Ff+oazL+irOIVC5p1uvYi3+ItHUplvASO0mDpHdyTGmF
qHYCWQTPSu4MQG51u+5/6eeUGeZb/10aAnYSfN0zAnyga5ZU9lxmSTx7DH7t3Bs9
Y3aJfC4izbs42S/grNwZgWC0lZ8TOL6/ajCnoT81IwymlJUobn+dQyQbq/eVtyRq
mLpu7Q5lQqw8wdv4vGdOqLmWkTy8pxLHjdcO1HoapM9pX32gzoX3PC4gW39SJ9Qr
V8mR6s4fiQ7mzw2569QGEHODhnF6pZcohXTrxr0kdc7sk8BPOq6VX7rtsMGvyP7T
kFm7sJUh1E1nLqWJS7WjkQqm+gSiCwfsKeFj5gqQ28/0L62SQqLC25r5g+NNMThq
jUF0RfJp2uWSHSoGY3v6lRszsoixn8xbITBr248jPln2Sye34u2qsqA/MlNiRFlt
vrT8x0l+hlN7htX5FsKebfLrBPzv0ZGShBansXYPbrX/FvAtGePvlGv0mdXNUi6p
J3O8zG5czMmAxA8umn9xQBAWz54FqI1YbZIeO5WRk4ehGwRT/nWRL3C3PHHS9Je4
lCsgSN8vebQTfBefBlaTSVhHMVRyfasoPtOv4scxGXZ+Hin5PtmXXpa1LfbVAr4F
SVSIyMQyKp5a3oKwndKDUBWoHcjVh7vtAjOCYQ6OMPStzrES9Emz1YKWGYQn/869
DbuiHP+3GsnGKEvQrLq45RzxStIgrLXOCUDbMwy7u0c0fbp7tWbDpbeE2RmAesCA
euDoqVz210LIaFy9BlYOZn1jnAh9Q6KtkrTZ2gk/ugmzK3oSU9WLsWN3lk4K2VJt
62WLv9SCMNqg8SgzIHbVn+2aomk8pcFKNu750Ma2DnfJ4xTw4TglXG2y5Ihsw4zT
cAh5BQHEccXQPySEyjiMXutPx5WNlwOtqgKDjRQAjPcA98yYBtGUCiDaPtJOdSFD
gi3JY1KledOMGsSy1HCkNSUxzwSGhwepO6wuLpfq31Kw2buqxXQ/+C+ArTbqenvL
wzfR/sQl5K3fqk2+SapZM9tObXKbppn2kh5BM1iU3lIiPP2Iz/CHllYTor0cFc10
BYry3eQniq6TOVkRg+bkWrvaRO+I0TjkpfeqwRrakFU3ogWR80i8CHSgEkjMpaX+
qM/C9teMpYx5/KZEY63o44LXcvRX6Go/5tSj0XugsaOXwfQwXj/3nEyYKNF7fopq
Rmw5h/w1U9n2vTEso055atyPst9P8ADNivQf3oWzqEJYLYWtekJhsEs/3bAyTNgf
jdvMt7XruFrUEsARzvGcNHEiTknMR8+MlfRJu3oSjSk7JFVp2RRHneZc8QTM0gX5
HMsK9ysw6pJbcPQg3oTyvkTAXCZByQNQh1ZQ+ShZTILl27i8M7Yybyt4qkWM032s
kYuJwO56qKmJgzPiGBYMZ5pICE5qnIeAjYH8nwizX5VZo9xhGdgipn2TJ29RJ/4u
ZZ8bGSfYVyztv/O3UWmE7vlWRdh7++RaULTX22GAx5gXPaMANDztiovm1TXhO3s3
wN60UuSnB//5rM7sGXukutLHJs1hb/G2X3U2RS13oNUF3ubtLTfDJXKt7Ft9EbPM
yNAhAm+qq145mdwPTb+9cTCgevT0aUjiK7CC7EnY5cxlP50Jlu63/6pzkpT3gFoC
CXv4Kl9z/gKDRSoQa/s7SA4VSYq42cuM2J2AEDPflLo5LUa/7cfXqDiLjVoH53t9
LN8wN+t3IFQtWdTbas0UWcsLAi5lnH2oXZa9skDaSQnoQxrwvbADgAJcRfgQWPL1
DF3ANo/ww9skH1s9FtDIYBg8NFVTrw+kg2VEIbkyEsdv7N2MyFSf2M4dQDWk6SdI
3J/Ls/aJW5zddf6itPeJEa6rUtu5CWXwYsiEEXVw+5JjpdBignm215uZBlVevAbr
uI3CAHRHwimibeePAsPelGdXvR+7qdwlBlirC7PleX7EtB4bvv8QPQyMcnvQTUIs
VCT9ua5JRX//U0NzZE9vRXVEhUXY64BD0nw1/UKampEoDrXGAdqfOAHoo9aJ7I9A
WH1n6t8P+tzp/CDbs8Pp6fkh/uVqZvyGPeE04vK5Lsy74qhsgW82IWReUcwrm9ZZ
QsJY7C+9QK4pjotFeBz4+1SX47GdK+95qoGRIPYGcMA5A44bRIHl7HcQT1KYwljM
MPAykpcr/wspVBdE24BvWSuG8cAqGNyuKdtpyM0C7adDjGTlyUVGayRPqSW1+XTb
xmB2sVKFGsyjnEl0hVFN2Ds+DG5sLIP4ZMbw4qQ2M1kfMwMi7RyNstc4Q/+D7w6x
9rVAShowXJTRnf908RwJ3u6s+A+9naHLLkNz9SJTjmIZJVt6e4eb33lklvZNUuv3
iU0Hgvj6Q786+HFgkQ7xxpdo5lOGo551/qRO7xxy8sow/TktJHXWRh7YawSh/BRs
K/uJWREwW0rfyMaf+e17FQlYFISylhKK2urqcqFcdeqj//93GaQ5YdT6XaTiRFOD
CHPqNaHeSX/SDtBPHeQftPNwWyd6x99HRCSeNNuBcsUtDQrhsRXxMJLW5LpbEkd+
RdnaCp3CVDxCNu5Z2GNa68RqNmdDFL/EawjfXRQWB8NIZKdbFqeBDhUP6KD3/hO2
xOQgL8Q5+5NBLhFcqXvaHOJnz2I2Tp/qFNTp5dc/+yxman8liqLRcfddp1nVu5Ts
f9b/rTePKIWic3Fbq5N8z4fWxqhbkC46uGnF7u/qwbZGlCmLqV06ud3NWndw2zMi
uMxvVhNA+kzkuUkAIg/3YABWuYTDbW2SsdZ0Kc+bwDD03VeC5KnD5u1mXGsvMxTo
Z1TyYSvXIy+atmsIS2Ai6sF8/TZSTEQaC4BnaYGPzvmeOCkUEpXQaI1GmQwgIA6+
dYfs6DAOo91Y01x32L5aBGAAeJZ0KX+q+DUhQdQ45Mr6iOm1WQEFMhK7NRsuTxc4
NM5DfbS1NKuSYkWCkk4p1f4aWfg0Uuej8oGz/m64Xbi14jt/rLxWx5bGXamKij7L
/+HiRsnlqCPT6IKwhf/21rDj2UraoSpZfvE1qUHgjHwfIjYDSXKcyanU2wap+lgA
ylJCBriXraS4M+IwLejObDqQrYIsHBC64JzCy2rUZcUutPRfjXI3ZfI5bcPPWDoq
j0Y3cUE/kTxDkNv5BYe2MOW15EZrOT/wnLuUTUhVeQe8v5NSEKwUA/z+EKeJLBq4
3VYUWu1mgK2IxP1MB9kA1bmKlZyrClBztwlqhcOcoeDV6SyKJWvvrRzxEenOHKu/
TsTfoEHxKfz5nTHxREtqjZBkkhvzYzPTNGJN772dp8bVs4fcLgtbo5IkDiKAEC7p
I7ZrVmrRArQKgfsu4HZSpPT+C41hQXtgGhyoTpxHZLbpjfgi3+OfdXwDUPQ1JP9j
rcofnclHjx9q2rV1asqw4SYbduhi9JbiHrPsDR3ETY6/Lov04FvsjLRWWwn2B+Lt
zbvrTT1WrCGd/DGRF+9LAo89dmZTherg7xD39WfSYdZsB3eTqNbKR+F6NnHtsOFQ
Tbt3SgdpTYVBrTMd/76+g5jtzc0g6Qp1nLRvCSzWZq0R94Tl57BQa3PAyEaWpU+A
bHrScrb/6Z5nTbSJ7xFOMjeYNHZKYg8xDXb6yjuilWidSTZPEATkaDCymujt650R
3jmxGws0DfQQLAR+nImXFAHEjIeBClWzXomipV0KkMUp6kKqaZRzGk15zv1YQifj
F8vubPQFAwoc17Nk0FqCTgqfWRTvq5/ODC2LqDsKJ8RrNIYRFp0D917HTfOffw6I
9wlQbgi3/qu6AyLiAhPMIDMxzbR+ELdtiSGO6aPSx/UdKZwuF2bZPZ+QP8SrX50u
ZvgIQVdqbZ8QKa3lhFxolMkPYQAgyKHE5bauk0i57/1X05BcpCs53ANeHOqXCwb8
41d85jxk/ofa0pMM9vCFDGL8tzSagf8T4CUJUclCzZ41NIL5vExumot0Plm9+OGP
119SkBy8+cdIqhWKgORHTjis04molDiu2q8JKhm47pnKKWyBzGYqNR7A0vFIbvGL
I9CRB5U5somTgx0z7TDxDbiyx0VMiZnPwUN6DRjCVGMqQ09NKY+U//pYtXeukeBg
TVl9EFOh4f+1N4KTTWrtbiH6HFoCZpqMerGio3v3Fto2FtkAv3bOauzuXRl+Bjpg
3EWQShWS0mssVRZU75KwXAu4p0UNYqqFfQV4BkI6XhOWRM7Ky2z4w/NoI5xUnO7p
h0FzNjsvPrbyyuFFpBTUWT4/vtrt1QvXun9Qm6NnATl6pv185VRw6SC4KsNedlhJ
cmnC1G140iUR6GyEsh/G3pl2NvMUiWErC3rZS5atzyR2ulDLXWhTA0M8OLliucH/
gfBB4o1emCCxr3pE3uWJ0c8IytzhWC0ZDVXqEMBU3NvYeb2bxwzpoHUuPkRuVQcE
0BY1Rgrs9EM7xhEzuNCoF5xVDohuZOjlVJ8/R/tK2ZQbKJgPgf+uWEq5dG99q54c
1sqvW6g0z8Ne3OGZXNoAqnOLCRJ5hZ+JI8TJL3zEr+EtxXNpvOn902wnRBXUvl0A
36IsL8HCK8tiCmOJm71pRJT/CmsiG1x8uhyjIE5m1H+kdq4l0zh65A2syL6H7fN4
Q76EealORwamCvAJXgXp76EX6k7HqHbXz+8b+A8b+MuG3jvNuWXi81tmd9Dik1jh
gbL7AQT/r+xbDXNTDmgls3+w5ZKme/XAQSymKmRLtPOVaKaU6ued/9TGuysu0ciN
8w0IzQX5WaIBYgZyAbzzLHlSnXZd7XVf2nyEvVzrl9QW7+r6U64FHOhbLqwVRkRm
KVKSIcJyiQfxSLaiV8BxdqApbsBkUuU3T+B99GjOfZs0tdDnfdD+28dZD6yZu7e9
Zp6dNwcNBf3NTpjBNfhzRFnmG1XgwP7Y+4UwsQtSWeU8TuMbFUxK3SZLKQ8V+4OX
WCKuViDUMjnJCs7Zqh2bUdKxVQTeldJ8HAe1GbQmNUjA6ouhZSQ+vxXfg3L+ypyW
EHfiavJk9jtyUH+utLQeJT8BAP5uISP2VnXAKyCM9uwB00N62Cf0+9UQgq5/Nqhp
hmC8G1nwp0/lacCP9AqguOrnp286vM3B6NR3Gm9mHoMbaXbqx3sPSgz/smO0B6kb
wtQiDtlhz6tZ9ox2LASsW36UtTTbGKwy34cO1LlBeOR2eg73K6BZDneoZ4TPO8eh
sjVaW4o0qn7ghjM2DWJnDPU+GyToCgZj2gCId9mgLZg0bpurNx86A7Ap1ZWQU7CB
zPpqoLsMhsyrSrwPsg3fPkRRS3YmTWHWOHQgnf4yQ30IzsoO0ZJEPN909e6iSpuT
1Az9xmh9zY/lbKeBqUQNcG1nI+IhYMY757NVpD3uhcvtHQl18+QPx+Zt4QxptAqM
s2yy3m7bdd97Ix81JORLLu8y65LKTQf7kaeWF8+JGEG2gPy+LMDgCsjNw3hOEkAd
O230M3tPCXkBe+ybM6fOg++PpVr7l1cuF4a4Z5Ui/ssVkb9AsaXck9Q5PnO7XmVQ
sVJSDQI2gPyxUaAMgDKjmypEyvcjaNQBNjYOKNKPgKBOv8hiMGSDGVQ28cmDuLXZ
TQP8plGBNzmiprGLx4n385gQqMoauWzSG7B9PABX7JVe/M7RhJfhDKeQVjHUzWan
P1UTJdkGrjZalHVmWe2b7YNF6cJy+Qf9nGMde0mfwYAQk0Pn3pQT7cF9dX23rIkR
vBb+Ezmba42iFBDq/Lia2Jl5pTkX9dFMeyL527T9a5yFzCZ4jNCoTjGPboYt/xj0
ggphEnEr3aOTQpvFxPLgFQpNbSxx5q19/EV61suHVmtjgCGZ2LEvP630JtbfTWfT
yX1o3cyKgxbBs6i2S85sYuY3m0uZUBmmNJ0ymh0E9pfhrXRI9sxSmUY1E98So32G
2jhxCAnRzKVf3jb7GoGLFQUbK8qx5Kb656Evx7tNwAPj9x3nQAzgBzLvpgfW3DfE
RM15yEups0OcJwX7AzooM3C7xMisxxw53n3AlNYZd0r3HPQuUtakv7Y780xkylPY
BbIKshCEorXanbky8x7wnESeboXefZkp9jyrBOxP7OM2wZW3BInqlQs3/gXOyqrf
yK+1hfxj/XKAKAyKHwtajrdnBBj8wn324XdNZ2cA2LlRD6NxboRoDILlR9u3NQMo
84/TacWQfJTR7mRbEVemgR4Yn+dpxz0lIL6cdwChHNt9VL3D02UO1vayeZn2clzh
k2yY5goKf3mop6YhcqCnOv9XWcYmDezj0e8pBB4nC5aHJiJFNR216ShcAeaqqW6I
OnWB5IBFHLj22OoIoFeZBBzKc7vS0Nop6uJxdmI9lYHdpz9Qm+yNBA5mZ2KFStAD
8Xis4mj/pVBnHW3YBObkHQ9niI3hoboEy+km7CnE8Ie8WTuxMQOnjj9xHYiqxCQP
vcHlXyfjMVtBV3HHvuJE9SIWubte2ARm8HrdQNfQ7XMS6tqDQDejE6LJk4Jg8+rc
hZ6v23HD9MW57TsP5PREqmKeiVcDRmi5Di2/AvN+QHEUlUACHjKZn59vCehKgZo0
20nRUkWql6AhfeHo9zN/ilx6IjDX4QoylFr7Xlasa3E/8cjWk2+edtlTicEqvW3V
zZzk+BTWdX196ONweIHypCOdxvsMdaX9m/nYJ8o6Y1FpiB6Tj2Zg8KZG1c8uAfUB
KW5m6Xs7CEf1rXQ6p3d0cvhWT4jtN3JkSOqBrwSQe9LseLT9kFYO4ZPeMKYBXYID
PiB3XIoUF68qL6KogcKaHTF5pOjo95v2TPAwFgN1+72T/VidKyujFPosT2mzAtla
/m+Wt45u5xMdWJfB0kU7G3ffz6A5BmuCpDSpjeH5B86G//4VBS2jA00QkhmTn0Lp
l/BZMuxAay4qoFi9trEEm/NRT8gEA11tU9aSA9m1EBabmCfpuX0DZoo6nHjqJYDj
LmwwCw83UlKJKdQnw6526uFHaaAgR+2PqPcBKshAHF6QaOZMYxaSN1Uw7usP8zNq
ECoVdh1nD/3Nhbr43yowlXXzLdA2PSSxuaLcZeuF6xsEwp0XKOVBg6zSVCn63Gxj
2JLsETjx1KFwmuqC4Bj8C3rUwP88YoX9vFfMs8FzcsaQSbCSZLkDGzToY3TgGv7O
96klQIGw6rg1+kCeHiROcAQ6UILNHlFqBLJaWQC1pfIj+FWl7oI3r9GX36vqS+7L
RRs09x0RxXbxRUHDDIluERmi4kl6a/l6sHBaOSZIZe4xNuw6cawKgA+js6aQzKho
I//fwnmggYtGo1xhHMDv6FwoXoZmQG20qlzffpdnfOE6wN7V2CueWcca8pdTMBLs
mBPVFmDdHSKv1t/J6K0vwzTDrR0/rBAFrTO9FSRaL6FenTgfwTcYtuDoTv5xNXTa
7K4VbaEEzoq7Lam5jecFar/ewTT92BHRVE++EJwDPkTe+Du47eKauZFqKFSwrNJ6
nkoHOroPYPwJFrf4ss6kD/KxOobgtEN/6jdkI9YXAhNdVuDbG6IAS7ilwcKB3z7U
2fEa8jmCvpHKPB5vRzzZE8Yn87y2/UJ7UHZLFUnyD0NckZCyuAW7a2ibrnJHGAAi
y0E9v/2KGlYF8nnhkubB507E0/oE+4/pldQmQr49pI1QlPgY2GdFAlM1DXOOiV9P
gUgbNTfjN7vFBKB8JlNE8L7HLmeji9JFeeLZS//tnCfDLL//Kne+Hv7mm2HByA9o
cOZ6kUApSJiaRrtjZ88TM1t3D9XZ/8xv0uD+En8Ok87RXW7A388+VVQTfnDRhy00
vrFPQm0f+GZuGMGlB6XFKWTp0+z+06mv1j3y5n9hOLs55LKgawWWaMa/uaKXGdft
27PnMuKA4pKEeG7LCOqXZZnhZkShamP60BhBP1bAASMWV0bU48LXXrEUtY+YThfV
N8Quxu0j4ejcHpSzWSbp98JD/0oxz9Z+BfwhEnv5jxItQJz+p4yYRkaZPv8MX+J7
x5bvH4WP46eY6d4T/5oux+mdH+x6dq1BXb6zIjuW6dQM7/f0kemv3Epf0HovHuiv
oVo91xpywPJE4xXyGXWV4gqvhMDtcn0zxi/ZqveifEXH4yYMKilu4i3kMPu0LsN0
EQVhuwAiG8zRvyTwxVF3CnV/VU98wudpVgUSi4tKEAHZUiO/vMkquOnBybIv/D6y
COYzDA0LqordU9zPA0saFiNlmTnigTteRkyLb9JqmbFGLmfTSuWudqMd5XEmqXn+
LSn9f6/ZOMitqKqfpExWw3qwZy36XmPA6TgX+lADgNvhhLGQcfI7z5CogdyKFiqm
jIlzkT8baxW46BNzSfbSm0mXJxp+szEW/biw5cyPB40mK041r446RDFL4nwM0O0M
koYEoQXpxNBMSGEPygQCCWlhd2aHHa1HU8oa3lsOo0SsOLAJA9xJpBouV4tLqgFq
zD8ec37Dwrm8rstuDMBpjLLeewzy+sb/1yXH30mMqyRs1amsVpMksJjrkuEHqPUZ
0Wr+tMSPmHofjX38ECO6xlAYIj77T5KASCEYhJS0c3SNenpP6lSgOYfAPYgSG9lM
A0yJlOOKFiFelbegn+secJ6HVx6vg/pB8HSw2jpTVEwPcCF+2KHA65xggr6isyZx
zVckGA+56fvrbgL1wS1GINFPzH8pniOE77gk7lwX1COEY0rrHyER4tKDZnmFs2vg
5fAMfYRS3olB7r3LoN/kNfxWyhjqaSOuOZoHRqAuz/8NB6ZGi9zEmOCBPl1O4Ycf
J+YH1qr3/OeGxJhgh91c14/ba7x7Cx53XYM1PJFnVDoSJ8Ba8a4H9K7xAQYKvCfA
5r1DDyRIXkctJoC41wq9gmYKhArELEVURzvxHpphqgOVTDW2FUueHfmZVyH0O2zI
QMr85wk3Tg85O1i8SkOy3dnxHsITm7rJ1fSt8zTJo/Wkhxyp+tM/+MkZB/HIeiCO
Py06hzTMCPgk8UIasdZnJYJionykofdWb4CaxQKDDYlmNp4YrbjkAeQ/sNwej1CA
JoBoJy9CGo00IAYZZMx54fzd/yywExaOAnx/TGN/rVFiDoIxCh/R9Wlzcht5kJTQ
jgVV7rxnY1CcUloStlHY3kdWy8Mf737X4a1UdI0sq1zm7RLB/eWKT/oY+HZOVG07
PGjnN/LSDPtivZtlBj/00TFmvxKbnkUq0s3xd0Pd/NzcPty7kXppSuUoTxmqiVmg
aX4ubEmFIB1wQMQT/5nUC3eJVQ4PZQB3aVubSKUxbI82I/HNNb+2i1NiAVQ3b/KV
NnliblmSHKE2GKrxlTTtnfum/OVuBB/MVZAmLd1UlBxt6mFRmQXqkram+bDGHazS
ncSEsCQ6vTeAPuaaRUgdeODTbhipEYthh6viD1JeHBcp++/DcCBgv4nytZAnNzXb
jwFysjggMMR/t5/AbZa+7ky6Xanq4x/tSsTlEbRE9EQzJ6uUdkHftIEqAtSDuHDo
hS2owVh5aFI0op5m/WTRN/3+FkPE0fsQdsBYDbRDBcgQm7VkWyXWSfliMOhZrpuU
VKc/rHJixyns76P5RqC2M/X4gQjB+rGb/Y17uLmzdNpN006ydb6Rksg2wnzLNLBq
tQh7fhm02uYfwVx5h2+zRhsdBlbf098DV3aoLWRntBWuDR2++0T3urZCij4b5GFa
0m90noRToC1tZobn+W23LSelhrt9YeYvOTJmreIeexSqiFrfbyF1UrRXQsUpgMoh
MA7NRQP9eSGe90pjSbNiYS3ZE7zYn97L5RSAjh0FGeQGnee/66WK6g9RKWoVuQY8
5rP7HVXY9IR3DckPAp1F9bath4+GAWrz+K/+2TSj9HqxYHWVuGsSHDortOyJ5aCf
ecNUcmobeIU7JEAURn5NKBNN70dK2rN3C5o1GO7A3n3lwCl3rdcxZeaOtyCMvTNa
5z2dL1xUUdqjhqgNUYn0Ike5Jlg3Wz++s+5BXE+CoYOBIbWWvW37OfFfr7S5cowc
eafu6wSQbPlO3l+OA+orLiivRvA6w2WM02hQZW+FlnxOQQ1ejRHrlu5o2pEeTKzy
GcC88tw3u7xLg+jvSuCZ+cln3fxOtIHMI4rbHofShBxi0ZuGc20IChhmxtL2b2QB
nZ/4oqMqeoMXkR3x+efJrWBpaurwm+dSbUt38YZKhS/3LW6YBCjpVIYw6JFAE6gm
Xrluu7ChGVAvKs8iqFtFcsThMC25F2aIEOOVRK3wE5VPL4wTElxvBFqXsgnQMThs
SKMSDnv4OICLNoN1SjZAodPawk5bn8D/MtgGt+ZLumUh1SxAmIe9qFX0xGenutTB
nJvG5xCPbNj/p1LjPg0P4rwWEX5lELOJgiTfjYh1ABbQogt6OBebK6L0TLKm20Xv
aKmWwtpi5GvqV+mYTY1KI3D7O/ZSW/aQpAgBjrNdyV8ehaLBXLG4FZ5tKtHME6LT
YsVnEd7VuBeF8jli3+G3Njx6END9+ylByjoy0akH4AfP/FwOAr//amFJxuPkwZsb
JOglLHWELWVxT9iu+lBoqmehxTwZzlyjw8r0wWrAFJfts4HIGFD6+5g3zqesjjSd
s2LvQcwI1VrJD4mlbTpxTzpQo8TL204bF9HAkgxdCWuPBzvW1KWkf/Z6mv8yySGe
qiOAVgtlHsuaqtQK4Jjzmg36fTwkXmWYsFRzCl+hn6QBRhrojFmDkc8CdbKGB1kl
WHNR2OlJFgh7HeIf4pSv8e+t/yxpXB/tFH3XRjn0GZ3N7m/XSWeZXd+hD8j01TRg
ut5808rmogY7L16ucDQxXpvWBA2K585MMKbba8Ys/2RsgQcDXyyxDyFavmYnn2KU
EiZFkjUgF2C8YEq3q4DGb82b0QrzxlF95l6Tc/eaSreQgRCnu02N4xGC/QvgBzmV
ELl5av/g2AtS5QrwBu/V9vBOnQSl0A6KDBfOGu3cMCyuXcKkqK2oLqF1GXsPrlvp
CCrgdlDVOEhaGqPDLA0X56jmJjhR80xUg4Stojbbm3PiRQMVe7jLC5qC2DKcuN7a
4uJbkZrq/wvbCxtNU1fy1GeDRkPGniX3d3ttkavlHKudVJe5NySkDzprFUzaAeIn
hhQbAXVe/fPN71nPse9t5MXhcO3nxuF1tzPG+PLAeZTyM6VVhOkMh6z8GazSQ0fM
pHT3G3dq+p7iqs/AlO0kyy223B1boz26cSGT8WBtHJ9ms+rwvErJuxP26ExP4WlJ
UpbLciQSfqzKm2EZIfhDT+MJmMT0alJpeixoV8DyrpRBVep7MWEH3sk3TMLKnniu
tz8utWbaHE1XuffByrRPz7Py34eggy9leA5BB18dj+oYnepksiBG8Mecth00IP/4
+ba9yyKOhQgiL1Wc1r0nDUF0JgcYDCEp+VkHMqXxAqo7kYW7llivXI3py0afHywq
Ml2FUgfbyjkWBIbYPCcX4E+m/CF9zzIdHpER3xs4pUp7hUs9OpvNDeb+i3zTpayV
DT/ETVjwCauqhfSsNwGIVoupSjFBEMYwYiQ+azw61riRwmF2bxMoKS2ihkVqmw2D
B8oIJuPAeAmIS/mwonuuEDEKndjnfDHRzMqXfAsYJv4h5JdDE2lqBSHgRywsnpL+
zlyTkHxtbVn7JE9ni60Yuj/4iaqzr3UDiHfcbO8Qu7qRzlm6y106BPlxM2+u4W86
0tIHeCQRwU5pdf+5Ufg3eBuj56/RzXuIH8rvUWHHvT1vogfm2X95YvsWIJlo7osT
z4P7PGCK3B5KEYm+TBtQxi9cZpk67IK723q0jikIlRvjoH7u2J2lf+03xVDOJSx+
6f9Di5yY7qJ99FqxBK6ypJPEGCJiDKlFIqU2Tjos4vJLJ3UQVfp090OoI9MGuKpS
GvklojIfl/khx4moVSGRQkC4aBeqWycEx0ufiaB6eenGaQmBP2irhexm25X4Esmw
eNoiJZ6v6P71iiR4QI4G+IqQBEXz0ec8lUk+Xt7jYnkqY7Mf8tzHaShj3paKE19x
IlNQ0diNhZ77vANvzFmCSItpHG44j4dY9TH6N/KzRYxPelHIcwIm9mhGIzLJYKCF
r2kX/Ow6obtQIGXfInBr7ouRgZBtf/Z54UMVjNfVl7/P005aDwcDlcPjgh6vAKCZ
emQuktEyEGKnv8PE8zYt+inShOXXr9cZi7265zge3SDiU3xtUDbXAAcrw7exojV2
cLOY47ZLfF6UIuGJbkhqPtEzHWbmqxbfOEUC0SAOJHh/kqHlmYb2ZAiyn/bXbIft
XbOO69HYl3j1eDWrIrKITU9Or6xbBgl6TqO1p/+4oEO90fReIkhkOY8rv4kOyBmK
SkSSa1ya9GviOMdHMEQZq1YzLz+fMnNRJFER9+0m1WRwY9QDeKKsZ4zpSPPTQb8g
4m3F2JloCHP01BU7Da0Noh/QUumVP6WNbvqferv6AM0m8NT9KpXjxxRUwiMDWY6U
eL3kNSJqCTGFlMdfZ/wuy2PRg/iFEJZqEYPGo3HNLTItZnTU+Mv83ROUAzNIou5h
m3r0+gHG7flIdOqETEEYqiEua9NUpSjhry5WxA81NM2UnoOnib2E0YMQRZa7maNz
xonL6WqjifYhZAiYfg/g3lSQUt4rmPgTT266Tgh6ondt2wBT7WCMBIB5QXdUoL7R
gIlV+qmRGdOl9DO54U7i+NALSLYkHgeYMLRjH3E9Z7r+uooW1AUdZH4xaHjn27T/
m9/nXI9ezOhWQwYpniCxeDwn3kbhUpFWGhX1wLSsvcJWg0KBdEd+MrYFbOSTi5Nb
gCLAFY/e7xvliXtATE/boltJKMcZckTSxgcYBMZcJ3sHCEtDpcuZR0sVGxF5Lg0f
Kh49WPB5W9e+AWoqQ1Qo64xnqbYsXpNzY6DQfQie1zzY+kpJZ7X350KAEgBhQZvW
7dOIfgT692FISQfARJNsrgVS9NOJ+KleBkc3k3wwOUjclAYzYLsaxsDg0Mjviahw
AbhtgKJOWQAbDJlqkGuySg8HwiG9oLdyeD0DS4lbCOkjpIVKC2q8c60hilyJ5EwK
KU1NynvZ4vtRNhAdIXHhBy+0DcjCkm0wJAVxKUbLbU9RVXG8rSWhjea77IiVbbsd
i9z9NwNJVjI7Aep8N8KI9iSAXXoLJFvdYFRydyLKhta35guxyNKqIqh8KyaIkJrP
94dlgjTv7Cy9qDtsOkorJ7MRAUASyRGuKgEaZEd8EQxgY2OdIY+sG6IL8+b82Awu
QPFdjp0qerr9ZVl5MOs++jbHpAgP+VaIyKMrSLr+dEF/7X8iPWhcBWjPdiSjhUKI
TcSdpQItKirTTXIqH0KFvxcG+9tP/Ewnb26GvGwuyzS4gIwMwPzm5jZL5/iEv4L0
/h18A/6Ekw2LrVP2u15vlPzu471fkrxYEdQTPmCEr0pUFrMhO+Eg1tuWCUYhV6If
qy9KGLVPU3bPp59vfAK5OO87pBpIVLEZB6HwpNl3z8j8aRyMEBNyrnwylbN6fpU3
jd7mIw6Ri5OzRGF0GzHFLvNALhbW95Ao1Ec1Y/PnzSEcSKKTj4pg+bMqTTlmeL8z
caYUYRwEWCrY3mt98QF5KbdaLY/RdkGTIcv0fdOEAgZjRAHdkcTicCKfBONJQKV4
q899VA0tZGhU/EQtDynsnQs1A+x0CC/SPGP2ZncyrcEKyXcOh3UKx57gBj5nAvCb
6+jDWMvEXnaIMPfvQRAGBGpp/QRdQq3ArvNk0ycBU/Oo0JRbxAkmNhO3OdybqqNt
YyvxEhmmWgSAeXPmWbdMm/v5ymjuBj0EngIlI0p+sQwl6AdP+WBSJ2afVuAIakKN
5USQhvUI7vBcglYHXCloj790GuxrC2r9blV6zm1NnY/1eX3W/CB+0LN0ahbiKTvB
vgvQI0J6t1KOTNyDzogjrKuZZ/TFr29+tQ0oOPQg2gZw8S3OcH38nLn7ZgCDrpPq
dkEhvwdFs8FdtEmBGhmdfa6Uj8yFdrtF6hcdWIMNORZ6pgQkkOa9lOnGP0hK71Hc
dDAkpAR8pl5PmVWyZFeEiZmFrKoifgl6WB8g9P2bNkTZ26c60nSsR1rlGom7b1QE
F3405PKxRpRDGtrFvCudWmGhEihA8RuCdBSncVteGeNXa+4is3qaJ6F706wSnfM/
kyI0kXkJWQAaMMdE5gMdE9fopmmXRB3pu8T8caFrNZ0slFBAFeqrTteJIBUFvDKa
wQVoGe7KRGN/33/7wiyJ2+yO5ofLjJJMs+7fsbg4TSpUpcBIHe4YkwvCmQ3H7/3r
fjgtougmY05JJWoVzu0JPUjQgASQfjk0jEKSrC3FDu/M9cTLcoJNC3G4ITPDYDlM
XNjlV+peB0U83UYb8GEVMrSFK74KH3skBYFRmyhHYqjrXUL1n50LRlLRCdRQce1X
uD7w/zAkEJlhqZWfoiU8Q4H1qHNCAZbGMUWZj73INVpEo52D4uz2pl1FL8K70GlG
hzEgTD+e6BqKK0JB/DTYQPbQqPZ3iScpygkF14011Ml5XkSPFHO7umtE1kLSdgDW
Nd5sjJChP/xcE0GN8ndWx/bFRxJF0BEb0p3D+nDfSwjdDy8oU6aTHpIjYuL3f11Y
hlAfbzDieX2NOSAOPS4q/NX69lkBQbIsGbEDf+rhxRSHbJvYByMFMYeOIZCHpzES
1dH/Oz3r0vTDDhnn3Zg6xHoCqDNQM482BO76q6XZhdtbj9BiHVZdqMdQH48mikc5
YDV4OH8uFbXsuatYQ6IfAxp3OSrQd7+GMV8LfY+BXmHibyTBmJutEb7MlSsowUqw
ciO65/QWW9iDsqulWLujJFvJr/bYLO0rvTG2vOf7ZMLdDiBBQkchy7htd8JHAJZM
bmtA928lRAYSndcfLc26A3yb4ywllNoQTcqYIMk2dnmSuJ2G1k4TUaryct3eaOAk
unLVpmc7GW8kbV5FjrTGfmZuSCszE+ua0pOjxBrz4srqpKdmRJYea3Ae7prVIKRK
r8fCnKLPBa1555lyQa87tqgtA+te4EbEEjPmN9x6dx4H8h1w2CRxxUhDlkYJko3a
ecsv9+y7uHoREEy4LX8yi+04XbaWdmC76TVDnlukavF6G2DXQHis7SKjNJ0tPexx
VCum45aYxjNdR3xbM3rv89V7lKXZOPjvKT1VBIDMYQGISTuQOIaG7qcDdjRM7boJ
pfjkV03/95Tj1GixcXUh9CMDKUoPIlKj0POzmNW4MBPHQqj36acINlM82qakFfNz
rKU3Mrp61wb61SbaYhiOlEqsS9gKB94KlRsEPHMSZQ1ZdiX2RS3AA6ftS4vAdT+B
dNhJbBJfbhXREyHOfjgU+QBB9a35n+QecT1cFCaA1IjXE0M7kBkkLEw2yoHVAX2C
Y3H4Ya/K08oD2M6gTINOWthWDEL+gEJpIMAh0eCPGpsivnvueqRiwPdDRrTiA2RG
u6E/wIO+yNlF2SzrbuOJ+MsZWv0lqABGSkRVSeHjWFh4LA0IuvaSXEg0JEcvo1WA
lMeqlj9kLHNfTvCpByl27RrPzuv9c097Fwevl5LzHsIkZztiLjZeU3oNSJffoaFS
2krpdJPbgn5h5o1zXeer/ga84Yy885B4xGd7Tmok+OTjTi0u31JjGRFsC+0+YnHi
FrDftdtlSpM/NsDYpmh2cEQBwHK8Q8bhW7I3TxfR/USsO5/co8FM/FV8JhveWCtD
ApZzu+cvKaOnUxZCTfD42kGq5lSUQxGKrTTpd96hpzWk+n4TCJ0lPdOOEJJuMYGK
DcH5UPXSbFIWMp+y2mTJs3lTQM1XEcBrdGovK4Q0I2Ul+iA/Ib0Fk0YCyliLKOcU
e2VaFxVCLNFn0zhuT2BrpwBcxUlpRWWV73cXrelfweh8kVOGAwGiNhh5zdUta/Vo
rxFlTIVuYI5HndJi8BtCLW5HCuSW+sM7+mGRphVDoNZWQknd0aVmYYkJn1opdLcP
2yRCqWD4q15hxKMOoQdNjfPZylUq28XuqyJ9vIzVW+4hOaOK1QwDe7Z2Zvak26b/
KBicgXMr5Gf6rY3UX0p+iX91QXBWnwYOl6AUGaMdIN471YLscVXsgVCa1VoXlqwk
4HKprn//CrmN975M5Hs46GslYF+cuMuuFOsZr2d4dXJyLULDn1+CTtRqyRb7FOt2
h3WfP0ccz1pH9nWQVt5XY7Axcr8W/MJiHP5dV6GxYuCGCrnRCOamirbIXv7wNGrg
64IysqJTJfkWcC4CEX1Vq+TUO6IM3JJEF1kjG4ZKIBcJGE3xJIPELAnA1zDaMoH5
Xi/BWykRkFYiZpVqai1Fd85loZOeTaPwNIEGnvi129AuxH2UKJDGJa0VM3LMH+ba
rU/5iX1F0/Apy+G7cs//rG+e/9eW8JeVa6Dyv2wnWMj4qTHDkxTmg8TzbhjtlQkH
+xa5CZIFeYZITfPB/VYbyicirar61B4/uN3BUZDoCTk92qVMsVXcdrPv0dbG0NSg
vNZgMY/XJFrcsV2mCab4xp4Gm2fDWH7cd7Es3E9inQLv10zvJGITb23/Gn48GSIv
NBoyz4F0QgnD3Mej10sNTAfn2j2/A7GfW3Sc3WUfmjWQEk2tcJ6PKDmSbQ/Sw2k8
Z66LHujv+gKMsDYU5ljJPYwS6opoyA5/lAySvVrimUBkAW8d2y2PIBLwtJSHt4VM
yuvCSKvH6eiSmGekRsZG0VuWNcZLLvQ4VVU4VWdcYB3aUxFHOsIB5JPF5KueLgwM
rFDiaunjVCpGKqUYcg2XaJ0gBr2Iv++39OC4WZ2AZN45VUOiyPDJmiDEAA9kmvyr
lxGb/I59C2Aj8XJ1vzDkOqfNvIlhaQdw+6Ut9YaloH+5M4PXYrvWdL3bcb7mSjAU
OxNc8jN935h5LCb2arLu2xwhf5wKkOFnM1SVmIbUrLpAYElBCl66AlkZ9UeM9yTW
N5v4U/DnT0UA7N+XnJE6UyojYXw64JSR5fJtnbMAyedR2mNaY1UtpIZf+SqAHfHp
0M6uxTad55yugawm8v9BpogPob1mLrYzK9wTKdFkI5RIuAYe/Rtg4V6deiPqGO/b
I9HWv1/GynCDEhxuHYW1j8hx8tWrauQyqvDVItVgYZNuZ8Y4fj6jyrhAHpmS/8X4
ZqDAtTczordErxMffJUFJ7knvEoeX9bSbcnDeY9pSKXq0nzxEn57pVYnVVCbv7kl
+SPJQ4z9MlV4tNJCKUA/8oVV619MksYlqvNFYxXdyCDYFPHac+WjaFXvgg5Ud+h6
wcKx+YanbjETJ+yTjyjqn0BnsAArdDbxr/cZTzJ6NOMklPd2qyYT4eRX9vs+DdTW
89dMBWY7ZyKwqZ5MuMwy0eu1pqgrO6dP2zosKzmvlt4Dcx579USWOAbvtpVuxehT
UGCeJ2cki/Zmf87FS//Eri1IcCnjDiDhMhpuphv7shku5YS5AZPcnOtBnbUYh8pD
YdooB9timiOGZZL0UWaoGmILXAsiDpnDsLvX4LGrSpHvyXlF2kMxv/2pw5/Fa1LC
wRPKDGRAVYXpWQZK/41vSDIDncKztf0umrnd7cGbaPmUwzLwrh7vWeqF/S8UdeF+
+5iFbQvelcjIgmHL1H7GEkloFQPk1eNCVdI64k5+4L6irOKtZD73q+tn2qz2LANN
qM2NzkfUQRz+Rb9BQErnhhR5Diwh/TP6G2T43mudneyKs2iddshYQcmdLVw/yFnv
hppE6FQSrj9MAMNk3BLQHRB5a4qTVBrLR495OmvqQQCfne85R2DX1acT8tOgX+kM
zXHYa43PqFYhF/iGi+Hw8cTK2rM//UbreWlpg88RwNWNPUq1QjRKUDoUcTwBdnoK
JRQqdCFxPcKgS8pi4TMTJpen+J7+j0vbklnbq3N7s6Uc0eRepe+06sgBat9UdyzP
q3b3BeSIWBczEuSlHwyEBilkg263SxRyBsrBbmFjgQmfoWz3tYhgFaN00C6JG3xD
MGNY+y4Al1wl7mtCZUnqc8PBUa9Ipiekuh91EmFyZWlJhxhXN1YZ1ubi49vkY2SD
EClH/LZM4w0mQ7wSEjhg3FDVytWFwZNBDCU079DoJZZgPuuMy8HT/YsM8vNVNIaK
x+dLSkpAOt8cGVhqVl91O+Uy95h2sG2hmls+Tnc48/j1e75TngEavHnnuY9lV4vd
oqnQRNip3W+8fhdhH5RiRLUohlG5r9Ws6W6X3EWvaN7m+U/BSFHmWFpXzPZpAH95
grZM1OjU044U/rlmzOEHbIiuLwxhdaNGI0nD+3HvAMokQd7GB0D5pXJ18VeptddG
bWYeicz4dOIlXIsdztbj/P81DiHaBY0IdaAT5hIfYuJCPAqHlM3ZRId8PZun/Kno
bsC7Kn04ZBTD6FhdEmtVyWOX03PX5UzYpa5dozMaUUyorx8Qon9KtNjhFD0eVTa3
vcFjzwAGpO38DZLTREQLp/uGRKQ5xWE3YaBGaHpH0TXDUsA0c2AYk4MAoF3komap
d2oj7acnuB5uU+gt1EPj5offaYlgfDKGRUHXr5AoS4c6MY4FgaVrmbBAUy998WHR
DINErwqsHg0OgF0RmKPuJ+8SuIb9kLk6ELBtBGzKaxMndmtBYk5DQCSEmmh0CZMk
KwBEPJsevrDz3Cjhw0awR4AKGr3sajGEvKR1BZyMf9jxF/EZJt0WoFJWQRtS2SvX
GAv20+3lGKbGy2RZ/gdS3EsGbAmQdmDHpa15Bwv/pLNgDU3A6/d6h65COJKc9evA
0Hdogpzf2lEOeiW0zxbFvNIdgHZhkmGytBM4Tr1/bL9DSHL3w23b0ejHS6WUhae5
jlvzsSUevGFCIyoRaJtF2M1NYhPSq0Gz51G9KIm5scxNyBB0yf0bJSAauiUPyACv
tnRgOVPrnesaumOmZ8RYhmCDxfnIPRiL2k4KFnUTNU6/l6L8MtlaUXKYw1/NZ9eN
86Vnrx4GP5fqn9ieuhTrH5HtnaX6jdsRF3TYkiqjGl1b1/YysCfAP48yjHI9xQjg
hLZjpFv2PclIHVh/jmKV5ToX6Tc4ab6n7ZA2iJGN9A1G5jauIuOxmLVYjYW6o8sS
hY/laoYJ5Trzwod5oChoFdWv3uCznf9yQga1hIsnyCm2bp3OTkC3E1Tt0jhGPLXA
ka3VcVGCJdwOcO1Z6rzvv56WTIQwOZzlv2L1Jc6D8LMURET27nzGnnYOSHAk1dBt
6zkSoY1DnHI24v0rLTqndR/CLCbmVaIbgHdmDVl5P+vUmPTxYl0IZxEhhEstKq7w
4RNFZyLaVfiLPwCK8ObIpew7mSNt/Iih73MPEQqUbtetuL03wGdaQ6FlFdbdUsna
/3fFtLVx3F70s9RlrcV+OTT7qWw8GdzAP7iPDTUdyzmizDv9vUJC8UBCdWIrM49n
GBND7VfYUWOKKG44+b9T8sANU3hOobdl4QIBMJWZvTdwQmmpPZKY4znYdC0vA326
RBEkJFucXDBwQsnLCP5zqnRd1YbIttcuUNwWOdai6ioHxKDSqOZjvUd2DmhxJ2ry
4l4eH+paFlyqX1WsHEqL43E7cpdhi1lGiQZf9cpzBSZkcrWf971KBq4YIqkW36UC
Cf54HmLh4B19eu9urp3xPYsYUyFxWwJAG0xDNbpMfD9hSyslxmxr2ydwI29plCG2
XM6YxQZVBwLZRSe+bLuMXkTBaAfeyyqEbzibqrPcCDLWC47dOOsMzsiHM9/VSxR4
T7lrcaYneIyjqnVcz8WUWZJSEflpboJBF6j2MSqAn71aNkrI27if1/DeO0ZHjB4N
Xf8cyzhKhqV42+hJfVYqAU2AL0b2VWZ86kf1l5hGVLpgDdVwr7RSr+mKGrYYK3eM
rwANchZx66NCN8S5GXfJqtPWX4JrohrrTXYJUzbUB1jH1TGxUpNVJud++9C8oOzq
VMLwP5kIfT2AVA83m+VjIQOFhk1LrayMvM8bQqawJOf9HBxPM66vtUOL/pQOEWQw
wRLrBYx8sypu215bkCXgf18Fqo8UdNZMQ6acfKe3irV0bmYb11/5qpfnMI8FcvtB
Yfd2TTdFG4w4OzzkOOY7gl5GuOE3kvL86kUgtxtoVKnEPwnxO9EBo92p5x+0xJJV
6hiUqPZ0i3/KaObM8rZeIAWp2WIAQvDRErPI7xsJ44N29+qQGOzpzxxeeSkbsQDZ
0BEhedsBnzggQqXZY0ADTJL4KA+cOT27FUoDhACPByJW7rG5F3XCNSbfDpLMbNy1
Spay2lL6E5K/0E6y6cv3j6fX/GvU/j0wFb9pT/W0xXCxixtccWfgHNCv23jUl+yS
fYi99IUv6Yj3BmU5UvEC5L2kAwvof8gfgaFjOS27b1sYItNTXFhdBujaX5dmmiwG
8LUkp7Ama1vwqbaIXflGniqYKC7JRxJ8m9sKmJOPexCQEf4UvUWK7AcaUvmfg9dn
y45/yijNNd2y4OSr3OwJ438iMZ0jgHHgd6hwuQEJqV1+k4GuHN3B68gX2jJ15h8x
JhaPt76yjz5eB63Xn7ldKMh8Mn9/cbxP6ex99fZWIzPKYA83yvIee+XJmMvwdW68
nG8986Cp4dwzs5ZJf/XLiPpbCFChBf/Y7GESyiZhs2b5E+9gr47P/s+W7oCcWNXX
9ULB+cY67bG76Mhg/5Bsbo7G9nOi6P8RxPLA0ugwxPrX3D6kUdvLMPx7a16qVmUT
lVojGdC/cMIbM8ZlqxYfgSJOigmHEThS9/nxoAke01f4hmd9iHphpNe5HxHitbgp
k4A5AzWkHsAiMYk9eITZ9gnfU0jIEBY8m9gQ2c4JNmkhOHSAf3WmWTTSiSrpdP0U
MXsnISYfxXw3hRw/zmURmvd9baTS16QFedPIgdXUuMj6hkb8YJAE21p8PV5FKGSC
RGrZ/kVtlq5G/EbKtJM7XHfauNQv+1r5Y2PY9z3++R3ePvY/5fuGU8uucBm2PU3u
9d6cf74820pkeFBuGk4dJfOH8RjQ631QGKuEWXr5slEGXciexBDJCzviNynZIDfj
dpOJWu93OFPcwf9NLZk4Jm0Sg7im7qS1kapEewUWl7mv7POwxsrfjFTdVJJqW8in
/srqKfobUm54KYgF0EY5w/FfWCccRimUkzMMaDdFR5bQE7W/giYlB2TwtgCizONA
SEt+vNs1cRJTgkJKxWYWdLfknwzPODmBonaJ9K6wd34/wZvOGClB9D/v0SjBAqDi
xRTltkaICjCBkEKdRZYTHYWuMdH1SF4Zrq7lCEK7XVaB2lzWy/VxhiPMZHKkCm3b
oW7/F682v2LuyZ9rAwUXcWCcTuoUpOb7Djiryr9t9fTW3/cH2oEOQ2RutaM0y5g2
+r306TlGsCCtpHTf7HL9v8NEsqrpVnJuyoDRl2yQ/4+yCENxoq4nyBJ2r0YZxXlH
qFQS05ADzaSFmu3Pi/wlESb2D+GP7hU+s/mH16zvHBY5Khgwv+z+OFKGG+w2MHxe
fekHzEjn0g48Q8MS4WmPW18zyIDlsz8cWJzCC+cXk2RyecdozAxeQ8W2PRIlipsv
fbJyHRS1CQXnLaIM1mTSq6xM2AGsT2fm1hMsXjDcFGyzKwXYXfif94npqNeXQ8+d
iSetbsn+DWtsGVAs961BXWlpd43HynXpKhh69zmdKDPCx94M1kHAI/ZnJZ9SNj0x
45LLWrZ8mxI28psND9tCTn7ZjEYUb170aAAP8gNgwkcKlNKXHuwbvThQZb1+12np
DFsrcN5tbSwkJlENWKT1bzQe86qX3QCYaZBITFPuudNqmLZm3NPR/eUoI2+Y2Xaa
NX/ZBAR+6xHxoGJBNChNnAfzbgTc2SSh+vpcTvV41bLnXw96dQp8I9fIHht1tCBs
YekuOiGOoHtkHoBaa53A9c0Nfsjv77FxIFK+iLoJVuiDQE61RtCczSSTf67k36K3
dZaGgbzHIfbui19jtHIel+xkf83jpOP0Saim20nNS96VzufoLDYPTtscWsFH6CbY
sF46LZ1tX0q8TVkyz95bKXIXjZVTt/6DGgJxDJ++WSH3BtGABzadIxMpfUExsYK5
EJanww+TtHeAON28AQ3Hew9iGXgfDHOLJSWUxPxqQkfToCg0rIpBxdS4EAO+qiO8
S3OC5Hn3cru0Sk9apI3d+s3ogoWbF/IiJEe457WMjpUxaGQhfAWvCy4R1ptLDddU
qzPKd8sO3Dptn7j8KhG+Kp9JCcqouILhHAY1G5QXc3AzTxJOzibR4E0F/VZWCk/K
jhkV8ciw05kaU6Xp62BDm7pk4p05DWNHXHEgBU2BowUCX8O/xcMk27OX5lTklbQE
63h09J0Y6HBQBVOmFXzT7OZM6FOgLhfV28zMmGJgCj+TWYPTnbA4IMm+GgLq/IH7
Pn+qHnqbPVrZA8DGGR11pMajQVXsAP9u5f1IbmKcyyE8iwvBpBtE9hMmxN6QGmqT
+ylSSUmwZjIcICd8+hSlNShWR65T4dilGuTayMpq5o9wwAPkAJA3kAc4pqYFZWJG
rL/UNweyDWLHU2ycVXG4leY15+Jc5uwA82xhpCxi0VBo3Px+rEMYypNjK8+69HV8
2tvP/4QbICvZDxH1PNrDZ0AuTJo0n+JjTd5rlaYvQhgjILgKxlBsbiEpklpUgzeL
s48yM4Nl32/RybYN0pm6IQ3zd1yy8hcYU3txTsjxSlNBEtS35pmFNkFCwWEmG/3S
YXhyrfdSKdj0rEuNPYw36C4Roe2ymRmXe4ljghmAmwrmgGzYiQSLwIAq+bv1mGUI
Y/vdwkOE82sMmxDLNsy3KyeFEHi3OiqO4I0XpYLmp8Kg/NikP2lYtyShf0j3OZV4
DeSwCIwd3TBUyfDXOIJNaJPBEz5zWb3vNZHod2t3LVayPoYXm/Sqw3t6Oz3SwgT3
kkoAla5mOGT65ZMAgI1gPtGuaxapFLBGL75a6782HtPTJLh4JBFiEAY/IJ3uQHSi
Ozqx1dYQdNDkHQcAD07jjROL+zlMrszQPAFEm1K045NmzzFzqd+vXY8dlLgPXFQx
gTLuKVXESmT1cIS9dUX6jlPrMdfoS4jGhz92lDtZ6uNG29r4pJbPtkW4w9tmpY4f
t7/nmKEub9JGT51VguLVFibsMBBKc0ObmLrYIQkI4n8fKvxazd6PsY7/BoQ80/FW
mHWshEzN/5QlvAZNVxN2hAfenQCdJ40Cu16PwV4RWXUH4PpQ5uLOXA5Tghaw9dlz
XKfjISy6Ruv9BMrFvCK6OyH++0XSbJLTcvRtETcgk/RXCThEQObN7bWyxlNXGv8h
Q5xVNWoeO08+NmtiSNHr9+Db6oson50m899t/t0PAY1w4+/d16RQvmXWRvIXBikW
1nuROwFYY9CrKfV0vqZBmouwgFf+SmGEV6OYln401zACS/o3xJszl4q70w9oQ496
YH4WeZDCg2S0j/9YZ+vrKx9I623hjgmBxKlfe+sDG3h2aEG5wlngikUJsnCVZWF5
r08zqx6KXVsQKle9HTDB1Wc/SWXpGCpYNL2Veq/d/FEycHw1TGj8DG3/IeiCpn1a
SBq/KjzSHRFhu0PTHEsklsczZdflM0lWsiR1Ye+9icjCjr4JQnHR7ZvMCqQ7HFP+
BqFkWXT6EhBuaIqTGekmiFEndM53Xy8dr3uBSDUwCeS0nSUaEc+N6V0/kM6nc/2s
Yymx8EO+t7YvM0c2bSv+hkhbtDLir3yCCm7JsIfiKYU/9T4bz2DNEvKxIC3XIrPX
mWiiOEoY9PoCWBmi1QZ8O0IH/1+LV22KyCsp3ZJslUa36m7AsTe9zeJTEoY7ijXv
oQX02ay5ij21gSYWDnB/leVZuitTkrjjmUH4zD7gqG72PMbWpFSK+aeRy6pL/c0U
gPQS2CcAIID56iGvd74lecnR7pCxwHTkzGzP4wwmxbPZMfFep5gV6TLsOlorh1eH
LY7yja2RiM2cxVTGjasGhfHT/kYqmy7WjjFgsWPypVHZPLFyEAHHp/0NF6J5mycw
0XBQDH5tPrWzTjzrotykKvTwGJiRQ3s1+Jdny07VBGhmnlNGpKwM7B0/NBIJN+qZ
jVwHoC6waZHFXkUSMrV25JARouA+E/EuogsLOD7d68WyHaB9oPeL6pryGULsJLVt
dA+EwYu3nqeZmcobzZ8jCJv9slAst9iIBYJcHzWWok0IRc6MqGaotLGwfcGXkMpl
8X9hELOKU3ue5jQ4ZdgaTaxXK06dDr0F7BI3Wvn77IftvZvwEDslDqQak9P2QstT
b+Oifpdzo8nl09NzGshudpVHd67NMvja6TllLRlxYtXZD8TmMCCkBAufD37d2+xj
cK1F5+fH8JjAq+Ua5Ld5HZWYxWxwZiZ5sSPTYlVtkxvnos9YViNl8dJkmQgatUHg
63ikilMQ/6e6RsdaQ61TaO+h4cf5lRJUWffoZ+xCs6ZnepXo3n4GmYDTgtbbeN4x
tCg33IPJn3Q33YkaQji4VszaSRKzQZ0lv+C6UvkmGV0N2QU57e61TvuTXvvqt5x3
8K7B60QMznoOxLZPqU6fN5QTiaolCzA3rnEOl/XmLY6NCL1HgIc5HcWUiLaOBoq6
Py0aQ1D7gRoRHXjg45T3QuIHRLoXVpmSmkNqI/tjtkD1F+0duVjVE3c6GesEVV6H
lo0ePmcMhsYuglLGPoz3fJrCi6gEpRbVsjUUya7GkzgjWovZtuUJ8IE6G2Ypys1b
YmqfeUlnRBuww1DxowSWUnJv/j7sfJjGjoXNlZ0VRa9+OcImwzJyssluxl71lre8
aeSedij5aTGnEwHRxQO7zYcNU0AmHi1ZXVsLxWubnXnFqOYSlfi4gTtFVYGhao0S
BE53GxJCxM29JL+nKG04Dja4vjsucSlPkJzi8m1F0fZFB/0kl3BfaVfJ0B8ayR4P
0AXmSk4TryDZSBw3rLU4gGNuEFSYiPvMfNorMyUBERFIDyzJSE2OYCxzQKsnT5Jj
6bJaPg2auduaIB+A6AtyZzz9p+TZWEZyoT3f9zOxXf8x2KOda7p880MTWbMKJIBE
frwTTfYkWUYL2kr7ZAL1HI/pCHU/kAli7fbyrORinWViPjgyqnQJQhAeCVL1S6JX
vD2DBlK10Y5ouNFPTAah5lJn3FDKmpAILAXB0LsAvzpOnAjVRkTKCeDahH3+JIyy
YAcOwGAAXMa2K5jM4HztbffIOGEZ/tEeowyx6ZrTieyr406ghufiLtK/59TnTeDi
+a3WuhtQfxyWaGXWlfGB5B4rZTxmUEL4NxPoUArkbIVkZH9JfvF92f+2HpY3Z6c/
KVPorM8KsiQ8nYJ1pBqQOecISJtSInmAv2tCnJCkExbz3hXVZy2TYi0wadeM1gde
lU+HEoBle6UuE736TADDapqAi7N6Tx7mFhf12dZP7Rw4ROPhZcYP5c33U9XqLi7c
vjadY0oQgdd66PYHCue02alBF14qf325cqpzQ3e0Uv/qIETskcJIRnKvCQLkGcTD
XxSeQod18vT9pfKyoa2JQb9foGCVw+WlEBgQkqGPyx5PZW7L537a8SrhsyFOennr
KkWOnz0//1EwbHpjmqEv9EF1NzRKpbmugLl86jmzYLtfiivqHH+lIkTtEFZ+w6og
As2gbEFOU9LHHIdtryGyoHgH376BWqr0OSfoVkY4kA/7IL46i5ZdrBrj8yaUfl7g
kKBAEYoNONTA5cEQueABnWWg7CK9FsXolRXZvMPOSrqZq9KWg+PPuqDKeFpBPuOX
RvOUI4Mzsb9UezjT78KBSB8lMDVe8r0HGscrFKMZ3CKhReNS5Xazwi/7+Elgw4rR
mS72F9ocKwZReLDRbYVfYMY3nrMvKI8qBpEJl6Q3stq6AR/gcIncq198ZGkouOhj
Xj9bAwSYjs6tkCaUc695GTWmOcrsYUYKOM7Rfm09fit2L8pr1WxatNNFGRd5+c5E
WiON+0HrHORJZq+AJa0+qvY12FU9UqCpbZi02UMddbyU2T6z46cx5Z3JgVvsoyrc
LNcxfSRZSsXO4vl9qslk6jahGCKbFfyIMrob3IOTvXxuwCYedant76KW1tzOZiv1
cFi5CFf0M7OuXl+PC6vlCsvxyKHcHnNe479nvRjQG1FMU3gIRM/td3mfdnN7rAky
pEK+XT8g36bInaoc56ZkEedr65ukPfxDqOZ/eHUbOkjfIO8swjaAva2FiOYTgPXZ
LHXHnT2ND9IJhMU0sk6EtVMVeo9h8fqPqLMdF/Ax0asMlve236Dtak3j4XQSsqHt
V7+icD1kCfv7XUpxH+4b8ptGAibjrHNF49ioFI7xwZPZj2XZyzSpBxFcYC8qgAFb
F2dL7HgejVhWvSZwykNCfBVVkStTJbwpqcLYuWT+KEz20Ld2S6EL3GY3H1s910dI
J5bIw/T06oZmRxiDEw/RrZdOWrY4bK99s5Mxdlc9/rToDvON2PULvjf+oegkmdRw
YDUg5TDofBBjj0fAyxs3VFaeXA1z6y/h4zmc7PzvLFCWj1ShphiO1RgZXHE0uCP0
OpXdR8Yd+ia1GBM8OoMLqvIfPO6Ow4a5TLYDqWUYKxNcPKRwJUZ+ej5e9LLpLI/O
cK8TSEbB6agmHFCvpkp+Oz8QUAI20C5iNitUhKn1qVBB6qeWfBD25kJeS+eQCSjF
I0Q8UxpCdEwUQgYduS4BvJz3Ejta5OtSF8xYyJtolRPptofolQ/t1lNSHFGY/xOA
2CEXETWt8A0Iw1kRMWOFyKWWfGSWkgtv72BYTM4o+cr4EVKB8RkXrBWyYv2AWGQw
rbi9xqaejYZIOwvGmo79kCdpitiaXMGetK1SjenLL58S/fj7qz8fWVNUqDY2WooT
6FGvmxezFevcWnU6dZLokuP67W2q1OEKt56+5gs1pdtzPPT7TgXksEMptkQxXlqB
RRUfiR2HlK+FmgGvWqSNuDEiqe/WPAVMf0/6Ir2z27oYehHwY7iORzyKnz6bE0Rj
GZbfFPPww0EzufknWE7FkEXp3DEg7WDLUPKzHD0i5KLJ9nqdCINwQNGw5Omt6Xgl
RBMRdhwvij1NSvjNPQIWE9rvy3sCMyQPgvkzG9mnY6vRqBTZBNXahUVaTR2wQ0FZ
3vQxcsShNOZjya3SyC/KnAmcQ2eYYdOi9et/k6mvzq+LsUsmovsxro2CIYygadLU
y1KkLqBpJjzFJdx2F7FWdccY9uVims/oV5GI6XKNECVDf3SendTwditHc++GPipk
T9ITRCh1z13vo0XUDVJwQ26WmsC1ZaHfKXQ4i5zTJ/N5C9QDmnz2rPhYMHgtlDhd
u1Fbm4Nyvb7yHvCwOj04suX7BLj1nKwoMeO6JFVoM7mOj1GLitfoZoCLCBXMsP8v
lyVV+kfbdBirkcMGw2zenDVzt1oVVLLrxrPlopEcj5QuRwO+5os586Taf7Qp+RBD
dTT3mCGtFgwmfREh1DmIwnzGLAHsoVE+jxMkzJGZd8C0lEu/Khb3j5OWcopuzNUU
D2OIBONe/XPO3Wd4sZaXkD3azxbZjXOVJvW/OZuqboaHtjxGzo5wx2Wach9a4zsa
iycTmLcpZgoeu2UY/MSprblJnPBzvNrysfempBmdBsyD+y71fWp82rvnBbI9cjVG
eKQGBNOHppn/FriHBwElLdtg/D6Gs3fspCi73MqRXYOfuqjihOHNKHkzKvy64yQj
BnFph4CWLX7UG/iPvS5BaPEz1ZK2ahT5LqC98XjbTLjo/W3Au03iSZKSFVN/6CJx
W1jD8XwR4aCXmlElFFDr08Uf7YkjQZMrG5srZAouEsc6wGyVwb0btobclbYJH88n
3g1NvkpLf7VV7hJHe6JLovziRlmDeB4TDXyYSxX0j/qSoMRgGPGZR5fEhuBKabiI
oaWMid08Y1w7wYcKZtQgGBM/LxqFfMX5ViGB5Nt9CST0GyiW15v5irioMAvwBR8U
L2uOUWhphdaQgKHuyn3Og2nFAsPXIm/ddpWksA0yhrnlL6T3DdoU1+/oRHoZ7spw
5Xq9j3w82cstK0nSGub2tl9WBIUZJGXICl+wOM0RnXMQ30oKPu+FDnEWp8ahv1lU
BeRO9FEZzwdxXQcHv8RQ7n1J7lFBOSHVFDRVjZOw+JKWRCpw7quOhGGgV0JcJ5kZ
BfLLqbEgFu2dUxdUYPH7OWCM+EUua9qR0P+fSzi9u7ibi4COymAUqGvjY14iIyn9
pxjSY2EUVB/NRqnSOfywu3UW3tmCdmnLPvYI9SZSyYaArZXZz8N2Zj9HXTA2KPvv
UqwgmxaFO1ufajkWOAO4WGURuS6eCA/wzQkOpkEQ++hcfwHntpZbM9A1hQsfq8ml
0t4dXctPBhLmCZyKTyGKJtftKPK74CRnjmIf/m+8HczsQ1PRLi9PTthdo4c0g8ih
yaqSIStoccYbanPTC3pSKgozarSk4EnnyeOrF0A/5mmVxy79YPmK5JedD1IJOpxL
YUtVII2bA2qjU3QnQqK67TFEeD0R/PUGaXiD9iEsrNIFkgV1pXrNVUTJcpD5a/V9
m64EGKfxP/slARfzVlNWp3YeqKR1cxEN4r203ap4X9XT8n1FarImXPbDh8QQdanm
WJ3D8LZ2tFdJY4xyN37F/J4i5JJdbLqk03AxU1giJ66mUMwGiN0R5OtT+WHLrDNM
g+yKeupaSt4PSCmjRSTTkohYKWDc1aYnPdI2AhQZQr5DT2FPmX43i1PaEWzvz0bx
VY+n51AQZ9TcGARZYmaxLR2EZc3wOUUjdouwmney1YGCJxTGpaP5G/GAQPp7+wVD
gWCNHJVfdI5EfzQyJUJqaE734zWUbNlilvZ8f273ULwxboEa+wLmPpXxSjdk5ql0
QDzo/QS1UD2h+Kh2YzD2pRU3nulVVow4ujxK8wDpdn/Og2FXxNKqRKEGeFl8VUr+
VdCTif4bZncVew36oNyiOg4qrABl1DfK/7OsBuszT6imVDEXGnakZl2MwfBVDLcq
daJ23dIs91tG8gI4LFj14QJSFwX/ooz5kNEjpHk6f1DTpKKR3JBhDzf1wSE9JQ5t
0W9aO+vxrrfunFCXMJzJQYGKjavSzig5XOMdne5x6FGE6aTo5oM0fo6yUiGiD7mN
lun8mh9rHQG9ieK2jH5Vprc675klNx9y8PQxvu+Om3wN7N14PlTSt1xjzVgOQg36
9w57fE7mWqPddpCTGdi7+BIuyKBpoS540bj3R3bn7CCf3TNkNAjXu9oUTc/1H75Z
WEJQ5iHWiZZ8zocwm1m7HV0KNC9OweNHMknbDUW7J1BELRAPU1v641BLMKHijdXW
oh3s1uJyZnk7uv897qICEoOTfeP3arKBbcJ/JVKDFe6O/YT8mzeWSDi/33OTIbnR
C6vuuZPrF4xWliYwGeYXSziC1B+bFx5c991VbyF/9Epc7FLQ5GEpPi7/ZGcymh92
RgKCMZRzdjF6cukcHvUh7J9vGsQ0d/ceiK3qLpn88i+imF5ai1lhYd0UEWP9an4d
KOKzrkTI/Tf1TpfeLKdHHWeS7M+VkvXcWBR17oMjnM/LPQIK9+V4sH+4AiwKq4lc
TWIihC+5+kQsuWa6M05B2eRpNAARvPw74AawFSoTJHAxdTfKantLEXgWJoSdD19q
8fyroUfHC3CJZ4nXZDGYLQgQNXITt6t3Zb/tX7/kUbKK1n29VnCVwyZIbSwYCiSe
v+OxPC3o+lNmcwOYkjFyUlJBo9BHl7Y/aPCjrhULXPxYae8iI+PnzaQPPuNaC4Mq
KyTZGJKBkcAv4i5NbEI8nwcmIee+9VCOwMXyYS9e8xVezreVWwmxsh4HsAEZYEl7
qKu15Hp7j1xz3oJZVybQC7P1lk8GjxdxcnRiWKkH+6+xw2RUv83aJWjt7S5oB832
2YZkv+k+Re16VeHfyU7Z7vgv9hlbNs+qYqxYJOY04v4vP5Ya1EYYrdeCFH1/Ao+G
TgQ3IN3KdTKnBKGBTDh9Jw9h3uSXwY1egbM0/6OG++y5tp2ws9qBuD5Dkukip9zG
wjkkQdhpHKCAZ3ZdPj32lQd1L9drcqGjleCdy70cPWibGDnaM8u2mK+HTIVbUzYa
yGKWNxPJXeGQOtIRkAx068zbh8vytJ9K971AQylyXJskRw+FSMq6V33Y4i+2BA5E
x07BPkhpWsI6Z5kLMogIp5JlkIslh/5UmxExE3894sMAeTGKgsqL00kvKhiFOCAg
x5gEwCxGVWwTJkLKH5vKxhs1SCvM2FGFDreRbKrsMOv2bnAC0E94hLbb2TnxHQhx
rPKzsjxO7QsPl1+X+35lEkBWaRuA2sxo8T9flTeW3Ouu6/oPoQH5rfOenJqQRpu4
6w9zXTctEgiTDQWzNup3eIq3b4Cr9F+Ddx9H3gtmo7rHeFWJW/6KilNvkt9HQonU
viEONuSUfzGXpp5gmB4eyZuOQKsnQ6kz1zioEapFRZx5LKDM6aVmZoRRWLxKcIJB
yOwHpw476e2cdRxPmOhl3GHIJEGKdzjpsW9iwLAsZUZPWY9iqq1H3k4Vvvc0dqL8
Ct4RvLvK98WKSelpp+JcH3NpaMErzqjdcV7C0wbK8E6hDvsQuZ9Ve1oaFuprf7IX
BUc1EPEp9Ygc/44x83NxrQCQl5UXtQPpifJ7i/yOuyFuLK2RoOfwSCiUVy0e4nbN
RZ/YE5aa3EmqHva+ikN2KxtWZ7mjGkCMt05JTSPbZQ5f7mxNXIFo4YwcHCxVA+IQ
ruDYsJcm7lCoFAx/Uv9rog0qfeRW0Uy9TboPWqBbfJF9j7UyP8XrdDHnGWwZKtLZ
5ZMKDMkAK+yrZ7ENr9gX5EutX2I0YkSJ0/Ay4teJJNYAb3O/oKBLzeQm7JbFexEy
3dsuyeFu4osDwTT/9/ThR0cSLlvfP5F+PP9Wf2tZgRb6P5W52K3DwsZcQGaGD5Mo
suaVoR4U30ukhRztfKinWEMqk4z6bM8T49Q1Ygw2ogZc3IlHdRCPRmjJoGM1HIq5
rx80jTLaowRNpP/Nd6ICJa7zBhicjqNKu+4QuywWSTN+PN9eGeqDQ/ssXr2rgTOH
w0VIzf9B9GJ8qeLQwFRGLPpGkNruwJusDQWrynCc4CgT3ESf3dVPZFH+GufHAgCl
m7rgmNyqzGk09WMd2Mov2ZiT3vJeIn1PXuTZd4Mo28riS9oBB+7welbR1UD2M9Lz
d4EYhT9loeZZulsmyCOhH29F2ZbIOT3pcyruAUaJ0/tXRygmD2AjlAdPT3YwWO5e
hoE6DqV7pL/dYvPkdCreL6ianU7KEfNLlC1DGaRwN0oxBIbfkiLexSEs16fJOrUV
CeuCxq4Z7C6Ab0BPNdQLDUHxBM2JdBq7BmvhXtv92TISiO1w4kLWkwTZTX0zkOot
ZfhAmPiHuLyJRkXDYrVREw+wTddFYcaXCgI3NRT8GYVoSZaJi/F7miAtsJpUfGLS
w7+JoNlHUo/ozB+7m7m1gXUYiOaRBDHKK9qSHpSol3DfUNtmqAlvFMiiO+jSKg++
tWCm5DbW4lfI/yD1VDA1FYBsfu6CUGLmTW2VMaf/06R6Uhe4CSUdw8dB0NzjGuho
H14KdjVNFUtsxBhk2jXrIQegz9IqZDpHoWfCsIGef9tGXSXdKR2b35EeAhNjYxI5
koI1qrGhBdv5o5jAxj/byG7IZNX6v1JnBuiOsT9fosRJ9rrOA9tqjJlXzUaDOoO7
16g9ezFJwjoGSEH0G8O1XeG9S6Zm9jlKcm1zBLAs/FrGKpFzsTsNpseMShK1Ti+i
WoDC7fN/iNqSU+4rYI6ydl3EZXYOi2DwOjxQpE3d8AlhMKLflifU5uPJdxY7De/8
BsNCeTj2SCSsIgalC7aXf0wd/pQrkuoRjBLwBP1d2rXBFWp5jzG+sTb5xFDn4yNH
w8+Mj4FraXRiEo91mzOuaqQroTuSLIy0JY2179FgiC8fjgcUZs3van0wXH69em8q
BUrqw+aaijMeWHaTuctxhVTKkJZZSR/gbF+SG5F2X8UzSL6ZRlo8pPM4LRB7eiIs
j0cYh2EpW9Nt7Skgl1zQ+tJT1hbBHz9mYHfNXnBBTm4mxsoB5rGKIKPedpOjNnap
t7DWCmiue8pg4ZQCIj38lS6N7HkRn8qxi2P4wOS0jwwYlpQDMUJIqPL9bOyPbwLJ
S5FDlX44nZZHPy4gH2nRWn8abIbdYurtNQp9rXK4ruN2j+OBaXQ2/Ltk3yuVOFOa
bw+r6E8ZKsZ6LmiomO7K6EaPozRUz5lMnndb/JUQ/QHjw6EpeBvuwDUK3IQC3UMK
Csfpj2GvY4cfSb0eTeRhvzppBaaYC4SzE06ir69XB9LcYKrmfRuAptYkrXzFVPOt
9KFt2sfBYMYiZYvGd7lxqzjIiAK9eCDTqP7bK9rdtocnKMD9H+87E5+conYLAGjG
fY+lpIF/uSaFkWgL/zz1o2zxbuDuUc2FJKP/tKWZJDSIYfoQrtFgncnX3b7AFF+K
JNZQ70zWuyHoI9iUfgh1qYncoSgOf6N0gWO0mdWTm3zOR6J94KfMs/rEdTTKBjAB
ZGMwxsV6yiAg+Jsd3Di0uRH1gAcAgPVE5flj+hhWR2l+EVUCmrQ1eY/kfRtUynK5
LummPBhMqRTqdS/hUt5Hvi2CC7AZA1caU4TMrXeH1MmGD7g8sHFSPrMyMUXINL1U
3lGOVkNvt0e8LZaQacw5YGzZqVtpzNTxRyUIOhtBhO92B4NrPV2wAIhsCNKHEYud
lZRdG2sWw9WK0I2in/jeiBns7HoA1lwr8c8NzCABTi2xwep8KM2DGyw6FzTPci1P
LcYWkC/uCAgOXiFQ55cerDNkhsgoRpQ/7MqsSsVdj4w7WCa2Jbc98KX0iiJJgR4g
+Yq+rnJkal8jvRnoBemxA5jazIop64SSGSxOj+OGZCPdWOZAJ09LYZh+ScyhoHz4
YI9W6VAuQoyR66R/4SctNerN3JL+2npJG45rVyU7lPjUGZ+VYeQeiIOI+87DfxHz
5F7sWl5RrxY99qrvPyeyhND+cCLK+tqQwwryBntKHIiTq2Vn+Vw2zz6iR3oQkroe
w4suHXExkb0/I3ANx5sykij2QK+gDqmnAsEwQcxJT8jHgVhhvU4+3w3zEDVZmADe
yj5v0K3UQLz5S9hhXSb79+9c0QiBMBqRfPX0Dh/FNEbzLRyVLy9PTfuq+1VYdQys
tjyK8s9jjKaMVEA/Qr6oHwcRC4CCiUbrpsT0JFgpLJE4lTJAejvWfqLC3jOg+REN
RGSXzfJ4+EQGeH1qDWzzmnApqVsYPhAN1B+6R/D1Y3sO6vlBwoS3JWRfB2eYLqWr
yb8ukJMBxh2XS8sMYyGH2Qus1AZYkwKy23stdsDAhlIeLqdHHa/SVd4ZY0E1Qw89
svFnlA7f7Bzb0JyU3N4yS1+TDYXM2jzU8fl41HL0UVKqmxxM8V11R3oVgfmLBYRH
ZY1eDM9bUKIRDxzPmGMZMCVEHLzGf/aCSR6twlGKtpt8GgSWxtiQSTSRIFUmF27K
EPc0lZ6xbQ/OqVLRsfjsvLBs1fvw2reFM/0thUCiN4ZD5s9HOEHTvRdAAw2p54aD
kGxqLkfKHq5xAbk0b11oa41DqAMROs2jGBY/VTYKntdKOYLeRixY/4pzJWdAzK3u
Obsrq164C5UtPiEwuo+Xep+xxY2JkZVGrhdoylOfYjn5osM9yDCTwrP+p5ALrz05
XXBCN+HhMaRxwkQ8mCebmDdHFN+23MR1ZoPn4iC36HQb1gLEzVh6jbPr84MqJtIk
dBr1lHmilo8zy1wbXqcFutNOnRrYiTTCZ0yL9hH3fPefAw1y31Kh5k8Hc1gKeb0b
wlCsezA/8LyQhtMDaExC2hvDduo6HTYvm+5FJ1s/hdRlqUutqndAS7hZdEOgtDGY
szAnBLEbx5mD1HXktgqV/B/jaTo/8PyVeeScrbVGFbdDEd/35XscntmmhJjmRZ98
gjovJuIIgovMtrHTpsKlINoRjGqGzoR1I53ds2IhOkOYWsB0t79Wc8N7tgbNlKNp
X7WON7K0xvM6k8rjKyMH114BXMASThyBj+CULA8oHCykqHA+/W79Bgi0fvhpep0K
Dd6ToUrzOqao9h9mMX2nhbkSesM/TNORYWmvQtJ6TBiOUsXjJdR6WPCzgMS0ypRE
MmTHLph7AZdYLqCSr3qym6k0IC3ZDH/ANUE0bMkUTqZ23ovUW88v3SptoOkHgBaY
a42cPLMd1riL6N7/yCqyL9YkqU8UYfC4SSwKhdJslP2Z2++EkGTaesJpkIrV6zIr
m+Nz6Oa7xVKq2gMGrHtg6tahA3ZUcdLbNBESKeEUBxLA8UOZKjkgfBNzUZgPOisV
x4Mt0cb4TQyyKkqesHRhu1TFDZ5yIUD7m9KzjazFsbYTgQPXWMKOpMW9QCivdeFj
MdB2yKyK+d8cuSHLJdRFMyh7cOLQiv06fGUULrm0F4zAqatl9uRNnIJURVUZPf8C
MXcDdrSjKrVluW97621H+jU/gHNG5MJyKCOyYCrdFF2mMnJbNg8X0gI98naiWJEo
AioRd4hLLEzuDVNr0O57YIub3M3uJO9sEKduB5MPYWDJ7YRS0TJiYpnDKx94ybY9
RNNFYcA16fLgFQ2NntS5h6ZBAzZaSu9JygZEMbDU+GPgoySO03RmP9BY3w5gNjLA
eLYxqxjC0r0EE63LaMkQY8u9SeHSYEjxC5B/XB0q4WJx8ZE3P+Zdg4mJSUdTHkAy
Z2jGkIVdxgcJgOdcwKoaKyKbtdtaqi4/sfMWzfnSe9J807KeO04hdG7iC1XAWh+8
NDFG5L6UK4UKuBP8woiqPMiHHLMdOGczVw9JylGHBpC16VuZ5ci1XHyf3X2PUepO
ygepMnaOtZMKmdndczzyiuDYFN8GL29o0cc1kzvZK2SSW9WD+qhl9gK+3lLT1wXV
28iyt7fIHPrMSWxrwdkvWU1Ndak0R7bVdHOdX7yGhA7qzAP47IihP55f4GQesmhm
a65rwWUcq5DpZrR8k4AZfHuJdS+LtLmUMZFtHBPDfuDSD4P5Y9i8ZiuEJWIhnbhY
tvDC3ZLLLOYOPPsvCGEeKC4SgQRrkp5EKbRBzdf+AKYrKx0MZkKP8WqpRJmdGjgF
ffFYoWoPjxDfX4OZlTQ0jh5c4RwYxg2+47Z1R0aU/Xt0x/r4nCtM2scQx7qUUwtj
2k6UT6vJJemKqKIoqD//jQJYLt+NlC+7lEXkv0XApKyF0mPLbpSpZe776tLshir8
UIFtFemmesHTyDGpLYr1wqRJj2kCEMR1lndmAesRv71vmdcQMPlDaRi5OitN6EtM
7zo9+MRNqkHQlArj0KoflRpexDcomTzm1bIkqDnTZLl7PhLYPFTlJBx3+bdnIQu6
Bu2yf7+Wx2YAbzTSq3QqL/JtNUOI1oW6YiyVZBO2fk6naSrcWt+AQK3wlvsLTwhX
FhBlD3vWudiIXff6BjWOWuxATa5PgRVAoWYByW0o5PMWdaAU4k0DF/AClzzbHMKV
grkwYoEkfoFRguYj4idvi8I9p0sYq5MMT7idaOAuKatEPYpOGUAzcY6gRj3o5R1/
bUaMWk1DGp6le0nVla/iDULbVNo4yaHh0GV4lDuWRrBPv9QT2qu/cYZ38GZLByMl
3gkgmlvwHgndvX7H5JEkKoPRIzUsryWMIj7G6Mp0tMBMAI0Q1kTJ3O/8j2BDnOIA
xAdKAXnC2w0Vb4UsK7gqe4U0/iRdt/KVtao7ubmvE8ouS/QoGCh0o65Dy4NO6QKs
MTq98yI+NeIc7tRaPxXMd921834UWBElY43mhOMEYbZ+oL6fZCf4uk+dY76LMq/l
0fMQU8zGmG5Uq2XIwjB1AbYmDzlJtmsPAE59NjW/J/7z/+rqWsKjbV0vvA3uoQAr
NzoplAKcRJp9voV8poxjtWsMB/kn6RfxosLSiDqLKw6y9KH9K061V2ba1h6oNIPa
6VnLNaRo7Jr8oVa8a/D5i72YlkvHiztqRYh5r0SegcRTyxxuMcGbKHGbOMROr43Y
WZHvtV58svzVxHXg9c0j7x68h+bbQkGIa2368iDZbtATmkUllRVUxyioz33U4PIS
+zZC6TwKCxxecdbhs/rQIQaIT+sOn2UNNF0pdJEFFVZdwvcfUPhR3uz09BZATbs2
XEoN5XKcml2/rhRhIfZjSGBoIfp/6gt6yRQoBnJMAxpXWlL+GIA30NZAjvGtIjFM
C2EY6sQFXVbUbIilUE+RG8Aiw4h9AslPSZJXK/s29cBhgMqQGSScsYlTUHSh6hCJ
uOz6UAwOYhSp2sw7ozogxAYNcSCDfr71197g84UstBlDb/cS305n4Xm3LquDW3r/
fZr0K0X/HxUwnwmkKtoAcJ+yFaRnIY4J+6tfsLo2Rhg2JUV9/2wfmoRCuvOJ6UnT
4v4gEE6GDjsXYpXMlLgykF9U8B/tTFMW10RjlZaFELhfGmR0RMZmAskeXrzYWJp+
cQF9Q3FlRHqAeoebNqRnQW8YhYSunaS1DqkX0Qi16zGQq2dxJrEGWOplqx9USwL3
cuW9SM+dGjyYkiMEXskRietZN9ttz+DsJC96UkB4S77ayz64hz16tlNeXhKV5btI
7px/Xu4Sh9I6aOFhl+5hkXYFKXhxNmT0HLE1G4q7XNjTWiA8+riE3KLjYtH8UoEJ
TaJzsYMoUmxca+x3uOw8/dPt9XWrObnJsIacMiNBKPhBDKblGEsrtWmR4B5mUwa1
TwcWnTaLCJtQWgxxJqFo1UAjs8dHzFE+fpRHEON8N9qaAtuj0yKORMQkycMwfGmC
XRA1i6ynG+d3dTCNHpse4l2wCPvPA9jPEGMA9B7GiKqGRs0/fTmE26jNdgeF0TaN
K95jqdHcdcW850xI8BEpmeuxEBkUGihakXqROZs+tUt/VNKLtc/o8c275PvFcYwA
GIyVd1KZhdmdBexmiwHQFW9bE/8AQSQOTDj6n1VMHIzaDjbC+33HSknwA8fNP4Fs
Ub3SKhuuBCBjrA345YQ9+YrcNiM7StOxF3/wP0WjVZmYgC5Av+1937heeZp4QpLp
JpODvcXCHQJlbbncEz/U6WgiMPHfg6fKvfRH6/OGwWx5s0EhQgfy1W+EgK7iCXaw
unLG3/IDB/jVc35LJyYlGMe1ZZcf2Q7aTN7cWZrGr0B6CxuDAgI7IzlE80AhQJjR
4g9dWnS93t4E0CDQYC4FNAbaK4c22mtDJr3X57Ir9PAlX5ABWi9gbT4y3SYcwo2u
2sirYorqZ6EPSHkLEevDFmiJpW1ajhT+NluAwVGdPtE/GYZcRUGdgLFdyjKod8gO
b3cHXtn9hmrcku1nfU7BEv6UP1/ba4P6O6isXp1PrkJCYIZ65sag5XbPNv+rq4Wn
XLuh3+w1omr+OtEgnbF13uCb/pzC1QxLIrtM1um4I9nuwiuvzwgwh5I/3MOBKJWP
3TsTWeBorsyFDlB7mn1hsTVcypdNBfSx7X4EEenYOwhE1K/Vg+BP6NIjN+uD7M4u
wkbiNa3Jpp8iahu8ASOEfrRTuQEMKHTeA28yN4EzmM5+AZnqaGZIpnwyRR38uDlU
q2rY3XgHXyGH10zMSEwhGXGcCCesVt1NZw1iJ0o90G2L7yH0SPVrKZjKfB3lUHto
1eAohC4YeAoXNkFLaq5bRFUPew5mzWk2jel8fLRNSINPVKWFlcYd5E5+BEOrzK7T
whNc0FNZmYOf97fF98pZrkz/5NCGunx8MwtOMu+eQ6WVJrYx6MWO6Mr0y0NIhm1l
QnHQt7wovtQqiqSTAM76Dlk1FD64ZwGCQ30/IkDKrf7GiBXPDbUvM71uHaTAB3pS
X9wTYJ7gSlB/OJVho3Ab5XRysxanGtGn+Mbj9gKzskvWYeZ/+y8hn8eDJmrvVu7x
GvUSJMlaO32SIlhB44lGIUZjC5D9+OT8Je4OAS/fwJSgWbdlQBTKlvQphnHSuwaW
yafTl1tYhESugPasks1Qt9OBuOZttAAfw8uiXIdU2Ei0OWWLrTmZbKm0ZA33WB4J
46s5PnAr6xtpglZmFaYxnGlRJPaX+0GZA5sz7rY1W7ZhknNVFbb7tsa3xNKchxvT
f7GLXVrswvPbkXhBcx4UcOIRNUKvVDSH6K/w/PUtu2l4YYABXHY68ACfZBA4v8j+
a34Hbzhxhe7zeVRwbC/qedR9RYA5BScLn/sywMrxgi/Bx9DzwpEzvX7101pG6ylO
0i31b8LctxwWzEevp1JHcEOs6B/N52UO21NRkNR5tsxZZ9vSl6dcU6EPoK2ormWo
AkglmdVXz19rXFSM19bKelGnufAh0sys4DH6WPSbosUlIt6z6vm2LpKQlje3/QqC
H6DyFWy+CQuaq0Nu5f7rw7+dVSOCNtyHfQuc5ltwegBGX4hzRAT0y4pjf9LdsYCV
G6qQ9ynBHobjpBYtqjPvfpl46sqY6kYEN8kpoUqaXoUYfJ6UbPVSDIVdJh093uRS
HIFhjUaHRJ26HX5wul2b7r0OipvPpQxbINoZqHImXFFyFH5DM4IAFiVH4Ak+jp+i
5DwBK9STvg/70socWkQbAQoOWPnHVoNhYvEhg+vBfLyFJ6rac2V2CoqzV1gZ+1z6
Atzw+pJ97fitzhSKhrwuZkoQt3JU3lWXRr4cKvhq8eI6boNLpOlMitIrK92xOi+/
6S6K5V6p2NDoayJNCBPVdDdwEsrb1GaJgs1oDunqn9+vHmY8mxLPliR7NEvHbjBR
Hhz5Z7k3dw4FXkGrZG6wh8MtZQQZM09KLn73GKnRp6riNg80SikbRU5nqCBv53TT
ShkT64S8LdjaZ9vlgHw6d6c0cY02r6HyNWP2NtT7s8ONER+hqvhlP672ahxign1b
P/woyfVNGbZA6YNyzCk3BkMT+rwgwYU1zLbMi1BwLboXFNVlR7fqEmkqzUkkw9XR
zdsDEdbVNeata/3PkN/UDaJ6D1YnKz6yrclVR6Pru9x7D8AHt5rM9HUdRidTY2hk
+/PhoxGYMmWOVTOsHGX8NbYAP5IzWoZumnZQo4iNvq0eozwCT3ipwmpMEBtssMM8
74KpHpjT2NhAnnmi98IXoo2nsxOGBo6a8oGKrvhJtCVhv+zqcA2BCIOiqPdzn6Z5
6AcFuOVm5+7uJjjJ4CGF7X4axxOD0xONpNTNb6JYfL/xw4+gXEklPzPc4QjNivA4
NNHPs0sH26OaDI7XB/NQjGh7ZancMFXfsiG/cXrYAtKHW9ENeH1nU0nfHsEFYm6M
FA3CN7vNyf9bfr2QT9w/jLUMnBEfnyIQswY2Rq7X1ytYGXdeHmUpWAPkgthNBuKE
F4fJa6qTrqV6mJDYVGA8cUC4C+W+nmRyyHfsoXjsAJRlIGSbXAQbJ4PTG5bC4kxo
q9hO2XN9Ha8hnQsum2Drrom/dxd9g7Gfhd9teCP9QangJ1RQ8+0n/vCn9nIIBtyL
BNFfUZ7QreHYERJTdjG93pQpUnD2rjsHl0/8opWj1JhAGrxUNEMGDUza6ye0C4dV
GZ6m62WmyzSRVtFzMhcRI875qAqDilJ5tjWEM8rLpRTw2NykoQKeyeQ091lFfd27
3OpKkas6C62YSpcaF7HO2tHwHRKbmi7oB/77C/WFLW7ISSFWp+pYDDq3VNfYJnV8
Ek2jvy5vS0jYuw3/T3gDRzL9kaDXGgpmAXvMCUrSsNeXgE63WM93OWeH7gNsbGez
aeagGrfGs/khI+wcLwHfmQxx6OMLEBEF6v7T9VZQiCFqdj0QTsZkvGG2RJQmfauT
l3BBt5yr4m3+8l0O7U7t22Q34qW2RW7O/VpxLwTTAek2a1YPxCHBTZThx71Bm5++
gmMd65hzSGdGOLFMYqdKsB3Aj+n4fG6+rBwy3DPxrqD7OjQjtsnNBgVOw3ybuefl
QJCPgqRKtoGmDfcH3pOtSnF7/6iCW1ZwqqRCZC1e8oiVnx2ZIthnzpH7wsthW300
fVPNoE5Whx/9zE40+mfmA1a4uHXkiUpVXY1J+gWbTtZVfVzBv/Mhz3Dr1crkPv2M
CdCRo2A0L4zcWYYG0NG+KdXycGzxBbyt3Xy0uJTQtQPa2FL4pdaSdPlULV+au1Vu
jK2NsMGd8u5Otec9AlY2Us1I5rUkufoy0M3M8fKH69xMqR/nO9xCqJNM9lUwafsi
BMyPiC/n/c9ePuy9Bd+QkvLMxzkk1f1c4d/ZW0jNB7Rt4nrWlQXrY71bplbAvD4/
E6I3ZbKt/HX5WHTbf1aXg5Fr0FSsNzgkcUn/WLwTpN8umkLJ5DbArbYDAB1A6Don
6E6gT16TfwFEPi5rtTrrvBKWvgP2Wu2UjGKIYxUPuWAfwSheQtcpBXbNih5C1CoH
zkq1tcWw5djOuB+PMoRc6eAqbD6DVNRwXklARgwDIIRDGzsxDi7tHbou0usqrnOB
b7JfM/XNleRxoCIR6AlIJbz57e9EUkgbifEzg6HN93t2BIwicp8kQ41qwyNhBggJ
9WyeNM66j/cO8jt76Oa/FMaltKWfw/4c1tGCZrR5svQxMB/6Q2nI/7R6/XQlXMUQ
+hl3IOzGhkl87oNa2WGvRl54Ad+LVLgJW41+XEeUIKf6DQ0t7kI+n7D8GIxkq8r7
JRqyqaYuLHEChqBMJ+sImbXiTHo+RzjedoCPvbnJTgYVGp3prP2AAinPIM9IiWvS
Bm7oosm8dB3Z0xUpr9IDJZwP0ETPlHKHVunlnEAN2LDRyDXX862KXtvF7qBoC+Xh
/7BpSJZaBSzcoXdBblr8SyUDJnDJv9pXtFq6CjwVI7vBY5mYHR989mi6Y7pq/IC4
uuy/73IsZokIi1LnfD+qLtgnSV3uSvh5L44s2FEZuYGVNNUnxATRlv+lSRv04PYS
pa1GVpYU4A+fsQH996TYsQfhA2FllrbyY7nQ+ieJ2VamvYjSggzgZnIVKb9EVziq
IaNmbP7LyFFSA61cjATHE8zet34PnxCBLZ4g4cvpQlU5E2bhHyA4fhnSgd9itoby
xb5EHL1g5KCokRHJf9d7iqlDIS3o06pGIj7rMP7od6yb5Ci6bGokjI0ewADjpZGw
sfDvCYx8MEVOcLOjtSTGi1/MDVbDIrAWrsTUHgCsjJFgaiFa8pHVb4g7PifWof/Z
9BzQH8hwDCiIz736HaDTwxGFMH6OmMwQXNmnRvgg/yzGwnas0qBc50wNGPMsL2Vj
ckR8tGp/Qi9qWqvPdtQ4qX0b9BCDt9M+K5rM8Yjf1738ELNP6JZw9a26ELX42vjj
QO6TJtQ+sJm3u6c53oZ5PjxZtdyruKtGgdsAOhmJSt7ThWedNY/0U6U3xbU+7QCd
8QcKXVM1XdfudG/+NV2gMvDrIxCnxSJzFjOxZoP/kJlrryOdcbRoPTGgGUJf7/yR
6iikWifO5Fqx8lYh6yVdoK9nsLBn6SbRb91oC4NymaGk0xtdJpFVIbWsafjmj8fd
0oDR4VXWTbNhXMp6/mSOfqO3oDVlpr4f0N/xAI4UqNPha9zt5H/XNFUPPl6DU8FL
8Y+a4yZHVj34hV3HcS1S4CDy7CKtbbcYg6nukf6WaNV42WENr3AvmwyjrdNBPVNE
0pyhEgxQ2bwal9SkQ7v1lPM+n2/6xLVOHbvShGWn+/CVnuAB2i2eI34fw5Tkfa0E
fA4Z43/aEAqmv9HcnARw4mPtMyqdmf/l4euqo4KT9I95h5JE1L31TJCkKuQVlAiD
2PTgENAEsc55yGzZm4nIDw27s/gw6xQAesunpruDR1jz1o8ZWN8zJTMzFfFtSX3A
swHPKeBMwRMn/zBfVrYsCuD+Qf/0eHlxo8AaOi8EVuaRNXsrdrRbvTGOR2NnzArm
XfpUInAF6hE6qtKEw4wzfympyeG4v84f7Mnlxt5+DOGujAjd21gD6pA5bW0pGSaJ
AjdpYxm9rcSTR9AohD4SxlgE9PRJlXDqT/r+QIilFim5qn9YNKAhi6jznp158B8+
AOTlei0pCH+xyXn99A+3m90pI7/oDe6H0gf+Beozv5wELOv0g6asfQBoX8HjB4VA
6lOQUwVDi4I1waPP4Bm+NpcOMAcWhTA6xL5g1NllO9bCQ00W1ql2zIjmxecbt/f2
UmzC1R1laY0nLJiDen0E0bmRUjyn08Q8GXNMjahMKO/wpnr1OQyxRVsxKGlW8IDD
Lz/oiA2HvjFNsGHdGWYV0pjiZN68z7OFwChaiyhWKe+hUvtTTKPeJmH+f+kEIAIh
eJQhf3nDqNOIxNcO4l8cuku4/P4yZ98EltcI1cVVhU0djsoisqO+iEWD6t7S3YRc
YzXxRfYZ6UgSUdggLg/oS+0Y69LnTNEX15+s9UZgFBstmoPWDdRWQNVdmmFHUX49
+h/VUTxKFPUg/YAVA2RankR1DiWyYRIZQYcSCGhoDqN67t/zwh8JTWbstnWpuJO+
jvTEHJMhaEh8/AODjGMDXvPAsP9NylljYdkFMBeGW53XxUrqtID/QjqgJ0TSBqWw
wvynZTsYXYKl5UtEF5r05VfjenRiT6y1XPoG0eshMA44xV5TMIY4QDpu6ee3fMvs
ysWgUGiCv1XgrjHKxhhGOqqr5UDMzFgoOzT8Gvi7dcsKHNlA5xMc7iLg3Kz0GgPc
ngooqzDKk4llhBsovSWuki2UFjo+HmXXFBaHtyStTDHuoqTsBKqgZHi2WA4NYufG
YcnbLsriP5cD0j6ep4VarKZb647hmVOCGil0zSH6u1P3QV6n++p3oJ/q29ZzJnU0
l7/zv8wdP4SU0fmptZELedpP//VxErk+MiuiEh0obnlLDrKsYOCHuWBQ9ejdy4P8
9E/qrqt8Z2yBEl7CHdnt9lzRvXxCjgKNzskuvtBbe+rOPuaiLtLy9BzJsuGqn8xT
j7LL2SnMlgoJBHwbz5GQwgofEoWkx86xDkggMt0/JcOzz3iaXnwmdaj9y5QptTd8
IyMGah/qJjynNob4bnmmokerxyw8512l/Kq/KuVEqsV1U2rkgjoWqbBHCEn4Wb3K
09EkyFQWb6dbBh11djGskQ8i1VCGdbBP30/TrgGas0JwYWgaadWQIBOrJrhoRl4y
rfoCyo3WupXXetZzF/a43cWuLm8F5npnJgiHnMnvVWabz2rMsOE0va5BWGWvX4vZ
Eziu+fKogKaVmLJMKPtSU9FtCvsv3ZVkUZwUIhqAxhZrS5sjvBBly4Qikko3mVAa
5yQGoUN1PjAtsLz59GKdZSdahQ4/46V/0+K2H4X9CO1k0oNvmLTEOJIdLmrCAFe7
0Y2ELB1HfRKOoLcOMUSDBY9ulctJ40foRAL845HdhVzUnBGji4m4WySihNwbhU6i
BoAIVLl/CnUhDNGA+XEb3yFtPu23lqveyiPc9C/Cp/GHF88dMDqT+52vpAeWPN9v
D3egtsT2NGPQcbmVSrWJPREqhP04+u/TGbjUp2PEbEDQNDxEDA7XIUHx1cd7je/9
j+Umaie9h32q9RBQuy2iNwKSGDv8ebdeJyVKk5ytf/LfB8JlG+Mgh/0+cBk7eNsR
7UL9AtY5xPqgaVi5GtjH8Ylv8Nd6qFMF3X2x7KvXPLbZI121SICFgucSbmdGi8xm
fEUZpV6T9riF+4ex11ry0dR+R9tladh2LUxi01Qrp2SpaoFy6pNDN+8vXau1TfW5
l286sB1R6SBSp9KF73FcayVv2ABBiYsWTnX6AysMaFCUEbGbflNMwWyP8SQIoQ9W
D3iNwxrFXW4pOoct1rJHAdm/RzRbRZsCVBO2HHPiX0bOROtmUnJ8gfz6hlcZZBZy
MGBrlyuyNFGnXy6WiATpItUZDU6q/hXshL+/mkMVQe0q3TuyCPULsAu4RKe/GZ8j
r6lxqeyLLg4w5XGwHT+kQCcCnSKrSjKvL3TVsRKLnuxlFbNLms/hzwkUP+mkY610
dlXhVK5pmEHD1iQnf0elTBPtcstT0s2dQ7SWkf7ZP/KNSXz/qcCh+tEGVjW5Bkfg
e2v+3U3eYxwmnvoIRL9MsLRxCnvlFssBTLlYxOjFesGXRJe9Q2NpX/5TP7mfPMZ1
+DGjIC4TWkrPY1X4InUiH/oA/zomjSfMhwo6zMBx8TGyZtbRSTH/UlV7tRaoCf/o
wONqqWy4vZJl717/q7Hx02BrT0z/gO9Wc253Yja90Rm8/WUi8GnE2FIIyJEfqWwo
9h19y1XPm9q7BKnwc1uNu2HgN1buVVajdFl4UmnROIeBcZ54n/2KeuB4mbk4WLzU
B/m3axuNWSABNQeiqLlbEd8XE40oOoHGdlu2BGH4+/la6YWVaeoQerPkath1hs/s
6wK154zSRpItaDJKt5VJTjKu/2NXl6xGiCWcdhEUVM9hZvfdQSIRUdT+X2zR6IHe
jee5aWb+PRZ72thx5K4xLXaW4scSCnIKXsJIlCsd5T7kZoetb//RXvq+jgrKqc34
U7RmVahPfMUsIOPqPiG7dyl8ml1CGgWlXKP307ZZSMOgFlXj6ihn5tKzU09dHMm0
fyxHhIUsEPqo9dXlIV8CvRx/KuYM7VoAxj/QRw2D37nnxLcleGQg6JjdbfUY0NTQ
QA22BwEDz9fxPDxzwp/fqMRMZeiFjKPrOBm01z3E3JS3gdg2nbQzWNUm99k/xbLQ
0CoUrgIcGVVLhOinyt7t+YUWHW/E1Og840FbGG32eRUm5yori1PM9cTCibewE+Re
KDIHRDS3vZ6diXKHr/pDlSnEjbMFVP//B499ogPXy8r6NADzHaw9+nGuIfrKahT6
pX00NpXrfkW4tZ2bSB0If3WUt51gnBh1plcHzDpo3lbn3KAubihhKx5yv4Lb11+V
36+f7vCPaohVD1s+jSZA7mirC6lmDSsg2SpyI5JXnZK9kzH3CHESjxzIexr7IMHG
EQeV+nhvrXpjRpZINMeee6U0cywUlGZkzRxVpuXRpnumx2Afi0PCKP25H/L85Kxv
/YMp2GUjanX9C1C2lcMVhK7Rb8Icpa4wWK9KQSCWBiA6Ekyv8D7fdAzntAH0SILL
K6h7VauLaVHP5Jqn9wcMzVNETv15T3hc1Vab2RPzqmTFQzymBGNAb5C/4bf8zTyA
CQoiLZs785okzJVBR7VGNamTX5fdhK45EbhB4HjWwzpqbI19G8Fb3y7H3OjE6441
LjLJHE6uYDpsV4/vAqsTGngNbyGDwTzpVpW3dSpTkKRQr5yNcNmOv/IuVGpuUrNP
CB1eWYBbHq0NsZ1W8q4kCrWGFO0sDc4r1dRVOQD3YNH9oVjL264Y5uQuQ2D0Xnzi
3eurjgHEpFdmYN624UdQhWz8PCVpRFvIhd1gL8Ha+GrjIugsSjxricrxGFXWNQ1u
/UwD/XbeyuWMD4n7hXrEqS7Eh9QZZal5sCFk21YcAoZArxTtTWSNGxLZx7jmuo2Y
IcI1gPboGDSEXLoUYWO2mR4hDscfXjBJ+1eP4aglEQbxNq/GC/y/taZtCC3SXSYo
rJ2aOg1eHQ6p4UTRoOBHd86juAdHzYo0+wV5DaOmOcmu2XjDHgBQ4BHHKEGQNv4I
Z0tfP6eGSPVpenYYKu+Dx234MEl/JA2aayAHVKwu+edEzaamigPP8+DPPpkfsNY+
RjRywHjhV+DLLKu15FA9Udzh3Sut1zpWTJHKWv/HPM3z+KNNaIP/IJsdQikI43jW
48c23DSCBAiaHBZc5xpVicqrpbUHHPwVj2cLpNh9+qY1NSbnWWrLxTAE6F07JukF
OD2WEZqJza0gkE1JlSQKUlX6N/8RrEcWK0G0wFZUk+ihz1hy4NdUtoZmyi8XJOtx
9qxMTu1p8jCjXCZ3Og8yXU4OmRLgazsV3686rL7uF3XOpVi8lM/wu9+zWIJt6dgB
9RfZt80EGQfE7VZ3xBk8QwtPIoqa3A+k4pqKoPBIqPToywmATef4HsKHQiSztDA4
LTMTePvM9PC74hJjGfI3ticpPFkLWi7yH8fqWYfL0Spnoc/HTItqah6wi6jus30j
W+SPvRUihi7pDo28psgI5m2pIjZQcKt30JGsQ9QuIpbIg9SVzskaEW9gwRSnEmQn
Q7qWeabTk8zNqjBx4d31nYUp2Gz/3BGovPLtpnKY8ImUIGy8FULeNj7Q/i5Bx+cg
2NBA+06aONYgHCLFMGR5OQs3cXX9j+1gmANhvojFu1Ch5xG9WQSdX5PTfgCZP20U
WRnwyxsKcX62qpMSF51ZYOevxbhENDo8YyPoR4eQxzlsz0si+9SzuVKNVAe5JbYB
UzPyfk/rFdnO9A320CocITU0RSs0o2VMD5AXrW0mR5VGWHxveBrfZkn+gFPIHjji
z5TfCYH4rqtQN/W1S+8PlMa1eemV1qwR565ueO4f8gqCcD9hynMUDAdmedKlaUQZ
SloO9LQkZNkphU411PDxhtRa0Y0mVV9AnE2KJBKPpdz13ISCA+rAQ4CayXa/OpTb
2sBg0YZqzHoay9kUlz8bLzxR5jWJWoopNy0reJtAoAprhu+MZrhmYr5XDrajHx7e
VJ6jYXdtQknD5Sw4FrwJwLCQGQsTRqTbXZn1X7KJdrSPNGKUe6jR8p0p+88P2dfB
z3pgc015ZsBWVv61Z4z6izU215q92LVX1n6mDdqMhKjveyePQ0EvVzMMh6IZBbnx
29AuEZodOfwqUJzoN2KenpxTN4uRPGpUTiOP+EErllfVBvcZirBl8XnD6WpgUgwJ
8iRjiRatKkAtHW0LYY87UB1ZLAbeRo1SlJXNxTqXZ3neFzoijAdrW8UA1ri6QNkP
X1mHYbDeoqC1MycvoPeSFiAZLvS57SIE0DSdvEsn9tR7f3BL8r0UfapYHhX2FOCY
HihdsEsa6/DH25DTbXqnCMN8slr3NhCxQ77GtwVvTW2XpOhZju+kdSKB70y4Yf3l
0NROxw+QUbXz44L6nwhPjB7pTMEOPnsx1wHEw6FZKNOcwsNgfCop767PW9uxkIYV
CvWrXhU3IEL2xibU38hmW//ErJPSNpfnujOxMUCJYLDJnryU/P21EF8zCAW2vJ+e
Jm9ysSxp+LvOnB0UgctpvbwGHu3mvFePgA1UqbxVi5hjZYbxzGWFirnyGDHeNWbH
TR2bZSxS7d0YYYvuC4J+WAwUtYv86WqDJj6Mp9pzkBuSdXAtQpS5BXcqeSa5sXFF
K8eleiX5dyv1R8rg+ctMw2h2uwso1L3VKFd+lngIWKnkgdxFkTI3R7a6MRD7PLiC
saBoXDiS9PAM5DCfFK25j2MLvppXsUXpCdpm7qES8OWhxqoKCHlyhPmdGA1rfA64
8Etgq2am6/inUJaY9zrU0sWAVJlhMHzCnUxoD+KrIYP1VL2TL2PjgC7hLPSgZFZh
szoCQOUWHC3P5QKamGeebuoeYfFHb9yg9Qav2OnGVdxcvZqJefOj4gTv227O6qad
WvVri9SY/TbMlovM8FczVhvmOjLLPg5lNjoP0gLMRAtfjG+3gBE/ihHRQIyTM/8C
5aUBwBM/8ylSHz/TWRjcNavhS7UZdO5ftoJ9Quqe+29QcQ8ePrCY7qNJofyuZSOK
CHQxMrRCoCCDXD7FdnvLk5MAwMOLqAZqVw0K7Cz0SWvpL/Yip6X7zQlseEzlLj5o
dE1hMlITPWmbpp2DtSI+cltGSRdEp3oXp76JnzF1Z1MB8tcUvotLV24+TMdqQQ0t
nrK2vnl7G94oVDLmN20Onp7IK4AwTGursrtxIiHHgx230Su6NEHRInlrpuMGzeTU
NwgIqKIQH7Yf58Gd6ul7nfWxVvvbpFmN9CkEB5KRXWIibZBBkv31/S3zfPefDo7O
DJq2AZnWrnzDULt9jayFDJTC2k7b398508BBKCvfhr54/UGBAy5DygoPRUstOvDi
Nj8jXCaE56lZkDoSaCGX0hUtRbBj0kJNdee0mw1ybUltw/qrzZlBNml+rpC3YZE/
4zTuoilm9qN5gLK71y/e4S/fSfrCFY/9SISzJyXCRikahM64rGiWdqL9Ud2jF8tv
rrXKZ3NC7HNFmAqv2A9lHVJgGKjn2EVOAsZQ2je0nd9dNCtGDn0/VgTP8n009uQC
BWuaiDJCeiU7U07f2f0sxDZGEA3AVe0jHsaaY06G6Y2401psWE7i1tERTHk/4ppW
F0byvYp+iCldcJvZyq9J/lgqwL0vP8zKFG6J8/43oHyk/g1DqyXbkECf9hDMqLIx
TeTzJSYixOurfrhQkUxh0YeievcP3YVNdyhi21Xn0KmDIp9szasy8mXMctBumK8P
ovjLB+odnQb05NUWgf+XyDEk2lKnDlhpU0vh8wlCA6q6ySX2yjRbz3BEmqEP3Q/b
975c293ePNerEEMgnmHfM4tK9uuYN35/F1ApUEP3sf03wuJcBavanLf4e84+9Zd1
lF4lCOEB1M0STqQRBeUhylNN70wtfks3vgPrvqP3BcUtQWVKfhlZqHmHF/GJgTAA
Vl9OvH5v8iIuP8ImBxx6Esg+c0lPLrS0l9fZZu6qrc3XRObWeyHlDly03hGtmZ5w
JH9e5QS2ra27ufX1sFFZ0jQ4JC271FnOTxfprDdRmyyOyOfo+pilVaQ9XS4bqvse
P+zSoxjPgjRWIO72pN0We6sPqgUfUsqxT/mf8IyaLwzf2uEBjkbjSd5kqkhJvv1C
UJtVePtKVbWrUhiLzgizdJG2+g5s1M343W5x8Su9BBqXWI8aLEDg1V0wQ/2i2syn
LZlqxIKCh3sgwktHCFZtXu8g7BucgSj4SKJfTTAbn6fogWCJcDPAfsV4PmpcCDED
6ZaquI3xZDL7ypLXSJmvEwfkf3NWrwytwFUVwhA52HQ6F5/gbo71Q2nEKBOybb4m
xHt6zJFOXfP/bCMtOUlHjimJss0oRNdQuiDW64F/C3/RP0L/GvjxvHKdmtV0Cz3A
oRw6B3VfaDBiBV3Qc9sR0O9qP+shMobrS7ArTTGW90u5+XD/t6Mn1o+pJLivJyjf
/Ck9L6njZPGrf/Dx38Vqbqjy470hLjGRcKRp5FiQfT2IHi259og92e1nkc1aEJJX
FlGjzUqH3l04MeeOr2EABJYPjHDFhm21xc/3W5h5CrkNhC/FrFMG+hVxaPHOTiSk
FO7vNLSzj22eRYFDXYgXaOuX8VfTguoMkNy/MgBs8Xd8MxA8ToA7L5J8wrPp2vIF
WengcG7vqtgPC4hn+YmKsvVJGCL8t6CAIgs6SWZmC0W8KltBhyCKxRVpjRNgFhwW
GjF7hwGIOs1KKwXgortKkxzxmlgIQEs0iigJ6i6VCvasRDCVoJHd5ptUYNDooCsz
MoIvomRxU7AmxUVsAhl9buX8OTIu7tLgwpgd31Rysh7pHZjCkyA4ynDdKVHY/YlC
Vy+KCFtTm58J7PYbzUlv4pTK/E87wRaxfiGyKqrrYb/GguLJej16qAfkfuSdqJkV
J50a35K486kLMcxS4TngvtmdWG5T4J9AefRAM6Speqh1VttqfqPkZtqfOBcMJMNi
kn897v5He8OoXBnMK/PlAEWZZ5+w8EJa8ANvAcq2or1ZgBUcPYFCiv6U3pfgnEot
UDKRfWUNIcxyiTBifgdAz5wIXlFgdSk062oJ2xj5jThrYYKTJjzlCzvDa4ZieBWM
TYL9PH0qGzEfx8Ep9f0QPc02wz0nQH20eN7ZrnhNFbeM2RbsDuCW6RvE04lrv3Iu
nHqYjK1j7zSHsME/DBzYq7IQH4VrTH5Uq0jkLoIgNoD0xI2UAMBu/pHjpZ2CLAmz
vqXBHU4eChMwVBdUGmk0+mTwbG+nd3fU0jfR3FNsczs4fg6zkVznhP04MY4cbMSM
abXZOgwD5Zmy7qs41cdPglCEI5dfSzCo9P2m+M5mDP8clDjijtuxOTX0I+jncdh2
5FlVx4zzId9q/Gar6HHopq0owUnM3mXIRlbEPLTjKaThS8GwQVNdphNHaRfcZiK6
bdDw+tJeC+Jpys/qd1hLEiwFJzYxNo3WI2iR01FMId8sPRtZ917XDf8CZ4BInyfn
36d4Dz2/6ER7urI5JSp4f2PjuX/MeAZ4+fJLtcwk4at1rmuJmNRrEflcf+B4yaMT
nBhadIGKhNztcFKhY3fq/rXxEyg2+piqw700gFdHKIKWQtefCh8EgbK9Atv870Js
SFDWMrQ1pcwKgJvOt8jN1knU6//Z3rZsGN8KSP5J0mmvdUbqyspTcInCyuPrwryY
PCHGdSEuL/ccpUG+qrRBZ0JxYvZxCUS4LqxgbhU26Ap7LIaMrH7QPnA57T0BtqBi
0lbsiy4giHAkBm8coIOCzWgmZBNNdiCQe9RT/Oelg6p0+MoygeHWNQ6IiixJqvke
uVbNVwQVQlMVlxW23bfMslWf2xfKAGVVTLyzaZzhHxVIAcd5fCKMR24oCpDOT5eq
WF7v+d1d0RxObfVS1kGX+CiuGgJCMQP2P9guVXVRWSJbhWK8pdZbGtR8tOYKVT5p
zmypkvM17/hzcNvmrQJjJmkq/Eme7DZNEhJK5rMlQ+l8uLuT6lNd0L6HPK03A8T9
5dh5xKL2ACrdobwBE0vQLhgisp6cDK2vZSAwo5ce6OV+mItm409EIcNdA4h2KXSM
wKM4zSanqcDOvrX71AEr2fZr1OiuijeBafnWSHbA0QUcYFdrOd8VxzepjlvYPI/2
VwffXDZoHD/ynKGi7hSABL99pTr9iDf0m8TzkZS+7gb9evNtnipJ5hjSrmLNryk6
VVQ8v1BD+XxqgemV84ng0RbhysRlQ30El1cLXYOY/XcC06hpK3EUFflCuMGqp/ZK
/8EpNaI+ZjqYUL0MB+1/iyAQuTBrYT2hRzrfBE9W2vgxX2hvnw1lkAb6SslTdi+6
ac7076+7aAPUfNIpZVwgGZHk37teRKJ3pjCS9YwqPUvq/vOMxP0/AWR6SKjldWzG
arm6F3U3U7rCa6XI38CBwcUVSYNNKsDoT3AKp8aEislAm/dCzqcQ8/td4A3xSxno
puCYb53WjfAPGJ5jEGALsWTcaAagdEq7pCiyIk7BnQmTIoePougpQj1GEBB031Ui
lymnlNRPzcIy3hHZtF1WtKIj7NgCHExM7uw7vFoHVYvUUReb0TqiUbF2AWvHL4ck
bmCMKK4ID3vSZe+7HrTMOtiUnt0uNdDvuJoYXjoZw3YT50FAVJKEEeoeLaF2gXK/
XFr8t6wjB2eoa5BltDBUuIgL5Kc9LnSN05WFcqPVgr3e3+c2X/JzmHEFQdTAfnjE
OtqJ8SBZW49GS+kaM97D/RoFplk1xXecd/FPkStESmQwJv3CpwydyeddjDL0szbC
tLiAmLZzHcFt5juxm9ttA81NyS0qh02Ypg4Gl8e17kGe6o6a0MuU+YbpbPiSuHl1
AHJS6k5LfZlMZCRrQIYq+cWmzQypZsIqQfQ8HmS38HCAZLXoGBfh6SLecQBGVpIy
NGl9mhtQLydBWf6kirwvWxE2H1o0mvDO2fYfdLGfufbVBd6dMrhFQeACkNZBH4td
Q+/UrVr253cgzlZE4oHX6VhpFhuD7D96mCPL+uwgFXdWW0siSQG04UC8G1HSNiXQ
YtKo+vWK6kT1v5g3ydkbSw8qLc9beOHbzGk2m/YTBb5BLJkCUYqZhC05ui9CsocU
7b0GwiJ2cH0ofeAxfEGkmW5VmEtXfEHPt4NM54Yh/qi+6KhnRJEmfTwIFYHqEhEJ
8czwOQ2iVlZ1jy74xrmbExHo5UGqu7QRJ+o3L9nRgwiLAR2IufFK7gAxPd1cSwWm
2bRpkylCPN0UjdDCOvScknOnnZ70L654Zp0GSn3u/qH4Mx7yNEdQ4zw02xCVJQHG
iJ9Sm7PFfZvHOXCCxkfoNNwySdQYVEuclzPqg7rg4aQdhrr5jkAiLqbAgZOpAagp
PBZlvufYHYpyxUvtnCiNJPm3LBeUYVZVwFvDGeBRYAxR+OZ2fd79VgsLy9fFMT1w
UJ33bHVXxdQ9Ev4TFg3VEjaVqX+WsjeBxCWXsCxzSClwLxtjSpspFA/O3ts1ve7n
yOwDG95sVoGq9IZaWONDdfKXUwInz0fDTeI8aF8V7nA4lN/o/ImxjJMyCs3/I0ot
BVtsqLiMROcvNUcrQJnMGpU03gypS5VW5LfoQue7kLhqfYHOBMm5i0menlQayX5S
d03DxEMrQ239a9LEf5zMOcdaxyJTFBBQucDTzX2E4q6NIxYv+tcMrEkV/mz9+o2U
wRXQCaf764kfltoPkblIlRQl9vcoA+gau8uKKbtw5SePfSPshuJV+Ka2LKK8AZPt
yr59C2fgUrW7WZwgk1vpBRH14LrTu4GdCkRV6lbF94EWpjpMhC8lBny8mh9dO3Hx
ssNB81AfyHwuQFI9Cc+DC91PYSH7mIVNw51h/WaDYhaAiOrMfk65Ts7lDjpWpSbt
9gpl8vl7vG4JtLoVDoy7ZxIKcvv9kF1wwwyL+MmovAINmg6Jjy3c0jPFtY6l0fui
XGqQ0m8ccxGheNo2WOVrJUS72YGO82iMFNpnE7ge4pHxNLuD9YIYMJzs4j1shCgh
H6aucbmSvSAIhg8dyEhQ0PimTur8a4Kjf8o6AXZYrPK1QQdTzHOgCA4s9ZXB0LWG
c5rw0uXZMEtTiBzMX2sfKpvToSoaisCU9j3RM7HPl4JHzdW8HFDaZCB6txwzTeOL
yGitmAH7FmMhu5saJBQGBSVkWk2/ysluI4/O1HrKRUKTD/zjFstB9/8PKXdQzEmj
3+PGZZbxwVp5AYn11NUCFxndkaUDXuyAwG1qgwdAcCciYVLnRDecXW6DaoTDkf/R
u7M6D0NdevJl8JAFDS4Mnm4y0Fsj1bWypCebae++FTpMvm/vqNc0mfrPzOL8TSF5
gFBzfQwg2ozFJQZhJx+1oExud+oc8HB5YmNmCOxDBQun6sQZuKqVCA69DKU7pHMJ
XwFULiZ2GVLxQEI0J5XDX02UlLFnsAsf3IqUQEWhGD8JO3fEHIJ+GOKvC5FEeG4g
ovuNSHA4zve/hQlK6+9HfsQSiNFNeKt5Fh3E6wnb8IsHFOnbF9Cv6wUnghBp6QrT
NHpNhW5u82nVGfDpPngMEtvG+zm3o07lc/7MZwaf1oqUSmYp7T/yCT2X6KljbQiF
Nyysl3zkXldvNCTk3TAfkVv5u22/uPY3WDkaohSVwZAJzBPZ4ZxtM71rBlpMcoXQ
4qMr/520rbGyfehUI53ZLtqZqQy/L/aBmjqhsBbzj+KW8jYc0i+ub81VxmTjDULV
cB7M6RVqxmpLykK+buF+0pxvfW7QfobEoikMRIyjdAROIqIIzQTY/MkvneIbyizE
PpQueXLWza89BUs64nKnhwI43a9lkqRBXVWv3jMqdw+mrDyRrVQWm+980wnjT8G+
JlRpeh13d4aaBsDv+6utm+Z7EAjqn7hBP8wiEcdqgrxBA119z1l0oeWN76EC59oz
7R4GBHZQ3HaFYpZ/KaQH76+So0pw+8MNJsHngpg3GGUBWRQ6Jbxt2th5bZGuII0P
ss7lU05nYMMUc/339aEfHvL/goXWqkqKo4F9T7X8Fm5itwuidz4itSBW4/lp5cKa
xA+nnVkWZD+F8TaF9GsHgo+XU0U/il/9uu0Kgm3stA39Ktg8yvma1dMrm7vcoUsd
5qH/NdsrIEy3EDJNYKkiujPgjrCS2Dfbp/nn6ZpMJ2Mucx2rKG/LW5zioXGGmzow
AIQcQNiz1yZQsbSFp4xwdB5zArVcrFZtrKOmepio+rml82CKO9bhVDTokAD94Cnf
THEVxMyDJjLiqA3+aKTmmL1cD7Gn3yujmVqnPSCi+xCuDI0gpDCFKa6vNQp6GsuX
/5P+PpkLjPQCz582A7soiJU6sglj3mZUOpFQ2YMW5Eenj1ri3Q24fbICoIsT3aAD
FYISwpVhCQEuak5XQwUWMemu9WSOuoKRpiF5oMBRN/MDp2JSk/EOiwKUAD/QRGhY
4X/rUNKWXQ/J4Mh8d7KOABuGZ31Ps7ohr6fAw4fnzbLpDEDv1VPVLYUfwR5Vk1kO
0RpoNcAUQZjQ4JXxB5QkSSK0L89RYjvw8u65GMv1WY/S89DHU9jcnWcypsardIiB
lf7Re9esdcG4bcepBZtflLqnBP3t1LwaEIwtoK7qoAfbeyWpufpIvcAsOSlx1iWA
M3CTcHQ/uhQ+5/W6CYkNZE1bGaez0TXSX3lmHhdVayaRhKM97JQRTcm7zrGlh95L
elqeqFMLRzNo+yqR7aJJwNafIXFfG8WlNWWC8E3o8v+4iODPfrA4DGH08l0CmHOr
sNXmT4T6iak/CYpEOQPkQ3Zx7KdAvLpKnGOLFq5vttjLy1nOpXcjICw6zhBZbpzi
PvsfymIiYJZkSnz15QddLzsUCfcPym9qJQf1RiMVe0BCW9MB0miJ11pgakuPDxRg
k8fXrOsNIm7Y0noJ2s/qFdId5KXVNWB+u5JaHwTZsVOLO47Bd0ziiiaOgm4ok8II
m0JHoANBBj3RB1ajjvrfkX03YkIKpwuLKlOX4jp6LOTnB9hRXYBVzlVSt53sys8u
uD9hKukYUhm+pmchBxWAbxysIDAdmYkBKcCtXXSTxvtbCgNcQvuWYxMY8qfeFUuD
yNui351v64WsEqKkbW5r9Hug3SOj/JLnkFXXTmVVvdmtxyHrVDLOGwCqvz3kv03J
3lfhjNaW2l1XOqldj3kRPDyPLG8YRBzzVUYz0gqxoTBUrPVwDp8oCFkvB24/b5rI
i1CEw3lhgspqkI/PnqM3iWDsIApsxarjPVwVN947xW+M7f1wRFqauFoZybYLwAq3
lNjZhB0DZjJzGvKkSGjffNDjxJ04+PiblV9PbgNzobdsD4kw9qVmpeuQFoyQ1ECg
RTrzs74sSgpbL3tjpnd7pbvTjEtQeS90qV4DZrtQYvpGw22DRLGJDuE8GSHIJ7qU
qa0h1H5Ggbot79XKvAerF78KsZ2ePbNVuu5qRDTfR2xhZAmJlz2I/wh5/4NAHnN7
i1ekKpnkz+aD9Zy3cz34Z6tXxMKOD6HD6w5n22afdJEC2ZOTBchW+FO0Qgsy3Az0
NtExV77FwrVhWt0TxjJ+5I48whpgbMrrrnydD6SgsjJQrsJOdrkEGL+dSFrcnEdY
OpTzzSVUr4hGJt2ZJ1SXUL6XwzzYXFGXyydppQU6TBErPWstXHcBylvQmPCsi37G
oTSMr1mkWnoSUQVOJOLGxMsAq3Plt0BfrCBzUcQObSMpaMA8o87Nao+8uu6jQGXY
euXu543/QysRHlNHbjB6VPef7+2x/2jfZBbnK2I8Us6oX3NpPuCcQn7kxxUQh6lQ
T54Sc7UK0ISZdWbMEEmYyD9W5T95oAfynSdoIcwnN7XtIm6zgRgcW5vaTSiMPyRp
yhYdUojUCKkUU8z6JUhgw8p+DveSV4loG/6HH12I4TtP8klUtZsUDsYex6HVBwiZ
hl8dTEruy7Z6rFqkfE+lbCizRyanc3loamVU3xr2cFaADJGgjr8Y7OxHyI3PhaQL
1K6la5bM8VgHAiFIeKCJUjCo11KPYxtk32vxMtK26TE4IH9jC5yvDsi6D6mIsADx
xtHOUMErHN1QwQonnUMzXDOLRJUwTcB3EbUIP9aivHaEwBnrFg21b5z5pQYqOJBd
/HfCh8gtvETwKhVbu6VYKhurCU2hUWcEpiCn/nawBh9ggj7C2N/9uKKV+K7CM1t7
EtKPQWHeBYIT6plmtWaatHLgF2UVluC7puO3f/eNBN8pvrvtq4qsaixhWbs5FhfG
WCpXYwEuoyPo6a6LAjXxPvv32KHrxnLDiyhEW+8u9izpwSo8qn66fVHGM9H6CAgb
A4wihsuvwhavXiQldnyt/DMieneeOzoBOK1wQ1hQCA1+AnsIgKPK/aAuDAqD+7QT
Qx5c8Ox7HVsZVQISW1GmzjEa5pIkZCnMysJ4KC7BObjDZSu/Iitd90/mHuK0QOhd
2BMh5fOKghHPg3Qhc4cMEac+WK9lGlzEbutI+hPQ3flV4/crW524EBhkOFEFCkUW
XamF0KHU14SC5Q8x8ygE2SnMrKv/xeFeVPEQHSFANgbTYTV+f3lEVQOHgFaldYUb
Y/IXwgnR2ejQOP034EwlwozDbxFTeEsMTjUV+nv/EINC2PVy6kpwrG+RdPuYlNCH
jE0M1HDBjttK2GP/vpH0gbsD2VhQxUZ/sm/7U2oAv7xiCd/GbwZAiAYs08/Nk1zb
E8g/+xDc7oZSktxcf3comxsPDnE1YdkOcHHh5hhzkjmaSHI5DGJLy3E7+sSuZW6/
7TX6L2JQWq63KEqVH4O5h6k583/SlQw31Cb4TTTXp0bunRYYyIMt6MPpCukmU3NQ
X1siphRbhAXNXWnFImy77l7NbnTb+8v8m4LnCJ8WygmiwuRA5bxXmVqkifcR1Xpl
n4J59CikpCwy3XRy/CmL7+phDTOI2L/jUMWK7XUF7R9ooI367NbQlIvHIcoSTgUk
zUicEWJ039z3s6NlT1TzOC2X0TyQzB7RtSIkWugFKB8EdITOg6YKuUXYxUDNBFb5
ceGh2VLMtDNJCz+jtwU5iKZ2e8rng7tkGq1ofzLBwxgqnG2iakPFqL0YhEn5hVPq
zrZL630xqZMzFnl2nB5wWEUSz/z6ShV69aslm3q+4KP/wqOef0q5WCiPj4TUw8VK
oyMu1SPMEL8R/zs/4wg3yDDUlPrYUYbjXXNPCYbb9XZTvXqOP+YiOHweAZoLsi1H
aM3gES2/D8bK3DYxDiHiy3sWZhBrH2oYqs7tuNwrB8jvy4f2xP4/ZEObBLkjCuSl
ZPrBYH2XBQMxbDHk3rghz6A6YJIlGuktDUACIWD4zmDsm1hNxbbBss7PhgBtaL0l
67IdVvCTdSdze2oMA+v2aLmWTaJ5uErN7Ndz6MBQavsPA0tqlUU+tNLI70XJ81JI
vwkruyg0WRGLGsLsJQjEQ4Slz7D2b46thDd5bpiTzwdmA+sEC1JfwyRZ92nLgVNd
SK/FQXZS2vzadrsIcyiHSiCjRpdFfutx2eg9wTTOMz//xTDNofH4qtooGQuwCvEc
AVl9qpksKTInh/t7yNRk6ZLMpq05k9Pg9kd1mUOFWk8HvprRAqIfw7I2h60OGsQK
qU4X5MKYQc7o8M1gZvSG5vRYc2d1jXGnA+on9LMedExDCLsaXOYbhM0k/Q+f88mm
RHWTqyvZTYP0SGiP4upFaZx+cbGVRH9pXQo9wfjUO1ao4qK0rV6FSWUJ3p1qXRYa
bhHcaA8ljcEQ+/n/iODathzK+SL/2J1Q1zzcp2V3qgIul8vGDJEeN4rABGq1NLkI
6Y69ZAazhCzPD4/5PJQC3wLsauSYv1czf7B4BYaUIEUTL8KsLZOdTB6t6HDzuajz
KTUaA30P0bxr88482+cV7O18xaz1FeGaTzxsGe/UQE0U+Lo8ze9uFKWQqpW0wliT
U72JWuOl6R/9xPq9cupbBlAB5k+bqN1MjamiheDmKfvyPi/uG1Lo86vTaa3hHGAD
Pkh/IlgqQUqmH2KzZjO9xxLnJZ+qTtV2KD8BV0lNS2/JC6OGLSEEJHCjOEuZu1D1
/GT91krH5T+LwCMWKIBQoaxQQfKLZ0F2qsTQuWUa8JKRtghZ2X3eL+7FCw75Ik+q
3VHWsUW+7N4S4r5c3wecD5cr1m0PdHbClFpIDire2XIy/HYDhNJYTSJWJjavy5zT
M9cmRkH/siX0noKiQ30u1mCmZJTy6JlXd1TC0MKAvchlKWcGBxAvP/JFdhR33Hto
Hi66QHVF5mfSHkikE5pqmoFriKx3F36hZs9a6V9KRMe1SARh4Bb06/VHaE/aXZ9B
9f5Reaea+3saZBJ8huGUEv6KRb7IQjNOjWbvgJ2LKteaJJ1E27RAjkEA2Ohm1SxL
Zt95RI3SNiG1e2Yq7vIbDE7RElfOThz0lS5F61r/BOPSxmffXdtxzzSIpf98EIG5
wmhhv/pWLxI9Q9RxAUbGwUqRtyvmeur6IFyhO1cuWF8540t0Kq6Sb6NAh04z6Yw+
jA+gz0p8fpa9GUXPVoXkhMIVOVHY6dBRNYAJ0chgY5CX7GcZv9wX0+lDAcpuxjUD
UXIu8XtCANjhdpW2VOlQL7jsMox/mS+cMiWaqx2RNZVtNrpRXUoh/Ou73NdMMVil
zh6pVRW+Iqf+vUbTZhAuHatHwTkoUK3oOT3F1VlCEzpopoG+gr66oYNvolI742Bj
bVbKe3iBhSQnfJRVjh5tIprG0PUqgGCtePjibOmCwQQFcT99QwrsyLeCVcMBwkMo
tso1Grau+wcqa930Mcs5lzfsHku4cKbpwWgoglMKcVl2Aw2gaTtT36RySopHJsmm
Q91aQ+2V+xKUhuL3zHBpY21QsuofuudBALKSucU8w/ZA8Y5Bcer0LphFGKb34+HV
0ry0mHbNoiZmCgRtCfO6SEUjOsQItHNcwLIfllyoD3MOyUHpLCJRPA7K4Mb2TbPS
+Lyq1GoAP9mfx/+OXkrt+p+f8ygfaejIQVZLR9nPY9Zcy3i3USo3hCvT0wf24C6y
zf8KXFsJzmWfm3z7LBO2V2635YRw8Er2F62emcL9hbd1+4DrqyQyA95jFsIIZI7r
VE84FWi7l8MPgHIDBY7iIo5tnWyUPEXkN9ja2GO7p7mAe+hbj/JpKQLLbJOT4uke
+26V9weZSHRj7y07E6qb5RUwoZ4DbqAn9dNKj7HEQAiD6rTfAK+C46bCSJPeHlo3
a0ewMukOxW1uMCXNJmqlj0jV0auPhNQkd8qscmZnD7ZospePlwfghzuYQ9zgW3qZ
psPZjpen2vH7Z/KCE2Lj2d46DSmX7VjIosO85fNNDpvd2we915mBW8bAxq0W/V2k
7CCS34f5Nm7Dnl8H7IMUCviCOOYdSEZS4DbNIt1FLvghfeU6wE89rWr9g1zaJZN9
lbaQlKPFADH3TH4hQ2usfLcR0zNZfqUFejCQQLwZlpuGiwC0cqjcD/9A+vKqD0BG
5w2gXZFBT1VvZLkXA7rtodOEfB5T+thqgSOR7ZcO48eOZTMg1Oz9fq9hI+RR2jOE
LNar4Svgb0aoc3WAT7yTmjqgf4YTnPNjjBbqnlTs5SLP/kPLoasXNlrEu0Yf9xeZ
qMhCPy9PENwVaG4DDQze77JO2ErOsTULOgatvlHe0yB5bim4005Ql3gKZN3NCttt
Gv0WAfXYhHQA54V1MQPqEqt/+xTY7Q7fD9RdgdbLNYZgobiEnOekOYZ4qzHiZLEH
g5xSgo1g6zatnHYV3z26eqB1htLqczV1ag5SYDWnyRPddexoLznxtC5y23JXSpdG
R7ijAvuidLBXm1sUvhyeVyWu81mJKE2RUKN1k2pQ93pqIAQAWLfpz04wBJlqCZQs
8I7V2AvoKKsNF9JzmSDjIJ/xdggLAxusKVqz9lcy/Ih/1oQjXVKGlTpxBdPZyfb3
GAYbeGJWdbQjnV21zBgbPi7bsC3mM8qrcrcdQnnodXRWui1cWT+c+e77Gp4OD/yc
4/M4BGQGYrsHBLaV0sokv5RcHF3FjvF3XyAK11Ayv4af1oZOuETzq+0d4l2I5qmp
9WzzmSfUUKZAgkJyF71r++PIW5oKnAsvcnbFiseL7xa9X1Y7/z0YvmzoBvA95+MV
ux5L63SYxojWQrXGsqkpM3+UwWt6Wi5CCh5WZGCcVbctYadTyuc/stgxjjkKfVw/
2Bswg08SNCcuLCSsRQ9LkPmQgZGMO79URAqpAJGOIcm+iLVumPhewsWId9bsDUoE
2G18nzm43GhkuFj5S8cGZDALp/QkwF5VdetAwXBmlkZVtftPbXd1JLVli8cRt8O8
WMd+ailWgXazuJmkKOEpAO5w1sGwOyqaxiTYWqrWoKbu+IdJ7dYe52mJ0kReCV3r
rHgMzuM/wT1AFr4IOmaYHmBq1OPM+Gxi/SqY3Nz6UCx4THAleYddaahuDXlSFdLi
EbDkSvX+PO4zQvuLmXbpPwLWNZmtNfTq+W7EB49eaffLD3bYQ+4CGQGELDBzQuSy
9DnjYCfivWV/Ve12CthSLn0PQBFlJUoUYuwy3sz1VR+/3ndh4NdsQz+q4+swlTcf
oXLxk/UEIyM2+ExlQ4hpUD7hLTYSCAW2q/wQLI4dsrz2DIkgmmrBqiJIc0B81/f+
MrdXpr+7SQkvVbIv3ZY2efpGWC9C9zsDdxStLyd51Pb9mag/44tusKwkzoxqlTgl
3Qgn3H/iOofEnNUQThDvkeg1kOQAtsGQS5KFVnuY5QJoAcg8eKp4ZcKYdFcY8qGO
i89ThhX4aiaCK7zZtdNjl9muactpU6y4hTZjKNAoAWayMRtNrzRDbB6iHJPTY6/7
STGaD4mXEyykd5D8BiONOYAX5CabtTA3vYh04+CAVR+Kw7mcrLK7gv6GzDWR3EuV
HLTgUymcrZjg1L+kWIbAaan0nvnF+U7dcJ2FZeCJRrlwILDTi8iiMOOQK0cKaIyZ
LMCcSRwwFxfkgomX1oLz+D5ymyMwIBr6WjWGzxE5jdBOv37wasehjpIW69Hh9h/W
oQfmfFT0g5vMLpQeJzhXzLchCgD5jqV0jHU7P1oD8lCbyvDY5Bcj1Drbt2earvno
dhsq2UjqiXb2oCqbP/aocirOCSd5ywXlO1IAYGViZbgihJFCUoNduz8lzAeX23iN
O6Eph91aYiXEK8GbPVHJf736gCP2sTuWWuRCeCFOfMzkBk5qVr43PAvt7UoidvD4
YRV8P7Iz/xJVDV6JOT32UJHeugPSLv2OmeVwCB2ToXDQ4Zf+sTJPXnUiNez+QXlC
ElNsrD7v+Zt/LByqD1gGk+bjshoreR1xpYnmoGAyxKiLAPcQtNkLEk0ri8U5Tc4N
rRFdXq8kBnoFiy+DjjUeucTMhiQPK7riyyUR/8llVOY8T2YTOwiSrOR31UGt5AAF
6lNTWdXHOhYAmgmzoatlIADntwacH0uxzJ+YXEy1ArwYCx4TGgvDyHWr7I/qa5Xh
yqvYUK+bKBHl2A5hoFX5NgGYPTacXOCZCvbTv+9o8XXQzmKYECEByg9SaKxadC3+
/VSJjw/oAVJVBVwetZN11nahVZ2fEYrLEv19zs18YzRP6pui3m3toIbrS6KlMcHk
Mo5Ls45Ou8sAe6yvtLKJky854/o50+D7aJ1x+4me9QQCg93u6mW1yxIvxPq6gMCE
H0cFkf4kcuiB3xE63LFHxTByZEG8KHbiAWnVWl3YiL5aK42VTOH6g4V1Ia8wX7Hf
7PqxFk+GQ0MBBSm6JIRVvHQ43r2ssEeM/qIR7NRLcSefE+OfmL3LdSynXVffgMAs
2gOzzWGkPdLaCuk8GemwaIE6tqMq/JAbsXHLLKXDaLEfAuA5BiDWegyxsN6h+wBR
tfgNUMhQpy9FQrW+d4gswfWouttuOcAkT6J1hB4L392xM0mXuMGw8YxRMBsgpBeC
3awKDHz1lrzqOSJCuxZ3+gfo2dEj2Lsjzlch64tY4k0mZqmjJEX4PV9E+ow2w8MD
myTM6RDWxDRws1OmWVzGthMu5wF9VjmldTK75uUK2yullU8c+HPEK6GG7uMnwHo4
wqhUiSs3Crc6Qlk8NKY2TALkJHBxP1m9n40Fp1UHPfaX5nPCt99VN5ILJwKf/mdU
NGh8h28lyiW5Ua14smVio1aZw0bgVyDk1pFrwdSDZef70DCbVLypuRCMBwgi6Q3z
kGLKz/z+cpAMMzZuYiK7oSkdDwu1yqw4+PNl/PFgGxkn0BHeikvuzRsCVOy8qTdt
53d7QQj42p5oTudgxe6HOVp4L6qBDYKRug12f/DM+888GiknGwHwSC0cUPyk0uIe
SrEJeJFP4M8dCdOA78GVIdyaACUWiJcLJbupMtYqTKlVllhJMdhP7qnZ4xf34yLL
FfDFH1Kgjwpq3sAiVXcQfBdfizzNvpmVVrq1sDEw4ea5Vjezx2H4l+zjxZu22jfF
xK9dVqJ9W6k8GjDcuxR25CXF4iLVjAhh37bnIc2RQr+G4aA1hsAddQ9NkJ4adyd9
IIzec49nbPxRpgaPOe9uYkVAEljChr32TnhzhR1oJgSn/jfX8ykg3pbMdlUnrvhj
RuwjU/JhJpxP+R502RlIbsW95dNMQpo/zQ6WNAw95cO9QDuEVbtmGw3BxTKXWhVB
bAg4UXlCDNXFB91cNgYao/DIfpCUozAoFSyIYt6scwynoeM4vzpOf0heyO+7KYWY
r6n264BfT3fNSLvnhptOdv7WkixPOgPpObWPAmr62c0Ti7eCcYM54LVdLZFnKoQ+
vTOPw/plCUjfQRmxrY+Ln00vdu85a13gKjLifdWU8fKOJeOS8UtsayPZemp7Ypcu
Z8kOuaX0LcC8ReIU9GMPOu9/qRW3+BeMwIHseJB6/9yePky6Fl+wKSnChSGNi0ba
xD1lUXbwvsBQE3UUF0oDM1Gx+BBSSzC0WFoE0cNJiVJ7G6yRi58C+TzvsK6qkWa3
s5P0O1/OM4v9hvyWTOmCPhCvg7nH9ZhSyP9iFM9YLyEljsm8MS/r9yv4flcp+8SI
ueh5zupCKMKR5JygokcFM0M+/ykrOOzZlAVUDlYpvpyQI05V0MxpSu24Yw8qMh5t
p86lFh/hYtHw5mcQUOO2v45bfpVfPHFbyUR66DdU2xZB/70l86EO8qH6MTGsIzuC
1h4m8vq3xYdGZchvJBJddb3giYi0e3tLmCxajOBa9wtIrgSN87JY2+hjPwG1ERB6
TEkbFYYCJRrczHrSlIN6yeh1UbaQ+h2nIzhESkd0cutz+C8j2y8Xs8k0LBaEmebh
P1ayenddYl+m1vjeNdtIKF9ejo3kIlkdeGNC1sC7qN5IJUKUZePwaBX3ag5QKBs3
tItG4bHg+R+uRzxSsXycWUkDGj8BBR9w9P3zHQ0Pa2MWxMeqIydZg5Nn9qcmjdil
cxw3q50a4pfwlSsVLi+bF4bz+6r/ouGmoL9A1cAUbgNhnytOxMEk2BLKe+xfGMC9
MMcQy3xsLQQ9jBf5oKLzPw33YhednT6lnQpva+o3pvNj2M7IclhUMCIazZpia+Lj
XBwJMxl6cpXpWnLQ6x1rQ3NPRznZbTT1/GBhY8L1Py4F5QWrgE8RynL9WyIWqdIC
F+B2unnkw0gRMdQVho2E7FHsED/qSr+iDSJtW+AEjWAtTRJPk+8XQSN+oYb7MBOw
338P7zKjyzUWuEjsBJ32OpptE3x5BeDNd6YuKTsuTkTJSa/wx2uAsC6MplA23PKd
+WBoZjwCwmEBE+UDLYtF2W1dxmqkpXhx0YoXb5hIM0iffVb6otTMPpK10TCoNOet
sJoJhaspidxXZZvS+KD2UAhRyNjKzBjaUEbMwhfkA2HFMEH7iP6xYLeIcZCg1Q96
DXU+rymJVUOPIZRitYSy5PAOU3eKKeoSCpGwHF4vJO3cnAHeBZIMNrqP2xddoeFS
ZvUpknfUjjrGbBiZbGbTVQrvTBnH4GgTOzQVNDY/ygysxHfjZrcsRxzOcxls9Ave
fqxoh/IVMJP7/RrEhMhk7ewfEXz4wHXXKxpA1QnVkd2H9qv+nNh+AkOz1ER9R9JA
eOoi9oLVoVIh+Jyp1jpvuC1H9YHKfcH1g5ObvugyJ8GlF3qSCB96GOGd/Ocm3wIJ
Y6RXPsfwZE6bhuwwbSsl4vE1CMUOyL2Al3c14yveT40I4HfjJ2RYerjE86uNVB1W
A65ZsvgzRbR2QLZ3+imhcj6l8+ly9fIea0LJRQ9X++52L/cFzvn+jWeTsobbIuqH
9krEcl/Urq4ce+MyA/3YVMcZLeUIh5yPL0MRfcOTfdS0fPMY8RTQeJ/cHJR/vTmf
H4/+VleOborWt7yg/D3ps9b0XmBg9L/o41nRC6NLXhOzZI7zgHeSRGkI4LkxiTmj
iAaSHOXoDdZzxuV+ZpbHmAlA73Mg8j4mBD1mMm0cghjXwbefyGQcsemZCTiHvUig
AUX9FiwAQvYhWQjr4esAP2Ab4ZDvB2FDhpgaY4s5WtnkE9GAgocxHBU5cTy8/RGv
IgFWsbFvtGDQ9qBuAnjCQyIUHFIOT+rPO+lvC4WncmZKsedqWDIqFsbyt/Cz8Mzo
iPlLFQ2a7Umk+pkKgFEY8/1yYowAPDsfFdiaOiG3QBfIIM8Ksz2XjcIlErmCYgcy
WPhpEU9yKWooSNTQBTi9FIsdrQ/Y2EMEsyiK5E28u1zSgg1lvNDJjdcdnzgNydHH
wPAe5Wd3Ij52O+LoVpghxof8WVNQaDnaosP1cAHy8SZnXscfEJzHqyaP7TiGLBPI
WhAqInBIqVxUljn5EIvg+Y5Tc6kVviBD3gaKgHUzkKxS2dwf6aVANr2rpKnDX7Lb
/TMJ3JkSRS+IWAacGrO0+w3f1ksHB6UqROJNBmH3e00PrwCLwNJypNW/hl5PFBzg
iJ4jKa4AStZvD31ScTbijUz1yQJP5n7api4XPP7yE6xPQt3a8m71ZuUi0U7rMNhb
LU+y3AjI0NB9DDhWuK23smoLQfewj5VR4CY+W60TsiMCoTpHU74zePZSJffd+TJK
ETvnWBnhDnUO7skNyrwQ/Ed5PLS+jWPJddl85LGbYyU0vq7puoydrhhKj14MiIde
C9InSlGNyEBJcWNAZgHQidyFqNggaSGxCQbOKr5VzSjvBPua4dOPiFlJESnAMgVD
yYmnAjuL435ss+Sowt8POhJyZVj16ePBFR4IIQTqNyvVM5B+4k2Is3e5CiKcAw56
9hcKs19nKROoTKyVKG0SU43vQby/bIPGozOlBO68mQ0x582cFl1zTpt8cw42A3O9
bYLDW7k4k7Ny+cq8nzBYvoVoNRLIRMuLLpvayziED8mtnAlBqOyA4ojh1j5sO7fX
gzm7fC1rMlpqWgR2VL4pW+aEN0p4r5OP+C+JXumi0WCYUCDaJGiThd8GW7wHyZt9
3Eu4chhVGvAdTQFBN+rKvVBUwy5VAA8V/C/DTxM5roUjr0zpu0AUg8+ALBIj323o
qICwwRtEC6GzuYWblRiwcS+T7FPd0VqdkOzs34N/N1WsqNFw6+DikwHTIk6tC0UY
TPr+m9oHXFn1ECE8LKNVXu1szvFgf71lRble9ZFc6A6ZOBFGcmfMaB8vwlU0MGM4
fHxyBVHfOOMmoTYWIhP6eVu4/BfqIuFaAmQtcnE+DlFPz41VxJrxcLS51sZkBeO5
gHX4Rai1syPTy+kP4BgCO2iHpC9LLx6BGhJPHCqypRgywzTPW3cNHXpIZhuf5vX+
VEXAukb5TsvoBiwOt0e1MURLaFAhmI3F2GPyKsXIzGCPG40jo/YWuSe3gJs/ZCxF
du8PktnYz3PVCpC76WtJjBfONrAh6xrDu5dKjtpVtklHYArGEP6grbLh3mgGv+R0
tX8HOzkFLcW1FZ0vB7lzyOO2jrBIvLB68ydnBfyfGeYYy3MvKyB6TBjU4+6OnMFj
/4pekh4uzySGiiZFmE2JSJBXFh6VmvTWjs9/pMeOx4bdS7GNLqcli01wHh2has74
2wlTPvbf6iYd1QP0pVsz2AwFutsE01iHmYsESivsIM82GZxrxV6S6PovquB5ZFxc
lBLQq0gSvvdRn8+PnLr7zcCCDhZyD26MSBMA/g8rxyXzMEa2A8o3tRWDS+jlwJ0q
BV3cuVlOZxoYhmfm5hnONmGUqf4AaxB2I5SKDTBVIEWA0u0nOV4yN+kj14eXptkZ
26utfNqYd93Hxu+gUGxpKtrj1Zz+K/9/fBOarEt+O0ZuP+N8JUVhag76mEr0Hs2m
v3rTrclciHthQ9k3ApsWJkKZRoPU9Vl6jGp+P+OJLeWIOYNkwOAZb45zr8rUfy01
5UHcPlGMGQFUv7uY10NdCEwqJ8bSK1ntlGWgdT8TgC63SIUDXiyZX7hV90DvkeI3
DHyDs3fR6q78scN6OxrJ0XbTrh21mVf0aH5QLu5ckIJmEn+VYaOssQtTlA5kz10G
Y+OvlDdbar4d6IGD9K6SX2Xsm2oC4CgJUz1yQ6phHP20rr1HtQD5lYUAPKMeBuc4
sMTJMDpONchKAD83iHIrbKmk3BfLbVvlrrom7QhBAxYj80rvNJVdLaF5KoyENKkw
fl4k6FpHW/o0y11FMeAr8jlFpdIlUtJX7Gie3VWTjhOlCLo1tdl223ivzpVP7Xp3
OhowRBEVBDZfQDqxpRGPv/cP5YubatjSiSJ0ip70Bi/VIYSWpwTDbHOD+3X2Sj6k
/kPHBogIKBrLGMhpV22YCAmJlp+QjkZsrqBVc+7Vmm1UW7nhZJWTR7sZwCeOB2rP
H+L6qjGise9WaRhjlLJUpDwugx/BH5cG2HRsFmKMRTLlPfiDFlUwfKOllPAKYceR
W2dg46KTKLpE/YExhtrjSynZFwo1mXbCJNWEIKfXdIN5pWhPjeudAiktXcrVnG26
fHsTUhSblosnSez9UVeJ9WFPydwc4MCr2AFlVsCZMDyhAnkTwmyK/YDYXoHBm3q+
dCe41pUXfYrX8I6qwsUI25sg5F2O3D5VGFtwBL+R6tH3QEHL8iyP7saQKFy4qO18
3dQd4j8fYvlyjiuNnrsF2ieKnZQ4qS8USHG71WCYN9AcEKVaH9ao0dbVnqs/9aKp
MOgxpXRu6pPS1hF8pdwyJ+Dc0SeySQb+9P6nkBbFHJ/OUpm8054NX1zrfKZ7GgDP
MvNB+Ib3B6gRBkvM1abh8Q6H5lx5mv+fvFpuaois9XUEx84AMHx0isbJ4jKUnHd3
tzZcst/m2wotNbzA6ec4keret8PDk2lEeUMwI8P3X9DFmxF7Y+RbYGDJ0RS6wwkY
pYWR/q09tY/l//nFxw2HX0oQcczcmK8WJceu1fFct98RUdGnZiLote16QJxVXYSN
6ldcpcPqXV7monO4TDJzH4aAHbhd8Xs5kl3yDUT9XMjZZzDyTFU1Z+PRYXOzmRPO
PmZUaG5pBFGMu8i23paXH05Lnq/C0rexicQYtb0cuB1EZUcjV5ODJJYQNN+eoxl3
S5A1G2/UEt2trfh9aWVjlebSK/PVaSEC0s98SB1BcphA2O241dx/Atj2TpA1JAcV
LnPnd8lMk3s/id3M+WhJJp5KG8s4CHK8zvHtHoXNSeRQ87kwDJNS6P5W3ciO96u9
KJOpYBSVZ0b02KZu6y8ydVMo13uKKKyJryTKbuFzPiKDfqt7odCtcdDW1nAzAF2Q
SUqPzX8QWSXgEHtdm64DGo+UxmFL7C0KFgOfLWwTVQR8JojpvROQDybDCs11A8fx
xNuOjH891fFVK2eVoHT34aaVixZBKwcNs6OYljOikPZ17xZr7urB4xWnizELq8uG
hVi3RHEHXaKzYR9pHON5Yx9OZqkIXIepN4xq5ICvmPc4JPxihC3GT9ra/iP6ze1y
m6EfTh/rXo0Y4174b+VJjUi1SQW8SHyB/jmzZfjb19zf1cUr0fM8aibcS9qMeFxc
pL7kdS2yNcEe52IGTHHYZoPVDa/xos/u3ErjwsOramJwfym/2P2bNFTtNbU214G8
V8eeLQhj18to052sU/ZayWYrwasQj7NPcC2p19RyoJ01uC25il0nPajnFWlQLe1W
IqZGBK5oRp4+jtwHpIR0clvmmUfOgRuhGthurlHEkVMX0lxVs1roUNnj0O0G0bRO
Maaot0KyRNsh6JccVxFVNhm6kgIaaW96hYYPXSU0Kj3UuJSmnCizgCKKoK2E6Pr6
UT/cwWGPlNER1hSwrCW58dlAPWy4KWtw/o+Kleeyu62iCt3q+y9tNi8YbUNSSEQK
5MUs13v+YiNer63ymEIIEyBrM262YQojwPStwcVzcALbzYPQ94XXwXhwTVTr2gA2
QDtuuDhuzbmW+PwJGX1UxTPTNunIjEMYuvA0NlVzoOdYWNP+AfeLMRGD3QLbVBk/
8Wq/C//u8hArFd7WeTWniDL7o9TggRlnBi6TtVYpReSpzpmFVPdJAEKeKL2912ql
VxqH6E7jQziTKDrwzFIjjus95AlXFvPemqbxT+wnWcQeBozfw8JaWXb1Q9/U/ayh
ozutirUs2ObTSSWh4Xz6Vy4NtBoy/th5LqL7oMdm6Fah10pB+7MbUvk49W94OUrH
5veFqgxbnLWi99mQUeFGc6+YjRR7FVEMM0s8Bhe6sNVKBXVckWDYEcIRF+CoeEhW
o4dRk9zEBKKCH1jKI+jrXwsI9ulyS939AAsQkIj6UG/VawLynxLPqsuzQ+SIkGX1
BVUhtRme5KXQY8XIqbnHYtsKaNDZDLYAmc/vSHiagZjDugbSCTnSYgw4XF/0V2KC
VfnYUda0wwP8ckugW44UjQy3j7t8BRiF9m0FnyxeULRuYkkHmxHa1Leo5tPpM75k
OtwZxsNdJcBjytnq424/+2qPxhLLKJJayZP0n5TBOhwXvZqOEKn0sIgONS3Men0i
VxZXyiMMQwnSEeOxu+EaplpiE6YRoionCKc5T14FppCflxbLm+CLKgv8ltQrx/p+
o0AdpZO8h+eb/0k9Ha6z5scJolWn0SjdnbnYQq0VdVu82XvxQl6/As+FbowVslSP
ntYUqOKIranVAhHLlUpH8BiKI6ILrP4gWdABqE6Z/AJlp425lIjJpAGifVbf1XDH
dTJsXRnf75HATaHBcvk5Dj2ENtyqFARjgXyvGZpTTjazIZvWkrDCM7h47NgRzoD2
R/OLqjPZv4WCODude6Xs3po525DrjKJ+ZKEZGywyvMVBJwgfOn9DIE2H7sAY8Lof
uoi5sUcjec2lxo3ho30gUdp8ECL2I3l3TYSK0ZUg7ar5l6frJuL3RirMYf8LwSoz
cfk5SBTXCeSabIgn7RJ6KM/3wgYzGRRP5T4NDco5B7qEnxFyBwYOIt6Fbs7tSAey
6S6cBKm+PFmRRqvd5i/DdE6+s9y7XcG3vW+NcKpaOeyCk1bYqJV9ZIVGsiPHALdV
mkB9XPefa2MAiRIH/QSS+PF2wRV2XYqz9E/VFsbJFvT+HUQwl401rF83ha0HJhY7
+yJnUOU8Esl3yZezgSEZMlCi2rNY8DKbzocJcvvPM/Bnj57Hk7ZR50d76b4hrZD2
M94uLWOZ4zFjIXHlml86M22juIqHRPO+On4nxXrsjQ69YN1sYx5IQoeJ0hTgMRq7
O7rYNby9fpwa7SBHXTRixifcuagcGpCVZOM2E1tFL3ZZW92xf6zeVh6iyDoMIO6R
Oh9R6VOnirbHlJXrPMWtAf8PEJogiqqu1PkYXQuym9igZvnNasJgocMkGG0L2s9T
39e3QSVRrZDjKhnUdb2mF2aVyF95jkhmaUkowo5RIuBbzA7EK6rbVq2K0gZR5a1k
l8Mmeqfq3d+zQXEv1mm+hoYnCaHDgs0Aay5HC2k9Aexy5jjSEJel7kLTDp2qL0HC
eZw52iCktAx//oktBN8Y8JB/DKuWqGla1nlEtKZnyuQNrgr+AVxvVzMzzQFyY0t+
igwJCM0TlWD93NEVaSulXx/UiJfv+8LwlvHgyFGT8FWy7KdZNw2DsEHRnS1Ai9l3
VHJ70VTU7EIUjjuUtMRRi6iprpvmmBNKM4o+6RhFISKAezqgJuVLqBKXpIUPvhsi
odG3u0KGciqolI+FaacgXpfSUPIfeQ1TtpnQJRxo5UXLlBgMb6u4A0gEroeLW/yc
XAMCdtyjr29J3EIYZdKFiXvM47L5/NFuJejTYw9vy/w1fvKgPJPsH5duYOPp79Zr
Na7SeWZnZd+i8uJhoJerkD/BxJPQNz78hL8P5tucsv69Gs0tkfjPBYxFTlrBI6br
7OrTyT4Gknd5jMxDFxDDdYjTwYD6db5+lNGMZW6zFaKWd8C6W4mYxqPXPmgBO2Gs
h0kN/rQ4sDYv7ow+30Se3Kr0rmqrXHhRMSWinX86fbZ6gL4h2PJe5EI+jqM1OnD6
hxTJPtAWBFDZeZke83ljHXYqbFcIyjHvyzQSbI2+KVXQW3qCIZ/D3esfv/6xA9DH
AVFBARLWuwag7ZNmhL0fIOEIjVmHyZmtBtA8hC5LmViRRfBhkswz/TVFTtRqlD+k
6EtO8eFzB5a4T1xfCPkrXIsEaqOaMLSD73kf4n4JITnqS80yG5J5tOOiJUMuvDxL
bQaqE3fHbnQ6IezEDF8oz1ebKF9kX4mClnWPhOKSHndTqenS+KnU2ixDXeKndBc1
KawZFRjdCJpmVo3tOFsbEEHA1PUHcE7Ji3dc4rTVJXTJBf9g21DD1we0DnMgHtny
3/6rJ2l/ABL353GgHIvEzY+Q/r/WtNi6r+FpU0jGZeaiB76pywQua1OjyGoUkXbv
rE2dJt1FppXik/ATIzrOm46EP5qDgsU6095xwd2njQyA5yPV2Vlzi3kkoDp1zQDR
i/+wupXoOOUXUQDx8u1BXvkfd7zaPZWEBoI2DN9iww2oGNeVtzY8aaaK3JXwYIWr
vL9y/BdiNhz4MRfL5Uq+gUaBcm+Bsbz6psYGoA+1aP5AfBTABdpIif9N7+aFz2VH
LeNishH2jfVDX5nJJl2BRJRmgCTisBK0pzj1ykMUXQoVj0az7PddrwVv+7GUWC++
tILrbbLoDG8dM725+5ejNHF5N3TmPf8QiB8VaQy9ZhUisXeo+k2/qUShStegigBD
bCY62qoqpI41QzvkEkPPfcG32Co4umn4lAd75tv2Eirbqg0vCrTTC5i827LR4ikP
/KIXS/CsfL1SCo1OjQRkuXDP0qbJ5cqB44riWj7UPnwyPI+o46/e8IbhZBh/zDF1
EEIAnsBLXTgGi9Vl1MTfw3cJ+x3W4nfnDMhWK+tJDRww0/qJgUwksWsS8mS7LLHw
fsm8GIr9kSbEo4gWct8RypVVnMX7Hsow0K/7UT3yMjOlg5yklCOhTdNMnO+IDZbv
VG6SaJJVdzssLhvznSC4mgkzStDVdrSapRUrxv7lWFLaz2+xPHtlTCSwJY5Gk56T
M4ZpctWqBiTVvoEc0dJDpSSnRUElN4CPPoc4Gwna0oTeGmLFM4F+qjMLum5aC2MR
52OtnCVuVJYrAqkHSHwpOnT2cHtit6mi2MKwajJydVvVO3Ghupa1dhxfNSK6kCRf
ujcBntRmKGm6q8T0n9vkT36BXk79WLgD8Ji437Q0Rl+gCuaByhmpa+bqCJFyHsUa
8v1Y8tclgGv/U0OxGjii0S3VkBHLLFt4L8SE/Na5D9p5kyrmC1HEEzUC7hDK43GC
hQZ1Xk94km1850kPP5TlklYmCDIazOnEd76UhJa5tlJVXxY04Lgf/WG6BBQ5BIQp
18wquxq28v2A/W7/7BR+PTSRA93lFFWThCDxEODLI3+MP4ElBWmiEUIPfYHdfZUH
cXeL1XIWuP1ZwBlQO0Fqg7FIWZr2Qb540+wCxMQqBQ9Gu83/0A1qt3je60eLVb58
kuAWiqxA5RhI0xbfJ/d6CZmeX/N7yu0DmQ9bDI3jeTqQ5XWZAW5zKE1rXrPJg22Y
UQTkYGWlSs9LjqCoe8bCZIlgbdJvq2IuLDtkV4BdAueCmc4ikDzoCVc54e5QtBqk
CJpKYXcY2YU2xqwy/XPaw0lMpRPUAzyfzPT4nIpoLypUxdh6VFrDSGtaoV0DyV76

`pragma protect end_protected
