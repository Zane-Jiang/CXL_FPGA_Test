// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
b/gVUASrOnX3ITZr1brylRkm11OEmHABoiNPK4l6JxR7ogsw5sEAFBbwvFNvJZJk
cz2ZaawviEOmqNpewLB36fLJ/9EzfazKaRrWyfVJq9w5i51pvC1E67+ZFu+W9PIg
vKti8NfSuQqwcttuurcXqUOAlWXf4HkvrLWqGEaMagQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 34800 )
`pragma protect data_block
3VmaGQrdAe5zzuCVtaNETSy8OwrxAm7H9HxkAQAjFi5Kr3BzNl6fWB9LLPcBHjs4
BDOAazfQXodzeK8VC2/bASdQOAxmwawVdjyd3wgODANuoKINUiTI/+AD0bYyob3t
IvPGiQlZe3haZCYqgCiGHCiHieAC8rjZtfaz+2Z65knmMu/edDUuT2wd683gqrdl
qCR/gFSGr1scbohykJ8paRG8Mvhykf8oB7P6b+4y8+fh6PrqYG4uuCWA9gm6tMNQ
69cjkMJ+o9CYTTrb+F7QDbu2rX2fIswDFBRDc9nJU36PlSR4I57GrGFbrc13/3ma
JtGZEfG75yGlxCpoLiQDOODDfNyfCvqRBekm9Tq/t3zQZqU/fIl3+Zc7BDZvRKvW
u+5WGYrdWu1TFdg5ypdckVjiC2MKZ1Q/SLBMNFiY0iTf8ST4LEHULW4ZkiXdqQ0c
pzU4503Zrbq07DA1lOJn/wgQLP1F5aXvU3Vt2u57SGzkwGh3HdOK2KCzDKfUlauF
EXqJEjhAU3C3pvWfBIyO2YM4Ggd5JngFUwXv3WmPqeu8gGdUQwOORZFhgQVqQZAQ
H/lQ3uCs2gHxzAC7Lj8ksHb37TD3xXxE5cF170j9jBPymGX9Mxx5EcvjrscxGdRg
xCHUA0haC/u+3NCxUGE7bOzgD5iA4piQXl6EDP2nTo4+J5O7hA9riL4HUjS+lLjv
1CYfYnwzxFMjQx4mJ0DBHdwUDgaxN8k9ozlcSDzACRsLxWduyTjzeZrC48Th6V0k
i09f9K1aJM1JL92ubmX8/Drqecv6X2doPHSzu4VJzvASRDLEZA7VGc8iF6Ts7+eb
YZXCl4tuK2Bjw6rvystVFGJZ1pOY5vAp8KrqpXm7rGm2ptZEjfW+jbVPebZIgvXg
M1e7mWZ19P0fHc6UgkNK6oj8gOjLKD2aRHeVGevjkqcVJ/+R3+8YHzR4Bc9dmC0Q
5OKjY5eLRGinxQNK9qYvb0eIvx/N/buJ2BbnU0VCJRfw7/+yoO5mim6Ukz1cgvya
F66aAex3XVmpldSXvEtxaOlyAPGoWCC+b5BeuutmXDjvL9PJ10/GT1k/mmvIfqPm
RIwIG6xD+ar6xEYOu3ashIYIbxBsFrJ1ocaG9s+x0AKbGbmzOxmQAwyWqBl8tJL9
/B2Nj9AnRXE+eNhErW28Ah1n3gIU1vq74Ri6OLp3Wrah9kPzGy6/SusPFTYBYC+M
frM1EJucug+1LtAvoh4+SCgelWjctyNlOPEAD1RLJQXxpug2DcD6rSA+BwL/cSYk
H8S0inccx5Gx5eE0rok5v7qyAha5SIm2M4nbtqXlhIcillTrNPcdyhvh/rFV+Rx6
N2bKKbbAekOqUpAOK8GTIwrK1SsJsqIMlqqfb80ctv0VNL9vpdyYrWpY3T+RC+xe
uupag5u6QZU8DunERVFssYPo/MhCvjrc1rMNp3C8WIOc+6rUxQdSycHLpqD+T94y
BY+5W2008BEZgSDhg/sx3Lm8JLCmwy6VD1wDypu9AJsD3ggZYWMEKpoTfRT5v3RG
TaS39QjkGR6dA2fq6xaPAOwkwqCwV47cGIAhEtaVIPqWd7CWkDay2TFLkne29EUs
LkSOPFNgFVoG/iCo3c02a2St5me0XnRo2ncdklLERYfLEr4t5ZPmCx6C9C0wOcXD
90InoWZCBvRFdb1RrC/MSRi1YoJYU6F3yEfcuvcbgX/E05FdyWcUu8RE4rHuepD5
8gJtyXD3VBuZt8ZimtGDFBZQecPXXMRubXUpxqIZSl+XdQEA0UibZRQPYwehP+Sc
yuwrVx1BE3JTqNfeZhvBpl+AQ3/SKp4vxcPsVI0l0B7bS5Ijbb7DsXe6rq857qzh
NqpiHjpqZca6HHbzplO/SkU74rERcVqknb4iSSvZMzE6myxxte8Uo2b3+32+d7wi
tNB7PvtV+tDMUihEyiQY9gSanNLMMXYeWBxU6qZnSP7m1wUjbnhYUz0naRDC7SBK
50AkHaDNmjp6dlqOnzGvGYf4m9S4eOBfHGDSUFgc5Zy3dkicUuN8keGw6mXnmurM
202J+XKbVsJv/twQU4aleeMS6RIHdGMygO71i7JgFgSrGi9wZKr8LYccY2ipHozs
eABzeyEtlpht3z6JIGiWkbleOJLtYSKsw1rcT39Ue/pjKdy2sXNcobZVFcVHdZk0
iTJPOlQQWI07iQlQtA8zB8mHaH56UFppowEJlO9o1FPrV9b8s5RmrA06gVH+Pgaz
g/69Sqv484X7YC1SGfzfU/NpKCtdu0OykuzHTqHz0JcoZqONT7aKUPo0ssxLEbxz
6W/pII10SWfoYVPj64k0kdjRtbE8WQjEjpjp7fAleeLlmjzoqXirPL53ykg0Hfhh
2ecBZB8DgQ3Md70GV6hqjqRFLdzuPTAVTRo8GRL/tdv/6ib0ReTa7lJz3joqE+NF
7oJv5ejohBTx+Jll5Kwd5YVawAjMWjPDYz3ksodURtNFfUAGn/eLw0VrgcCa7W1m
cobL1Iv3M+wwljpPsY1NZKit/gfFLv9lUv/xF29Mv+6cLUsaTVB41qti0emeOk7S
vLAScjXO4/SaBnXhnUJL1udT5kahum0UC+9gZ6egNmRSUFEm7l7vK+7GhvC4sn7B
eDFEjaEszQfWB+q7EQv2ToYKJ9xgu2dC9jRlG+NBug1/Cy9v8RCuBNQjYQ4S91g9
LmEJDzpAjzifB6Ibe4XXBy8gctg1Yq30TFsucLY8mVCtAOFSEoyb9/INt17AfWYZ
3c97ly417YGy114b+fIQFXmc0CdFO2Y0Z0T5gAIE96K3VUW6eXiLdCMJ1fUGoHWv
JZXhMd5W8+lvsm2HoYysEXzliLDUKCzFp32DpJbQfAYe8zMCzUri6+OmHoIoZxpY
U4eCL5ag0XeY1b57b6swpQSForQmdgHxvFDWG1kstM/4NcAjXedn7+Oblf2c5jt2
c77d1a2lrpKX5VEnJldJ2jJveXoV8zNnmbbNTAG+2iX4ne7s3lYu7+m0KhaUuPmd
RDAP2aFG30kqjQC4uiDXQr/p9NSdEgP9pL6d1M6kWegGmkh9eNDpt5c8GniNoQsq
MeFvKwsYxv9sR3okaYlPOcDTnkWEioU3OsMGDVb24F3mEGJwdHDpQiHO/NFBpzLp
cuGclxHApPeEaR/QZZDLnqdbJlLBAWntjXALQ7xYkR/VYFBO2psQL8Jta/nOmYJF
nWnk7RR5pjFr4a2AJ2A6vxrc3tkMftmvt4cKkIrT4i1EcedFsY/eP/SCDht4gTtj
+jhVaw5a3LHxHpEYgmedD9Jj2Nmi8RFA51ph9Bn+5DDk3g6k94EXKIuxobEcpClq
LAyXy40bcPqanmJX3+fMGbRrMgLUleNgJbtsSesB3Apo0sJLC+Jf1NRdyUCG+t9i
xMQCnCG6qyVSF0UXGe1Ks2IBwgIEFw5zuPazxx1rIZ27uGilF8vAgq2J6EaCBWh7
YZLs6WDGpjrVQZQu20gactn0U5KWTXrXInIq3jYhPpumNOyx7YGmAxKnr2MtpD49
9DFZJiyXkFZFYAY9H75st+DBHTwbpPwbehv8Mba8Dk4kQhWUBNiYIXE2ziOSMRK9
gHc99DRz2WgONIXP4Q9n1Dlxs7F5z4TVsZ66l5J1ZDHdIbCa3Dy0nKSZugAAl3WG
uJP01jhccnDjY2Of/paLJ9QadzZ8M9EprfPXkGY9crVYWNzKCYDFRbpTjAZ9fwuD
WlNy15BDTueiArybRthiMZFB34NamIg4dKvqAKK7Sx6vinpW8LRVjZcCx/v6bMqU
jDK6Ln0/XUSzj7WIde1bnmWMnnEoTvGwzXQB9W/VRo21Eo6HjC1QRT6NGTbFnW9+
8qXNyEAFgdfaInBTj8CCTZdIbGYNvrE9XNyoXP18bfV4R/Z9xXcmvaU6m2aX0nPT
lH1mKGnJn+fbpfUlqOGNcSdqvIVnrsYpA5LxO6Wh4y6sI6eieH7Qmx+Qs8eO2rF6
OvqIm2l2cSgwMcFWxDKudZKeWnWONjL2b1LuicwgLOR1zKq4tWchRt1BvPBmKoU0
bAiMtcoueG336HCUOCYOMB1IJKHe81zfmu3IzgfQWRAvtZCF0KoSr6SsUF9MyTgw
N1aYQjUUQeAwUJJj6/wgjGKecubFPjZiAIBYDLQ3fYMOOERp/0TuL/c/YwuF7TKF
rv2+c1gcpQjWAftmr5vpB9ijAc5OJLnhBVGFQE4U2AeAbtUZfnco1Et+lpUV/u4h
nnHyHWDcLFkxK5B+HQaehYSmchkSdTMN98Vb98LcoW6DQw/oaedIoUIuFV3P0aic
+U8KJ4Cp4X5W08DTX/hODJVo2u3FdwezG+gIveFGmaxoxyZXm2CISZEjOiZdwzZ6
5Katrm9t8qCJikVDUK09uTM+O6B8qPP9GmcDKLdHVCe0/cvLyblQaieCNEUxPRgw
3eQ1xPT5LmlMTLob2CjvDqtA5bWloZABhVY4X230HPHDj8R9hCOKc7wSwPy10Uej
JCglwZdIyc1QoZeDzY24ljxwojDK6wdti8T9CDaxq+xpm/mBbl1dusEDNTKWJ0E/
J7IsekMwbsOziV1uyEdZNa/ICCDj8IKyDpRXDf6SpSTJJS2WZOQaFierbn7pumAP
Vv0QHoLPuofL0Os2RRiggHAUgVxNjGLhvIaSKHtiMjtMRyZlI0O/j9G8fd0epnhs
3dsapmL4Osw/07r5hGYWzkzBzsv1iwCI3DXGxypoGkQch+gKyzXKMDnJo+Vy1mQN
Bub/GmoPPl6S3dRSXEz+sBHaAsJ8v8f1UZxtcU1M0K04vDZ08lONdaofCmCZFcQD
mHRW+FsSbru5HC30HJzyGQEf3VNKK5TbGxyQyhV4BJcXTVfGIBEpZNgziRw9cx0p
E+N1syMrMruWitzwoLy7/9zhbEN9AwFGYoMp1bMF1hN53Y7gNluWazCKglBZopn8
kWQ8+UR0xw9Iec48INnLyeCs0gyz5pZCVPTOBX7c7uQZOov3rllA6fGv5N0zln/P
51VXFpWLhKcgZrIlFDS3H0mcbKVhTSKawveDYrafZopZLtKHVkIrrm+dZUutTbWE
5PYJdXNB9sfX3m3TitcV4T5UKSo5TXpJ8wLzuFIWDCgR47SShnMFTxxSkGMjjhQU
cDGuPE4mqBEDUdPKA+1X2zmBr62yQVm7gTSAv0RCt7uQbl0tDsz7hVUXSUyKJL0r
RVjY/q5cxS6skAUEBShUR7XxMQEIDsgT05k5x4jbOed9dAUZvHJfgOy9b3CbbI6U
CaEpxttqTPql5t0ekgRekAn7q5GoMhK4jtcee25jeTY1Tp+RvYHBIR9Jd/N5g3WE
QsoZyX2jrtPxvAonMce1O0jNNl5E7/6s8/ZoyIgVToRsa+PjOGwQzkjiyx5tabnv
FhYDfDBM0+/3jLnuLBlFqhgmyHXCFuKMswB6oc4ZSaxVUl+7Rr8PtV3of/7ZOVSI
UEftg30tsCy+CYGdUv1ePb6yB/phfGv+UN3waHUUz4LVr9BPf9HqHoyEi8eUB3jA
ZkTkQIPlQrxL/17QUkOONToueeoTrEDyrstPtEkxQSmSHkp5Xdw+XdkT9TvbKdWR
0IzH0OrQ31F10Vb2FAnlG2dMq8F+CUFzpvvZxUKnevmwSV5JCga0GU+8WiY23tvo
kxLQvLwD5IOQqQIo7BMS7Jas4jS4h0fiI3BfVx1MAgRrixSEfHHAGgyn642H58OU
MVRNiPbnpPX8/ZQAmlY+kJnyCnQNxt3Kxh8JMAABcU/CCgZtJ5rWRcx7WPAfxl2f
r6L/fn9Px38b58ACDkoTePKPK9f63I84NMsULY1faW6Pb1j/eUG3ScGOe27ratkQ
oyW43uIgoWjDAT8r23PWzPFpnzjMua0vwAD1886dx7laz0bWzf03zkfnYtGqFMGb
SryrUkQf7Xl5sCsxvKJNYB9reBm63H+jxM9IinPOdyUwM72ieDObzgABHorjwLFk
MmMMukQz+GRgDUn8rn4pVgTEYeJBT43LySh+8URWLySuZx8Ohkq52fj+M3GfE19/
w88otn5OnlV0BX5P2bUlcS1hPjPLssejuRGI4tVS1qRb1fe+6Oz9Qc0jXAEE9kop
LAZ1ZNoqOwFM/CsEsGRX/xwV6hxKJACvMgONdc0DuM4yyqj0FMGwt8eIjPMs9s3a
4chor7MMZDw6cxfiUSBlAdXx2Esc3VQGgpf5Rar/t0SGh9pafm3UL6hC0f+l79CL
axdOcMWsZG0AbPhA39XnelKeioE4RqGT3OpdjjKNHP+JO0T2D/8mHYwuIleVu27S
9m7e8CDjYbKV33lYKU7hKVppY2RF6b4E7NzjudDmBeyHVH1zC807CvdTFam4PwPZ
qr+J4Oc9Bf+ITT75wAPuE4U7Xyp/ph3l65s4cAZsmbcSETZRqbCev89Yebwke+R/
9zPhuNSYE7BifwBSyVHE4bEbinlcP4fSXXaEpdQXDZ3/dmZ+mr7wonGDQmSyTgTT
23Td1YGV8vrdInoJIN262cSXQibvFU0S+CRZi/2+bixfSMfqj9zolh2ys0GSiwsL
lbQdU+FgigDApV5aycvDgm0vinPE6xWZ1uVrQi91mUN1ZT53JXcA0rKXgitTa9og
C3pw7QRAloaQhIZz7XQMl24+pyy5Kvb4so+o+kSqg3ieZXeBQbsuVX//Z1xaWMJT
2m0gEzBdOXQn7S5K/I8DE3wOJqZYVNNgBLhTQwc0PMnMb7Oo/ND/N6xPp6Uxa7KD
gbru3SCrWJ5KAlfOm13aXI1DlSHp8K/B4gmPjisIy1b8mVughSSSvufDpoIZxDv3
gLkk0U35316O3AFCnx+3hTRDrHk5NLXHNGD2CoCWhQIZ6cGxCAhr43w7D1KyfVJ2
auwOaGmWgVXFSYeyVbGn/3S5pvc57+yBzPB0RXZsTHLDAlZ6YaFf1a048lgXyV08
CWuY/jStjDngWXtBRPGxZtygNl0pdnrURvxWmDzvyly948AF1UteCbvhnbn9Dfon
YoBpYNCmuP9PVEb6bC24dKu9Wdh2pJNJY8u04iJ4PHj7qbVysCkBlfF1nr3dkT7G
skzqEr7WF6kPa7sk9rh0/NrdhiYzKGB2hHPQf2G/WfZGdwzaXvh2ydbGWRIk6K/g
LCf7lFZ6Tto2j7LvJuzxxJoY8W7wJFcbskytHyIPSBEm1xji6MhtKU4I0IvaTcM3
TtT7GCOdR5PzXh7coSsAtSQH6HHOyGeARljHq8wNxY21Qk2Q7wkjv94eQMSB9md+
SkGDCrGLDGMyY3XXY4V4CnshhaWIBQ9uv2PFLBdOWK69c6htnceynuF7g7WSt/2q
onAK6wE4vhHwE2X8yeotrkkS+0N4DWscuvqxwezTuYyw1JOh17NvOQ2gJOIpMneJ
iALESpMRBzK/M/KAeAWiCwD3L7Cv1DmUNJ49sGIom+P2WAw5bNQ/RjSeIezP80im
qjMne6pgmxyYWF8z4GwoyVmpBXa2lfPDbwF0pWmAw5iPs2dInsN6fvrTl44/3uWE
xOToKjMjQDYC+A0HK35iorHbHgB9ZHx8Ozyxb2d+rkensestmaGtqAfTz5KWjmgp
xTGbM5VnS2n57qbUWCdLNx8LspX2SW4WdMpHujBBjjEkSM1flQL5EloB3wpcFHmi
bW58psztFTaRtlyOHe8NvAGzAnGhOr3K9AO+lb2N100tTyGYt3S8h5aDpypfTzMQ
E6NhnaSPCflGApnXAufCb23yAH4z0MGwOmIm77cPXDcn4YK7F4QBwjz5xRsva9Zf
+Cha0hDIjz9YuPP+XmyvG/WB3J8lkHcTy3OhDeB2lWy393rDKq1rVDpDnwG62dbS
rPXbFj2WkroAFStHxzmSNtSDyvWNlTdDC+98Vj3Lhvq9ZyfDrKwaQ2fOjREJFodq
M+L3GAKratt2zWneKoo5MMcK1FjHUBrfjmQpjX9LA1ktT1zb19rQTGzpUkP3INtq
rqIccSR+l3+DlEEICKgaeb+3kMjzE9g7X5r9KIVNryn+zAn/M9gusq+lGdaVJg6e
U4v1p6B90qjKvbYfMxvluA35mI5MKCB1RFzzm0JJd1zSSiSFbC8Jgu3zap3IGSEd
QI2evEVqH34/0z2M2mQKMoARjq6X6hpoErUyfSHqbKRbPmZ5LNVxVGJkp1Ors9X0
CEYnKSp2wbTnUYXSv5ydvg16vijdl5/G1FXf+IQnqhyHPHyrPJEvGFdzYmR6+Ayj
bSH3UPdRYfg31Da5yWxGa8aVueuHZKblxrLqzZf63BFaQsedjlLMKIjCRgk04Jcy
ADILTMslK6tQoEOGHiy9utm8r6yRmie0M6F3TACi+hRhWm5/6WdBepLYPfOBmw2L
A5a8iwwGCiyd5J7yQzxcWSIKFmHpTkPOMAllbFO/GFsUJBQXC1DwU8r1KHTjkNSG
ArQ5Ewh4p2GL5c36P65nRfeXVlifHdXQSt+bVb8hFI/8wvN58zuT9S1me3g2EF38
UVima5wc1vd2o00hn00kC7vAjdH7cnWP9xTLLZTJ2ydYH3A+XTba4ZN6MCxio/sK
nYvpWoJzlp5q9AV96svuEZHNIOMq0U+Ltqvh/OKo14doux0JNfCdOeVuhZMbyj0z
FQ9wUcGNzbgMjHS89yvAqYXrOArx0bhhcx1XgdW2Worl6HCpQbpst4A7hTd1ca6/
KBqbUByAPqf5M3YreMlu/qSlU1w0lyKSCF1H4QLy57tQ6k83bAw6nLUxOVBKaFD5
Z0sDAEKllzK8m+oCBDpjehSQWYE1UGkZq7IwgrzJ3ugx9FEe8Nbwb+0LWmy2fsGt
xwmQIUlcIxmZ4kArgiy7Q/+ALm4LSPzZA7ktvaQpUnN/kuoVEU0m8a00VRguMM9/
Yif4S0CJGjjecsN7/GqRFAL8Fq4bn/GWwIkga/9ICj2Ha0j8jDlp6njNEOVe9c2/
VQFSllbjOGgyqTpjYMyy40LwedMPCr3hzyEDCemqpDk3RwbHzswbw/pcpoYLIE8Y
upkUd9m5QcIC2ZsZVIFw/l1y2fWUrkfCozZ+xbX71/PYoIN2Bj8cB5gxVAXCgmq7
CsWFXIpfaP3sPREYcx2z57smpMLAmOD3Bb+SokgAsuQp0IwCRG/dhwc3R3FzYmdM
3po+SYqhmMYwJjy65cCUeXbjKs3dddoccUvpWCf5gm5ooMe0Gs7McfZmC9Ph3Mp+
HBCDJW+reCYSZgL0PkGw9pMdtSXhRtXUpmT4qsJLzSJQa0eS4Odk5qmvzl7zcDzr
9ByjSzvsYHOpv4zAvnrT/4GmoPSli3GgeSWBb0cjVD4pYJXh2SXuj1y8seWJ0MZE
MBYYj2vklnOtaKotRkBHtRqqGb8mDVN4PfulBw0dsBMIe8pFRY3B0RtfMagFNvcu
zaHCIo28SWNnEb4u6fGq2Uu2UPLyKw3inw/SEJ1j0aFCdoTKgu2dnSJGIUW3FX1Y
hlmUGP3nnTKet6FKBMm5MZRZgAvs+nipVfnEoqFfuVCg6a/jfB1bhFFdGuTy0uTt
lYqQDoBptbrScLdO1FqSbFTRn3ue0yXPyiSEDEi9+d2ZiGN7TFtVGiCMiVSao8XV
F25/VLbhvtBHdFnHLV/cixug9JyCO8f+IyQUUPqrB3ITtJAFVYjperYo25VemUy1
lfo3t88B5Nt00Gveuyl+vYD4dRcLbKIXWqWu8vBShFltmo6il0ip0WRV7Xxv3vB8
6Q/lh0uarZjtXUU7EHbk8OqR0WhNs0MoYNcrWtZjcIUKCOIH3PO5T4X/3R4lSBYW
gziPiNi4owed4ZNbgrtDbAV9wYXx+V3vaoZZW6KSefXSPO5uYGt3K/nPP8AeTTR2
AcqLViueVM4DwjGxbc0XyVxWiwHdkBVFQ34wK+n66X6u7sNleAU8+llLczzpWEqg
tFOg4GMLa9nElZNzG5HuUw8bNLaPaQYJeIF2fgtuUcosZhaDYPpBzYZuMnqi68h4
UXHiZt7UMi4auTRytH/k9qyR0JIGVtCkw95/pJz5SoSfFv+ghIoeRbsfU0aaYqY6
tPhYWBpLf/0fmQmFljU5oZJkf4UruBmYSoEr3crumkiiqUEAnCgjPR/BVCnzofTU
AYm8x5AhITpKrbUknnyfmw8zJLgW/9CYOzJ69CQ1l4ya3PYSXUE9NONgD74tzQMe
bhNpwJLlh29nUZf3jHtdwnjn97LH3J/JbZfS6DqjoIuUrWiEYnmlIizxFGZ0tkpr
Me2XN+cfZ1qHIcbM7tmzkE/gOt66jrhUJWX585VJSAo9JVWl4XGZ+GwKWpdDml2f
CoT2FqV/R3IsEqK1B/lXsVTCoAvLFbvVa0u8axgtfgiVE436ZlkGMJmPt0HQx8Yi
R1PCAbVByhiUboKVt3INodmx8kdDmEhUy+24eRnwuAfoT0vQEcUpABbpNQz6/n8M
fk3QP5BsSSsPMFu/Kg4tZOS7Of54BYxgVSoIlpgpU2tgSoEPcinawi0Rfpoheiz0
miQpjQctgLFct6bckXx2pR2UqeWAZeSWy0orqPDqHR6w46830LhaEJjPDds8dGvQ
3Yf3isI5+qjw0h7uy27t17IQclG69WHN1i3WClyEWfY3hEnFQwWOKOpjsDZcNy1L
5JOYLTA3x7/r7SYIzyQctm1BhyhlE5D50CE9O6g4FpsmgldPwuL+yKJ85bwoUWCN
+jbjfs78chntG3Ho8xcxGFggppTrg5e7KaAAQP8WTbRIt5mSkeMDqw3s0M5MjIV3
/SOigxSRQvIUGyNzBF/rzMqqhhPw7ziBBd+AP11tC+GbX9uQk9JcnqCvzQKyeHHt
Nk5TQDDgIrHWLXoxLWuNyjyAE7MvqP0Zex/qrF/qnkR57gF+JgMwpQbJJWHkrS21
RiKK2c5PAly5MitWsrZLpeG9gZ8CpXh7w+XHnOYSW5ergcGbmmyZDdgVE7VpjBrb
MNV/vzGhzkjylxj3JmBvz7XmgImMaTroZPl7a3wMZPnZqoxAEqHcPKphoL+wvkDF
2ePimj1Gb2HgWbFzeqV0a4LQ9NX0FvoS0U667aF0em++W9clx96Dk32nq3aGi2qY
v9ScPJGPRWg9FOkN7DM8u9+6+CXTEbExrPhrUbV3tZbSb8xy/6S0sXgNOxAWyvv3
YiyGvSs5rbCdsnbCu0PmkZvUO/oh3wiOpbHNQ1JyNP2qRDDstNlrr+YNvCVURfLB
bZt0lOU+S18VEe64X+1g+eLrAHuXOFLlHInVT4F12XdChwy7Tkh313tcjV3LjMnI
LCxoOv6PNRjIgGEI7ACIkQ1jHUGo8ke6bsDvkyQQbx89muyfqekcdhHiCQSGq4lp
f8ObG/v6/SLIqbsP46pTMtCVsge+aSkFJNQtEsdrqY5uRgEC3779Tp9VspRVMHLt
iMXw+zelSw4UQw3ESul0TEV1dezHuKSx79/RCeHif3Cnh5CcdFUNbByMPGuWkFU9
xGmwaXYCvLhgwsJyeDx898Q2LjVW1mtIez7OMxA7qMM4WwFcrwrQWhuKavC/WItO
2xWxi3bNGnCSRVW8LOkLRtXC1jEy10IYjhi6shWV45OfWthwmN0yoA5MYAUhNsIP
jM/NvZ83+OMR417XWJgTGmRganSD2z31nwjADeRQqKQ8WGFG+ZoYXzeoz2G6D7BO
lOQIixZZsd0whJ7kwhWKqMHZ4LQs0plEghVF5kCATqFFbfVoLH0EiKdDCw/rG96L
lXda2BLrwznsCTU50Nv2z3WfdysbGtsE/tRcCa9G3j5LvxtLGi2crk2WpmrGksOU
zD7fTb6gZaRnyuu4yZlDPMMo4u0Lxx7q8CYY7Q1qV73YjU6N2L0fZSFb0Oi+2bYC
6VSjqroe+RugT1E5mpf02cVkegVhsgd+cig7UPUdY2YSUSTYmlZZR8G/tX39ApVS
1QVS80LFVAJeDXvi1HlMyV2IMnHh6KYqcUWQZi8xCuivNwApYuhzYeRZJsHnXM1i
6xuLqquHjeBrDBJKNOyoZL/HTGn1+boUO1zi2DO+30pehveLb9msthBQn7MU5Vgw
qnHZ5o/CkNab6B08eNAwKkF2KOy3R8L9bVWELYWVeF89sooWuZD6qlAkz8bgzNbo
nc47FxbC1tFBz8vmlN0gcOgFgKWNatJScgtWSViVyaNYLDBfyCrGDlvW714xWWTT
UcZMA8ZdiEGV9Vany8Xbx/jUh1e6I/kkuiAxZ9SuUcptgCzCNeOrYMO/x+LeHO6a
SkIQUMgDwAzK2xWX8OOlFMozsK4UzWvpVnHVKHX6nOw2dtSGVd4RUY7ixJOMYKtN
BVRIArqHW56iCA4xh38tEyZErtE5HnQj5uPSjjSuZK9b6eg8ihPb9yBxYimKbY1y
1DIhGBWX02deyyxr7UF2JP2WVCDnqLsd9FGj1RgeDcJTQjiVwMhXPezeuI5Wq5sH
MM9UoIqJg6cslSF6XvbqujAOjWPhWIgOGFQ7ZIuAHJ/I3kq5o1H4VNNvEDZf+L8n
G7k90+9DV21azLsMGWuK1yp2oQGmYfwSUgTKY1r9TM4+Pm4OWKiVmnxkI5A3nNtd
hDW0nukse3dU1y228xOgojOwS7s+3mGW6Pv7DWJCa5sKfbT5OsIilWEpUV28/va+
awER2Sep3YTUYYT/fTLq9CsPsG5ZGhci1sQNloo9/sRcJhziyVjqEssgYsQlZBBL
ZfWUBLnuMV9m2lAAR2CeOzzpAdLiGJ/GqWY2PGJyh0OUX4amOnyha3Kgv10iTrp5
mlOCl5X1mjR/3SeYltsz6Lh9Z9tZ3Ox/2Q0LMHdC1ltxCT287TqWZhhVoGrwO11x
GZ096K5fqLxSsSmYiJqiNs6dMki03H6eKCo5j5C9cCMzlNgmpd1c/jjxqkkyr51O
vYp5uq/SLcpp+2ztRB8riZdbl2EL3sLv1U3NdcVff8uSbkRkRnYt+XeI2Hz1x2U2
NYJk5RhMfpvXc3rGAe+jyf2wwsj4e2J0y7thYOpmSuc3Dnl5+XFXkA5lPXzUPXxd
nuPuAk25phrT7dSG5uSdypQ23tHFhxvNgcQpieWY9R0anieA71ELa+3Qcv+BgNdL
ZB2GR8i5rz+EOvjU1YCUlo/pw/e4uqpTRbjy9LUpKkmrP0ytD4lxA28SlAzXuI0Z
5ez0ilIBuQQylf8oL6N2IhoXDoWhFc6OFnEYpDVY/pR6Hibx0yMRqoSxIA7XOkOR
zDhdaOfMM3S/RjfqZM9UfY395b3oopDeu5WuvPIR6tEmLZsuFNnQ2rQ7A8b1ZBE1
F+E/4W9bNtV1WVpxBn83to9D3PDGo9/Z/AcbPgSej/HEJaVowX7r18aWiyzyg9nm
v6o4SVn1jfGdM65UOzKzp9U4dT0FexVwpOCGd5geArLLqRcHNHZuTPzTaY44HJkZ
gdkTf7h0bs2ev3zfkp/dtqgIKM6HKSGFjC96uWap1jf92p3WHsEUN6ACuretCWBs
HZcRtNRtFThpckiCR4xf2mKNOodBDHIUE8YF90F5PqtMd6DXvhCn9Ik9yrLgXlqo
7PTw6i/CwNhH8Dq4IjnY5vxA/EuaTfC8/h8MC+QYTbN5Pj7ZnIAkbsHd2svDdCQg
uQwdW4iKM9Wt0stoseXri/Ur9SDIYRRCx0qdMz31sGCWV8ZnACXFYvFqEc52QVeM
+ga59IevO3LGRGY6HR+CL/BxWZnPBqprFPb5qx6CUKuUjS0ofkO2YQ3qEed/6juj
HtLYuYMPUuJF25mXCU/V6RtVTuEnh0vMVgrIExPUzHhy+jrFsAN6kDqR9lRzKqKj
n36pWYqnBKX7FsyY595KMTmQ2hl+q98+xg9cDsWIM4muucFnJwWq7e2gA4a1KBVo
WVkZHCATlHaqVjYX4Z/wSAla0mu7B8iQFMhIj4Q2FjceYVQJUUokJwh428iSuron
GkJNhIndMjS997jMlm9T5q9c6vVpxFfgx0rCRZTIzAnlZOVl3B/jZLJPph6KW0zP
7u+AmM7iA43FoteM6W4GM7Q9+juP1WWeAcsMFckWK8ZJEsZV5Ri2Ggm7aN3ZcXGY
vVESE/4RFvqfhHROVo5qdVhTrcSYHSjOy8y7gyYPAtMvGJbzWj8y8z21IhVH1zRD
+Fa9pqjiOWFN6hp436shVgqZSHdxGq/Opi6VpZ76vzzpGI+/jGrO67vWUbrz9idk
g++/5qdB+X+NO/Q6D8MsMw46RtEaSCQ3eY6CJC1o85UBFNxW7ttwG9awuEByMk7q
/rdmBoAnuWURIXuHu2KBCbRu8Q92O7FpDPy3T9W0lqQSTxiNOjq9jQU0YOtm4O3z
cCuI41EMiAL/Y/UBvo/mPA0BIDXS0cLvvaY72vCm/JTzGsOZDjgN06GBH4iDwUYB
V3k4Ad8xt3F/919Ve7q7kY87Nk+iJJGQbuClPhcn9RzPmQAIFWgxrI18ybKQrlif
EISrl++wxv4YDikTKgJKNjSX59VBk2XKFJeZGWoEuTA9b6wWc+kLcPYu2RZsGo2R
FpwaJAILvbKnrxnCmq53d04mYjLQ2L76FwBWOAG8bOcnYx9RTj96N5x2Xxb4Q/BD
awwxJy8tIr3u021ZldDnTrkUJ3YBTZwPL7tzUOSq//wXo8La/L+1/J08lC2Xqgr5
1JyjxW5CD8tUbavSPJfng/g9kmM+evPiGMww0nv5ZdF6wEdZPsoW1ol8kXPv0oWf
9iqtRf3eDMkJrwXurX/2Vfx4IHIf2dBcivHVRN15llTmmUU0xcGA1MlJJMvqLqW4
SNCFpMsEUWrExy6kb3ilFAb35r9mcIDrvkDI5Kf+Uwh2hCfxMgcTyrwoOKtn9xFd
+mrlSegdjcj28D2NNhuAz+ahBK4HNsP7vNK/OPxWqKZn9tLgjyOC4GSaGHn2H8nM
TJ6LiUmYHsdYzRWUFNGideNNIPuCWMN0N6tbnEXYGIa6c8FKbAxwCITi52Q3KI8o
DuOYNN/zk39EYsSTuWVIlegbCUJ6eU9Vxli3lv9RyvriXPN1Lue94r5hbfC+jfbx
K2zYtZe7R49gQArhDNcf+Fk+291bQ746apeIMxN/uNaTkaPkC3JiQVHHXDxxF57P
S0iX0A0/SDtUcO5hpTdetwGbzuf0tr+prjrNHLOh+bGzt1BErpknJY/uHcIKEOjT
y3fhb4Hu8nnlfsHAvNz+gJvEb20XRox6LndxidWlawIVqkGdbyD8dnW24I9aMxYP
bHCrRRweb3YuVZEtyVim+r2i+XjkyMR8GrivBBV3VS9RPdi2DExU4+cUkK9Y+dX1
OjXOre8NXZ+KuXq69eOtffXlj62Ig5bNw+e8RglD0WTqKjDT/T7twZ5/slsdn3sW
tRWxhLdejble48r3oeZjgp3mvT+7GXw/QCCOROQzjQMvEC5BXDj1JsYtCJA6tK0x
2BoyaysfWQ3VKnUr+lQ9hbdh7yYXuBjhXIUNxlk6r8AlSB/OoMty6bz+Ksd3Mo0c
UCllQZI2tmufersz5/mNqijd4tlUDx4qWCnYE78WFvuvzCs742WelxXPH3yyhLqf
/ZBz+tv8riUPMcn0vkP60gCVvZ6DmSCQ8qABpg8KbGiHUivAMaxkmUrxy/bY9bg0
ukbP5YqPtOdwqr8LFygBdk37v++UVYjozSAHMxPQ76HFO2ndkK9LdHUMdBzB2/rB
xxtkhvSCiw8ZaskUmAl9TperTBC85EUFf/yuqgE30Ee5iSVGwm6FIqe9hjTi7rDm
vok4kYiT5xVk4e7puqOY9emt8t7bcwrWv2HJ1uDZXtVEjF5+Y4Y33NCkg/GMdCLA
jg83DDyURr+XmlEv4O4NAaNoXzbI7vq3qq+Gtjy8NN612C5vkBfbBbfRxSTY7tR2
m8YqAjTNjoMLsS1bdnDQilT2QlhCRrNgF60LrbHC8WrWYDPVKt39eadty8znii3H
JoDbSnh2Y6DIxmO8XOSzq/0jj+BrkzUWNf1yaDHGbLndigumRo/63OUZ4thg203t
iYeHUZsklYFLaQBxL/Ga64ZX7ko97z/uhb7TJM4Kbro4EgrX1YRPopt60lKpisCN
h2ilJro09k8yeHSS2hWSSdhlcfHgKTgbmDcaHfTNNdQDU8h49RlzZBaHNMGo8izO
Xgk1A43o14zXiBQeH7GpnnovmKj9IjR7CyMsaZ9Jk9b6cb+mhcuty6EKqnX1SI/q
nV5gq6f+X4jXApFgzWwFybWBa1Zd+4j6xtqfR0OyhPomds9HlzBe8Ldb9WQvaoZR
blFvPyAO+0o96/rKAjfuQTau35dqmi3r/vQg9Hn4VjEuh2kzIN+WHQyO7VSfILPi
5+o23LBZcz3QHdCRFjV1BEVI6Fd8Cm2ygwJdRGYYO7e2YNB5BUxOX77UjO7hkMYD
vK2gxS3EWHBVQ5+b1PkRyW1MfVKM7n9rr5P0VbulrmMJA6O9wctPBM0jeybIuq9v
IwA0Er5CB+8lD8lhqY24fMPIy6SDNO4mP8qHI4b//FVywIPlQpj5oV9qQ9kOzGvC
eiV+GzTFbB9oHVCU65US5/YQpfjImFTs6NUuX9aJGBhw1AezX+zxo9H0EpahuJoI
5+hzlPjh/dkYa91eKzhyQpb8T95GLYe1UAiLPbAiErx7cB9qfMSpxw4hC2inY1Pr
94UR8EAJeYmC2SHZqt10LnN+xc0BT7dGZvWmxpoo0pLkjuYRwpU0kCr1Vhjk3iGX
qinVyK5EYOZDFFbWabk1e/fsTHMdEhupDX9GopiSEwpuJO28BXPNzgnZWLEQXdJR
94p+f8mwY0Ljl/ucsuFctNllG/GEYHHRIz4DdNntBYVf6n/1KLyucUooBQi1d995
oIHmvHon1TAA2BmP0/dRFCHv+34ILs+nYNxk94ZY8qwkHAJ+KKB/X0VJNvGRUB7k
FKDeO8oWnZpslOx/HFAbL1EMBX9NwE9lFr4Ga+xIvnM+mjY75XBUZpNpIaKyCSFw
Q6umBKjhAKRnOfSdpc6MldixdjfC5WsWYwCqz2sDlua7HXOUaxpDVt17BsBisJk2
E0+DV1FUGAjX/Fc1Vhr05Q0t+ZhhbFXAIISTgPsU6/BnlQfQjqOgRIyR6v1RHkAN
K+ZO/sOan+nrTwWhG5HrveK8EhNkShtsL4tt2z82fuQC/KNIDMAVGQ/7WcHZORXP
764J2ylmvlV9JVj6osAadAnxUm8EeoxhP84l/As1B9QCZWNdObCYewVDCZXqh6tL
ZgiH5f2TA4xNySrlG5+DtgokLxdee5627d6snt0jGORgTYOeyyJexISMkkjyUHe8
ywOt/IX38qtgb8RzlBS6HJLHE/3vV8t1xHz3z/tk0Eaq9SmjOeHZ7gxgrn5fruxG
fq5RiQXxcK7+E899HOPkK0t6rN0lHtIZX7PqCdMSgPs2oBAmmh7ez7sN2tRJhd1X
L84rb02u58In2pncUJRTiOY2+/01oMaKv3Pyznr2SAMSd6+9Z1+mSiBW7mqVS5rv
7ukbIRC4GBr0/QDEQKHOsH+x/8J7o+x+BIcqPxcgecnPRwK+BStFcTimDdMNpq5U
sFCbGu3gkK9TVckAxj0kHkCFe8t9S44gEhhMErN0NOI6zX4l4bb1IVhrVBl6Q87c
WJbm+eGPdC5yGl6BJsJOsbB7jzVXJ6+5cNKVUip8OCEv6xwmFnzOwRaFuEN9aelq
9XQ01iEGHKHDSFpnImB9Cb8yv6waDs8GCQ7vTKt7F+nx8FeL3/07abd4vHxMhWQM
BE0fqeKXJnxNrvz8+m63JPk0jSytY+MWzZxv46E2EDgfuo6r/4T6sPf4Zrfu68i9
WI5ccsGfNFXqPnXLZNkwWml45sz4iAc4jcfJjNnMToOcqouRbQr00qqEXF4t0Dkc
/slkYIy57Nu8kAVnt4EWxYhIVA7bXAD5J/geTjnIXq3D671ATbT3jaY2KbUQDklz
g6sOQiTSdKjjNKtlGlDHD2uf7IaMqIR737teTt93wOyu1eXvRluNUEDkUu/LcbXw
jG9l/Lvb9Pon41nsVh2rlCYqx/r/RIPUhnIu1zuD4CtDZ+wQzoAwX5gI4WHPtY8H
z7Fo0lSm8F86dmDwOtOhs8/I+PCJT7WEzuUDFpF6gqGKHweMMGhA1EUo5Cg0JVpI
+dZYLiPl+Eb/wGmR2VUrAoSs+GcTJYtVVKcqUEe66nF/GJ+Hku0JqlHTCUr9pMtr
LETU28Xch7sK3Zzp+RNUWVtTiX3bUnfE8ojwez4LIRQvVlQTCcMqrwCZreB0N9lg
HnIFCA/7tRIeeHcZ7FY6CRts3P9rPh3BGdR78SehcYrP1X8pdr9AB5kt+YFJEsaV
WGpPMkjQmePMBG4y7/5lek9cN1a4hzrLdxj3+5McZKUzg7Y9+jFF5avm8TBQUHA9
TZkFu8roYX3NchkxG+Z20X7t3nmqIza+fj+8mH3OyNZbCGjtyk2jMTOoDOyfDTj/
MVuE8n1VWGu5fUk9rAEhP/IYLFoZSUvIbPRy5Ps7m/fj0oBGpsnXCynHPyFmNe2z
NduzyUOM0i027EFoAtTayW/1T/OzBXeLkFpUjaU97vtwIGvyxVuixumI2odgvS1x
/qyefBTkq/guMKHJj6dqfoJpv/WV57k42dtyssdkBJ1fVCU2p+ftTGrZzlJ5Csdz
PTCi7NHC9pcEAPcDjqP6xuaXWRUSvQpPAx9Kz7/y+9j68YOe8jZ6AFkzIwr6LGrJ
Ul9OlS3gmncF+bu8hgy+liznPNcjDbt0yTT96Ao8oLgjz3HQMNrj3OUoQH7Utfo+
4bu0XFo5sF8E4ZXbVXLduFXvjnPnaFkiL6ovyQXlMir6dzlNwgSX2b+5lSKihc+Y
t7sTe76kyXhaTr+UKAMtP5nVLREFD45ffFbIf6bOI0PGxN50E+9jetGtUqr2dNik
F3hu18n8lezt01I/0G4OiSsAlV9XiPy9nYCHaKUeyrxkuu/T+DzjNp9qdaH2mvFZ
rKnvS7rFUIgdbfBvcoYClVo3mezEDocZRLW8RFPN65BMdLgzvgd54EUYYcggOHy1
36scwnviE5Qfa3bG3ppSKCj9ggT/HKXRyiZ5xEZgO3kI90XBZDAqkGAOAHI5wnw/
sQRuO7T1B9xJf8xxgz3aFMGmyFq4nYSUFJHo6yYiVpXg7CmdafinppSTJNcyMHh6
ExMBmnEzqM1HF+TYGAEOJemudUXW+NLJnHz+lKcVnzp1jZJQaoYH3H1R3uoDFB4L
9Ef4KW7C+Q7Hs7j6QjbWlI5JS0+8Xepg3h+KPZ1w0529gfA2kKSRAEonaVO2lDWq
DdijVX9gToiKEMvhtHb5wrY9eF+GGbNXUGZJta0i+qMXbJlRKFGOC2dsFnl/DOsA
kKyB7n1V6cE0IjO56sZRrtz9Dlroq3NuQ9nKW1rhwBhHWi6n54MXbgegIKV7/OPs
PJFkPGwAaH1y66GhtKdRVInLdPIWLHIc5LhzCC0jH2/CSGXgs04rQg8mXPdkf/22
Gkefjv7hYL20vdNFqdLhW88I6ghcP4QnEOMyAVJnaGnGCV8Tvj+lz14th6NEZ6Pn
0sbTPzw4bGHIpXbpbDOJrIBCE/sodoA2LUcjcOKlDsmVz8kPybcRqHLXmTPwSwK7
PNxfHO7t1APeOj6ZEUrgvKfeB3qF0zkfFdCRpHk+uhG/uQUfkXU3YvJ0DpM25Ty5
l4XhpAWhF4IHLM3R246bxNZWoFoPBcNInbA86K1ekT31rQUWpo5af1GKe43swDfc
AUhoo3scscxe52jLFQ0UOrtrUHG4VMbpVpKj+PBTk8BKbXzSOW1ghsgyjNlgOekR
pMK8ZDvbFu41nFNdgnOyoPTZis3twmwc8ukN+usM6qvNdtg9kkyl7+YOfOa3D4Q7
Nlm1n1+3Hn5ZrhRMOI3uJ5V3h6DGxXCi4R/Jhi1cVK4i4w0HB2qVYZztrefho77C
VVQpmOqELIJhISzWnyRRyQr6VCYIvqt7KP8Uiz2dKQ85bZDm9g1WMLq6pQhjXxse
1YtUnRcjfqPM8XikeikoPNsBFsFCcLREWLqWS9smlJwM1qbqFRkz76TfUDCHPnYT
tD4S4JEuhL1MHzDDgGTiCmo8pmtdUfeZNT8mnmo50q5jpRT0Y/sPZscvQIt/hFr2
Qh5hZudWgrK3j16+rjyaNvPab06YP4BlIPqmEs3qm/iDgdrmq3npZaY9KOn6y7AR
MgoWLWQd09FsN8cDRc4kxc/QbFTILPl441IUQHJM3kicxss5/LisjOvXDgyEjXPS
BSgT/AuNY4xEVKSb+jN51kvS1owo8bXNiTgwDsE3qK2/gPpI7KX1mm26Wov6t+Q1
rWKmeKyUmM5pS7FqMXaZFgUxNas1F4CKwkUbbMi6Aer6/p2sqrcDnhtZd5Qh+g3S
ZKiHozdJvoJcxqs0Wl8/uTq2XBRa2eN+IB7IVADlPBcYVSpZfze+zS6BElxd8WXX
6ffqHYYslhWb0JYenOuIQTB815sWoGYV5O9nAi1mG85DydiUTOD/ZnRFQSeBLE34
gBPInn37HyHAJOEgwq06HRB9StxeuqB7wD8F1Xtq86aaIzKgpqiVK4h7wm5fUb91
swRhy8uvUKN91VLS9uixosxL8Zre6DpIG833EXPyVztRKhgBikKHTYBAW3zPCZr3
/lmuGzcHNBwtIBaZAPJG6L7Jqf7gfRkwnyJuIsRGfIrayR+a3080fTCkP6azP6Mo
zbV8Kb3nDfguV8KIyOA43+A8SVXwH5mYujKohIJcoQHgOwKFHwwHSfGrI6kN2KUs
zIl4UpppD/IhHAS/iREtlcIaSZjh1t61wBm9DzK7oXYnm243oBpLxRcUhDoVsXdr
njfELM9BNQkLTFiuk5aEfncH4GfmeEmE6jaDxoPuMqye+eIsDMWGpeWkk9ry/wlJ
n3hXIV4krcUelBMVkUGWvkocMMNi8fESqrQHBkYrF8WE33dfTpd257UgKYRDXO2z
2KeZusJv73yTaRf0To0M1IDFdzfnN/iQeCvALAET/lzOVFTcWoLsMMads+WyHu5U
nq5G7ZT7aNb0KusDOomm0/bxgcLHDpfUITly9RMq16v6aKpJr3s7UHRya8Ri2qjp
/7ZPhlsuVvKdYfeAULwStNbgWXNvlytVQxEhiRCw1AS1DBOkGX9ew/I71W9b6loi
qX24f4wej8UhjQ6iH+9nT6p/UbwHsYuOuYNqa0ffW+UTmr3MXF6sErZ3Zk+FgiGp
1KFBxmghaMIPHIgTBVg03FwuXOcbtrrLJw6/sK/3hnMQbyqlWPc28+4LLfiFmmTk
bA0+SVlHEL1V3gvZ4o8FlZOwbXTU3RrqoR5HhSnVq+fjKW1eBKnG25eYSJ5FCtGP
dwVh7xjWxSmfkIC2gKAnAQ1ToLIWDoj++AEKDnx3ZV+3FAu3LPsOOZ5qGijpyGnC
QOeiOmw9lE6rHH9gvqkIcq2YibBAQ0L1qTgHp1gNKojbPV1kYuS+LZaKy6lcuNc1
aDpIx/nprAq+02P10hgfUkdF4EOXwwjG30TwjvX2iGVjIW+y2DYDQ8eZEueXiP6L
jjUidxxcD5kX49dKu7/luOWd++MGneFwGg9cRty09Ibt0yeVYRcSRVlDOi16s+X7
ICrWgRXKS4AxqlSKYZeKAlaWnlGoy/HRZDqjT3ov7X61OskmlRyRGigM5/bH1lde
fdsKJ2ol3LTCgDUfQv4VjKKFp8dFAAqAn/HKXvz5Fmza1B8ccHwg4SiasdeQ/Q/L
kH/ciWBIKM9NUEbRM2xX9HixRtbtGkGYi4TbFebv9T5Hr4oxQR6UgFw1dKjNtRPH
f13mZ/HzUeiQCHIZnXcEROlXLDQkJer5Uf8MzTl1X3OZXWGmjZ+wPj2qwB7IEXZA
FizojL3I9ngNpErgBgP7H9WXYt0XPIzuwCx4YcrBbVrU69ZKhFhoMvQad9ykFGEZ
DYCUg8mvEJDDVOh3970N5TVBZDYZffYqRaAO1ZldFsxcO2RHrDJKhFfyp+D9k0iW
4Tl37F5aQKP3eYh8g0cq8dCHN8CSkswW9LoToNIhn12ClpGQxU0qjMHsJflor6ej
wQs0W0pTompOEnrv+344tPf1514YKxPToIXVrd9yFHERHkhqzM2c6J0bJrk7mx/U
i632sQ2p+q60qoe6c3z6NVAdHeKvL01Zq3iZvhUZjXvyV+S3XRjboGeCQZ5Qx9mu
EAoPaKA6MhN83diCn1sflm82y2S8QWzr0b9adVCCNW/aQs6iezE+2w3H6obmSe56
5afYVJXAaR/2kfiW6KWXS2CQZEGDqiYU4lt2gOXsD2zmxUl/AJnCUbsMw3BE9peI
shk/dSE/OlNYeUAWkk1ag6lc6rZXQHbayJ0D/ZG5hgDAahlxWSaOn7SEeAXTHI0S
YBRh3aNB8y5lmWYvmlSc0Te9Z7c1zK+bs6Fcnw/H0KhXxB+VJGvh/SkuGEkImzab
daiyI2MKZMxnf818PbGuYviqj9I0nVrxJgYCm1XwNwgpW6Kh37BshNA5FQKHBhS8
k0mlJX1Acq+nJ5Ka22rJ7VEQ6ygsooP99xdWXym//vb4Wxzq89Rr6O6LK/YrHn7W
BTbQKI6cKMNUY1SkWmi7Coow7VB8qU3Uxv1PgVvzz+NDEg5zu67V0knxUns63m7N
MISnqIChMzbYfRhIVSgJdvah3LoKuEOpEo89zzPtqo/8vbGg2cFKH3A8x3nxtBAp
wVqM8xD93uz8Z+mpnCTVkl3uY0xHJ3p2aYnFLRnepYlTc7E1xa33hFhi8tT/JCYY
7PHwh8fxfLaY8HWeMk/0YPTstte3J/8WE7wm2jPSlk1irc4zuNdpwKvNhDitRmju
9iM1x08fxIxiJ//CvJG3RVwPcHm3P9sr2JspTBzu3RFbxzQBQ7xe6zOXaNIu/38Q
vxpK2uJswcGz7CaI9LyDwNuM2p5tj46LrjR9I0PzLNxnzbdtZZKPOv8nCW7n3WMB
T7Jd4w0TOeIkD3hOLaxVQKugnnvnmFJEPcN0BRQNehmt87ffRx23B9AEVTP19Ssz
3EX26Zt3T7AqsP4dvXlmid+8GdaqGJSyH9CAkmGkG5lcCh9oZiXN+3ziMQG5dl6E
0UTUnN89uSj0/7mSqKtenRPPZSkR4fF9eQDWKqVI7K1RrVvCO7i+P/MySMMIMD4X
/a/31ZnYek/gi7E7VFhtFiTpnbFiDMSrDoYEIhF1Z6+yQnp3KzbreC7vLZLdxBTf
MEcYn4+8nU0HZY45o+yJPRdQBypdLCK8+XER0jNNvNct2r8tLMyu0YU5xROpQGBn
4gAAoq8wYiMmpRPneyLMPLLgrlsfFpqNhYejijw49SilCODIo9w+UzCWjv3X26rM
sc3jkUJDmLjF4c3plFWaYp83bgT0oEwaolkbcayT2y2urjSQkJSNimeCgvvgGEuT
HbvL4Wf7Vf/Xq1XqQJrzLIQHbm6V7QqZYoRFhhyUksapH3wErEgrtgGvhlxnRG95
Wc8u5ICBWYyiMsKF9nsGSIr+ppw/+iAvVdV9HQlhQje0syEOGAQv4JIg8xoBljOs
uKvGZDOht+YLKQwU+f8XGuDFE5xj88fGpiAPhXB4o7+ErblaRqOzHHoKAvz+q4g6
C51bbkqb7YWKiUcu/ra9TBXvGxufZsuYkv+iEzAUDV6XGtsVXEPOAshvzFt/RTiH
xYDyMG0t+u02sup+P7GeqqgXwVfa9OUKJ9wlC+i6UG+s7dqhCjG6wqxfn6EKo+Sn
uOSSb1sTlI+S/Ip6HUvzr6NBJD1sjUb8aTZupT8Er3X4Co7rfpn0A70vbLrHjSTQ
k6pgAYB0LAFiZXsxKH8/45VIRCKUBtGYaa6izElZwHHumo54HX7uek8TdMp+yw14
xnH9LplZ0rKXE+O7/t2D0EK3jf+Mod4aLZ1fNZh5XDP5a9aiL+NmCgd8eYbDRglY
umUw588y03agkrvhAt2qn4/wPfBMb0ukAt33+zurqo610q+qjtBCzw5C5MlPOMDq
vmbXPH7Esx46ojexHPC4cRoluti3Ub8WyN+uD9t9b0LjdzGDPTD8RcDPTPrHEDeJ
XbHBUpTo/D0Hxu2Sz14laKjsNikkwbvv7lFRSNn4t/ojAfeWCrmBd8xlR/DSsh2A
MaMKhcnSL10hFLedT1Fr0PgSFZXZ6OHS42FeSLo9ACRDnD53ymdnvycaj7qHnnWl
grgZGn/x/E7PLClbR/Ey1KAOZyn5FwCDHkBtSDYpBGeS3ZEBIW0K6/ODCOzRpMSU
48QFbXZIrqsHHvRM4Nv6VQlcNAUzpD7fnNO4p5oH5LMzzFDslV934fjbFhJ7jrRq
hdhVcOJrrDv9RCQ50P12w6UWeX0w69fkAkLO2xqmWVwrlFqGnlFH43KdLtgy4p66
shpipGUE7xguzSVcSn3X36LmseNYAUl3N04BqtxhSHL8BmZ6ZuwsMhurYPKYhFol
BP23d+m2APmaE5f8is3N0h2zi+2O8Dp5T/BeO5MqM1bSgAl6s1U4t7fn4g7ERbVj
zr2jNYk5YMxn2YLYz1KrvOUkOh7bOvmi/HusOcf/LjRWn/bkSbMVTKpStIAxUO4q
JhgV91+5zobp0AOJ4WnM3rlkRrQIffsW3im3I4CLyTs4w/22rWK/CvCg6ASp+QTz
pzNvZMKkgWuMgvu/EoRRek9RktSTjG5nPVtwS7SuqQjYONL1ypg+zllL+MsGb6yy
R3RWLzekC4vi+6pnw6MD2XheVgnls8RqEF0zhbKFLKBLiPaeOFshCmnIhC4UZ2yz
CzfxqKo+cVqp+0+7NnCHZBF21q1vPyNGJR/CwmkTTfXW+o160+7icfJuw1Bhf/Oy
AEdRnn25yIUZZFmML/ZYQOxP2112p4WJZgAFdod+eiKlTR3bfLXnmUhNB9e7GViK
QXC+rBpd8Io3MgU7qVibrhrJ9OioD6a3Bzfr1j5RiBUcGiU+tMyiMIG97ZUtEXZP
bYoODkeibWvqNZqrzm8XrmKO1bvRQ+w0AQjdXgsh5idVtDYOGZ6d3q2iq4dzG9cf
KSfGPQwa2ZBfHhpPGhJteBQLlaTM0JW76zYlEOJTtROodRCY4dZetkkZWsrkZJTL
SdKdRv165lENARlImrFZ6g/Vc4yU245/idUzE8nnwohtelD38GrcjCwmbOBJsXWn
zTIzxPSr0hh4iuPDPmo7/Ha23w4bXzDOv1qopdsWJBYJNcq82uJzJ1joYXKo4hpu
Jb2wKdMgXAdiKCnPvVIDrxV5JsCu1AQrhBMI2Xu6gt5erEeOTDR3zqUceUIx70Iv
4+UTZ8gbjCYv69o/vFf/xKfTjX2DQYAAHa2eS8JHvk5vR6y3D2+pho6YfXxCUpwx
yiCfAoXoqfi8sL9C9xrwtOE2k+02b2XVTYI+hI76R0S7EitAezi/9x+WXe8Uiksf
QV5oiHV434U26KA5PJmKlQqZ8i2H8KQ8jiPZEvcoA4pHBjjuE4UqfQdg8ojwdVKN
WPuw565iU+LJGhv+3YigEAPUwDDxs14jT78lqEbk5y66SoiSXM2BipQgdZpyPyTa
l6cMmNaEsdG0fIMGy9M7DjVtqm7b3Lscz5ugscOKlqenbKp3XkockNu19DXc7xGf
XE5Ou4HLcmIxw/FToxtd4PnqOQxU35YNl9O6vj0dL/LQV0MEj4iqls66LPfhknN5
srwTSI4E3qjpYTA0gNMHwC9O1PessqoYeiNY4t+MD8ho3HkX+1SRIP3a7z31bFDQ
0715qiNh5zkMObz2HL7O8pjNaaTJHS3KmDoym+J1XngL7YB14A1k3vjQYR6nGSll
cHCg8vCaL8WqZFvr0sDnpWiVdNRieX73+1G4veGe9tpxiSpVa8MdfsEtXkcr1YKa
uIwbPnklUNTXCb1TqM4v00EJztrEaRwlmzWdP83AvKlNzb/nHrg/v9U9w6fVwVUI
lNkzy8IZEbqa7bLJhDvBZPd6rai6GACaVObmv4LYfkoovvlM2/oZhUjUre3qYa/e
aPunzO1em7cw8gkKabsdWknZX0JEwf6j85sgCJah9hXXjUnu9Xrh9JahXsToRCZu
gZLQ7J00b3u66uTVzdUn5SdX4A7n6TPnUfm6GcNXt7MzGHGlP9/vac+gxe7hVnDS
Z11wGvL4pBmRTi6hLVTl0nL+pVmMecnx/ao+djH90glqEAkR5P0tlCcixHZw94Qv
78fNF/HF8orf8YwowOcAEhgrj6p+MpbRsogPanO+MY3RqaNZFhSDkEnEMOK99wEb
xot59rXQFoDMvKM9zpueknChfuqEJXi52nM7oGAHjw/TBbk7MmdNZ5LJU5UH3Y4O
f+/xO04ke+1hznR6z9L6aM9GfTajcvykovuaKQXVj0xQ/Om4qI6r/0QR2myKyG4L
rxrtRGWuOj07Z9axLPLcKAiAZHlpNfy5N0b/6n9oKiqh9kNQyixmJaXKxBJ8cKFh
C9F4I5D7nmhLFghj6ZoT95tFPNjSdng+b4K9CNu8W6eBoCUJrRLktxwqCqCfU2l+
JP4GI/kEhEKmkZhme52Y2m1esaGeYooHl+DHwtWSbKwDmSVYvt25iWBFHJqk8Swt
kQrOQFPBQ9Yg3Rd/mWbvLqAZTJSqJztMrWkSbya/NG4W4r1xMyEBSOkl3P5Y6U+B
2mVKRxkkONBeSGyOVTxuAmLf+WGFQo0ba7jdzjR8NdXP0RqqXzUgooHOfU1Tu7K5
lvUJB3SR3wQohzw6/ZQIG3PRew2qf35KmQeTZUjMMRvUicYjfiOYiLp8GELnu57v
AzxRADPbAt7Yqzn1EQtupyUQ34MmteI2XJ/P5oyjXAjL3hxIazB8z0F5bd5keGbr
alGwnzpH66lWKujQqe0ekWVGMqJzLqWKqr6Br93/B4DAGbzLXOejy6fVzRPeVfok
UEd4sKrwtTo3ArzXqZYvh40ohKMF7rnewpprMb1YbmaoFsT2PEc2FnpXQp7Y/sJk
44aRNuxS/LHthqv9skpEfrQF8gcGgIvu2XunNSoiCVc17BQp3TZ357ydNU1gWq7x
xSOVrBRW3tbOjXfYiLyLxFxDkovjA6hDWX+ADKykijo6Ao2PAVyMhvdF7a+dNEJi
w7trIvagK8plzuIT0y+wpQdQuJ6S1PskKEkemu76oTzXv6BcELBxL2tZX4gDkMqf
yBnIn7vJX/Hdib30/NOvb9JwmoLN6BCB/YK2nUXKC/riEg+ECpoVvJWbmVywfRx1
lt416ab2B/ESvOdFGrMJueqVegfS3P6fr7tGTbHeAgQ5NtAMnEhG1zG13IQup1rA
hJoeqRWoLSOIIM5xj9tOYckJ5Egun69lyV9xnEbXvh3YgtYpTfnxbg+mY8mZdML0
xZ+W9jmjJHxeFGbNzUMjs/zT/j4EnVKcW00vzJRunZoicyZEI923evfdEI5NfVEG
loovaVwVmCDERX3g4ZO7fRTdNbcDh1HwWRjX4GfbGInLzgjoAZKulm8x8sUDHDdg
SPvB7kyGZK8GeWYtneCBaw3KYAdT1h2nd9EKDfBhocdKjga8p9GVqqG2vz2RikLf
E/uvWNh2rsXUOJ1+W0PkYXVUdrpDfCkmm0W9/S74s95+5R2atNWIPTrXMLWqQQut
85y+u6Gps4F7ehKGEjdVz5w0gsklRQYE4KVGXgGPm03oO+sdhcPSxs1CbqVgjtIc
wl8Nw6Oos9wRf66BMn+ksfdmdw2CZkAzIoj6g/BPKaV9zSWuR0unHbSsmHJcdnuB
6S4AgZiOBxHBSMLXwhzqTbiGI/VhaWFgmWELABcQf/YQTMr5j0Ht9Tqviqg3eJXm
j400zU+LesPkDsDu1N+HsM0Zyeh2Se3z8jCP3o0rSOTOKjLhc9qll+TYcJtPVEKm
6f9H6uzAo066gqgpz/qa3tg1piDthOiqw6NfxNkN+U2Bm+RVgWMr4DVQH4DyBQx2
+2L6CsdioSmHeykHdZyQsj5SStESRHPtS8QTuamvoJ+Dfvvyk71DotQGXlOjmTEB
ikn+BDEyt7AYUfmwO785KLiPVSNDHz9I4ZODYxlXgxRkZ2F9H8Yka4nqMmfh9wS2
2D18nkx9xlTRFK6DRF0w8trYfepEs6iapmIJw7y/zr+BY1+6BMx4MkpeQWhzlQMM
qZWojPgpPqAvUb0vkgUesAexMvfOwSh0TUxx1bz2k7AMFDp2qZA9I1f2hUqdXiP0
6jOul4F38/+RlYWC0ePtkrJZazlt2Dy1iGmcyijsET8LICKNZG73c72UjUj/175K
seSPCQyiOmD8g5FpZ/b10j8gI0SI1IMquROw1LiIZcWOkb0nptBpOoqeyegm2m49
5GuypBIeLOFLQFGdzjlZPWKUVkxrXHwj/yUpvxosxgg16UvmFlTxbkDLc3n0XMkL
M9LpngfK5d1tQhb+G48Utj49ms5RWAvOITLW6wVBsD/sLb/GCQqeduAkdTykM1dh
ow8BLwfD/+IqUGyRJQNpI699FH2L2sDJf+9dOQAExm4efawVx/nE5uiOOpaKr0VJ
h25XIgDYOlg1icsQiKQTdBCnRYFk7HSVqTuyO6KnP1thRroMCrmISAhJxI40BjIX
RAGtYnnUkNS/UsagdPhYJo9JRpb8UfdV0zpUA5TmCY1C7TjPGDTVhb6lOdiLVUdJ
Tqmzj7430m8UyCtIopoPj+M0lFv7FqRNymu5fE6Tq9qUIMpVs/+Fu/5JtY2RAJWO
fqvUBuAh5te1NHbzjW4wrJF91JfV9XAoY1BQpC0KFmxALp1rPCOULSs+k2UoczZI
fa7k4AHM6Xmp9hM/DV9vZHZ9++ky2GeXoLH4etaSvmXt4kUCbREGccntOopTFrJF
CHNuJYWxaZr5wbldh0xggDQyJBRRdry0TSiA73G5ErJxS1oClaoHHMEUu3Cqi0oe
jwGcRp9jY56g2nHkh5RZzs+pRLJVt9g+H/o2r8VSlN15MrQIgfBRdcpYx2vijKrd
d2YgC3yIFck7UpLjXluDgS6JVQaiBur7C9ljW3R2viNx2cqWYPYGPl5e/JtFPZLb
MuAlcdyzPDoum3mGE6sT3KL9eokPZzNOCEud7MymqDylTS/67XJIqkyxmIShCqm0
wx+Wz1KgUPA1Fwtkk/fflDTeWdflSuG1IfEO6i0V9PD3xUEuuhTstTwwB/QCNZtv
yj4NTDIAGRii1fQPzMyzG9Nnzn3fXSHI6N+oYDd+2EgibT1f3ZoMxNDhH1T6wcAo
7ULyE5UCLLY8RMGewWtqnxaicrZPRVfROBdWxsD3mDWkKcu/A+6u32qR7uVL/qZU
yvOk75y1oxmKFT9vjgW8VXMOKlyYmTNBhuYuRgWcqkBIZSRJe8A23xMTfn8CqnkS
bIhTOvKWz+FEpGZg/olkeBcmu9U2AmXUNrfnInF29ngbD9gw4OegyRFf52uWZiyH
Yfb3GzKUDfirvEVxI6jiJPFjPkJGRwMwwt5FULORaoU4f9Aua/+m5kWDlTz51rZt
fIdx/7VALwjn/JE09zEl5hgDjfESvZFQdaORkyVXlSCpBaVRnEttI2p0ghAb636g
nkxmAbq89joLjpjhkR56CD7a0w+++02G4liBpQyDXhzunjOYRBolOZtB3eKz8A3X
h5mZnx4GDATG1x8NRzWKBWbaIapWdmUZgDSSHbwZFzD5WWwiRBrW7AY5eC/2LmlZ
FPUzdVhVwiW9n4RjTubzDpvYaBS0+q2NryZFOYQmTvb4o2KjudQUvA+ktotv19G7
KcB12Ep8012LAolFfOViAnueuhpMdLntiwWVZ36cGaZZeZ4JzIiFgzpuQ5+g8WSm
rJZ4HLrIN5AFt7IRrJdIpck/cJ72OFRTRy08Bng/2GCF/q9+Wdq/ButxY4H2fh/s
/NZ7f2v41KycsPFls1xRXltnno87nqFj0HLurynbkm0C0N6wB8o2/EW4DlRmMBVm
RrgSNP8M14eMBPVw/uqpG5QlxRMfUU2CJ/fHG9sOG0Q7PlmrnTf9EBD6dWFRUVfI
/P+wC/HRRCg+R+6rAxXPGclnSFuESIdALRFqiCaLTnWYTHqOkPx2rvC6/T1ueyvU
rYpPaKNLvq6/oMfJCC+TF1hi7rYJMMHL0MxOoRXrsbzTR87zLQN8DfPflleaZaIh
ofTzm5QwRVmuLGHGpXaqeyAb7JluiODIUDMx+mn9EwrZAqf93i+pDfOch8VOSC1H
ZqQ35PrXJaAf/V3bu7Iho4ifBdOsjTZ97pEGCJBAcpovnHM7rYnuE/qwS4XS8bOg
FeDgLxE2de00NtahD7bkCfzX7v1C0jjVAhUz/tFAWF5Z/HQYiZEImBJr2K/Ia5JI
Eqqt3JELcT7OSfSgmzVnRrLi3m6Rp1xsSww5j9NSKCWxQAEoLOEA3CPuGOFomN3t
upkx7M/1KJSmDTUEuCbWv9eeEPHbHk7lhkQ8JDfol5CTTYhigHnj7PDpr51MiTDW
Km7ujUjFSdYmdIIOo/oDpnkR2HHTuxLOx5+O6kZVSKwOiV9EydEuounQwd/v30Kj
9wQwKbHuBtLLuVjzp6ENecLjSsQizugNNPcZpLVlBm4i7ipBlX/uFp6PkkuP9kVD
j1kSSzmj9ClSi1y6T7zrzB4Gmrgxs6BUJf5Q97FeOrLq4DjWTQoT2hNoaioHVa2r
FGW8i1u+4xlByhRF22yPQDOD1DfyTJtkBG9OdPAULivABhi1cwBXAzJxeUCEVL58
ZCCpc89/Iie/X8Y2CVBKp8LPH6iW481tJDXjP1/jshi/syK1RWI+lJ7AItl369Bf
wllfotYl1+J6M22BRbfPZvgKL47OQj7GmuK+QOhc9eLvCDU2AvcI+IOeK2mUwE4Z
9t1OGhGDM6r6mc0fPw3hCUmgdcESPnX/6zpA4F1U3+w0twt7VPUmFrOsmZVOI/hl
coCBiT0my1+gYXzsva5tpABZmXXAMlMVApfSoW2PoWdRogmda94r+X7sAhVXFkw2
mdD9fJ2wLAUmF20r3p2sJcU8wc6Mvi7uJpIanjAxV+AqhsFH/xKJwgf3B9slHLXk
LQ97GKFRNIiTdD+DJTdSOzFqZx7XUSw6PDqtxiZ3rB9u3EfMFqzb4n9FhBJNIFbV
rHn1Q8NpFxs+15z3+6gteBJ15rBOAD2n+/D4row+S95vLWKJoV14ymgXxnxVO2VT
6WXZeo4yndD86SWHA7/u2DRtZIirr9L331QAzpcKAARmLyWGdpjGh+zmmQyYE0O3
zWt/x5xXjWpouwORjQy35jLh5cWIZ/DqxJLJzpSfmigwgK0UpJYLyfsVUxO0wx3m
ClT+tHU0ZBV0Nz4FbSH5jTruaSKsbVHl/jc39IYBF30ldcr7VoEY/lz+hkx2i5Y9
tkbJUIrPumm9o3mgLgK86kINmN+Fp8YIbbIAW2i3ywbxbtnjlSTN5JreUqu7lIN8
75t00SuWMV5Q60zbPB8tBVy3smpouE/B3xnzDbol/U8yZ/qy/0OKiPXYk8T1sPpe
wBXTmaZv+cR71QTWKaedubPjO5kYNpqRY/tInOlviEWByqokV/w0QvYgi1bLEbXy
qADE6ZVveNSsD9S/ZP7+tpDxaOKJcusGaXaXNJC8lfSn/jUY5qVrHT1sXGp/oNzV
pSQdtj6bUsCsjnSW3l/AH7wQKKsFl1iVRR8PgUx/VCH49MNmcd/IDiAmXtl8Vsmq
tjvZhzeLwW1gutx0NWRRihl9dvlgWIVCBwk5NTbeF0HlmVj7NX2noIvzSR7+jecB
5esfLX78sDj1FcvaR1oEIck00AeSe4u3yItll7oB32N3ch3PxmL0EqlbQWsoHrWw
Q6fnU/C9KGutzhXpBD+T2BGybYwcIcDcIct723JYB++ZgKGx3yOtRlWO8NOKvw0c
GT/RqDp7PhTWeOHWNQ4W9eXzaU2LY1ZeAv54HnE8n900HMoywiCwmBWJpXkLYKCR
NopSXNZehSTBP7zi9xWMMyiW/VBvC0WKDQY6p7iIi+M2gJZXK5DfkJh+cZu2x86N
IT0d3qXeFBRwP4NHaPHh0N6WEKnIqm7hHewUYin1API0hbhfmvryPmYm8PiNJmcz
bzTH0SlI/NJXYLFpe7V+vqa0TEdHFSupJoqaID2nIDaTW7x0Vkhg4ggHaneFN9tI
2to9cisZaWFsTxb1ieAq4xCKUWpv3rBubuPI3oozEUj6rvNFtWQuQLgQ3gwQBVI9
EhhM3rh0KDbiKNgqV8kxmNtwYoPhLjaMuU+VmNuSUEpxbeprBLeduGkHkxKNALWH
YC6cAgtFKcXVXulSZOp6ktrG34FioSCdCblUWCi/01QuNUVw3qce8cYtx8uUhY+B
WlSh8Rncal28Hf09cyYAVja4P/6yvPVPAwGlBeC0yVe4vY9pzRGHHUGjazA3Kca7
ABDeg3accgupQjiLvcDnGibEZC5H+HmWhmr7NoSRaTre6qLn2o9NCCeMzmzQS6Rt
lKgFjBxvp8cntbg1edscIjZEtZTMq58ypEkmrR2o0Ekgg72CfcLCzJvmhJek268i
QXzy79YUb5FuMw0rsDFChDu3UUL5WpnIiuXkv4ayo8t+k5om8gDsO7NLXusf5u+Q
GVYAVTDKX0qK5wvJqLLc79QwvIgb4r3uxh67ocNLBlaaxw4opx0awMsSGW0uyZk9
Tw+rgDRu9NBU3N90huBbQRdLJMVIbiSgKf8mhHYwZ8ErcZ+b4r4DJBAubx2P9TQK
fHhmOyr/UKIAwct5vrfcVyssZ2ZNFOaqLb48Y0kFXoNW/MAXSNT+mmdXgkAxEHbE
iCDSvurf8CMkkIlFcD8nHCmkroB6bbwjuB5Wu2XubCsjuxzKPp/urofnpFvBLdli
71k9Dnm3hlF+lw/u9/8Le/68rU/D7YTuZmLtdFND74lV9S3DPFisbnCzbjVYwTST
CTo8kUMWlc04hHiJ/wnrg5JZDRSypGsRVOTLDZBDSZPs+9TMACNvuZGxHC+6B0pc
H8eA4Td8nLEztclLN58xLreWYtNkjAUX1OghVdo8fNHoGGf2a2SFMwKHIE754KCy
hADIFC82/R4ndJ4LwgWKwt0Yq3PkFyZ3WUdOfKRf9WFGVGQ7hH/iB4ZJm0KvJrqS
06uJpR7zm7E/GDnm27GyoRxtefkAZPXL6pTLiidrkXp9g6645SMI9p/gdABQKUbT
LlxRVS077ZvYToNQrKXJTPgYCiKtbv5D1V0wzWNssmHlpw0+zn0uukbkd01ahpdE
u2sJZ0pwJ1NjCjBG3QHzVkEa1Qxib3ejaBF6S+aXyx8kfMFgKPbWtWjHzKD0gY3f
yOI0DqS4byAhJxhkMNFfFMuliJF4j0JrzPnl/i3ooqUN+wbpLhnfpKNdXjvZruLg
egvwKKMfI8oc7DQoW0BRbstwqIv0/3+H3d1slCkwPB8CiANcYBEtopeziwUw2Yda
zRH+QCG0UXefzhMxCKk1mRhxRFWazks8VADKfHRqMtwhjNTBziIPgBseRrDimzJX
jR2/0IXPEv2vTlQsCpfeYR2XA6EagTVb46kb04GFwm+KtLgjvVsgzPoLq2xH2hDb
xkHnPnpGGmoLH+fpH7eA/VznpsE2wStWLU/fRBNlaAoLhIG2qF3EjW7uMDrfhbm6
cj1QkWkiHg730Qp4k+r6X6ZN3NhfOqtdPKSWOueBBW1YAamZWw9Rz7th8rwHTnQn
45x0+ayoa60Yn0lJXokcvSlD1fIaCGT/nq6RQqBrPAoXCBBjxIwok8d4bkXE9UX8
HdYCc7XgHDP3CCZZIAj5FSK43AtzYxwJ+bLpV5kBM/QgB5PMR78OjRCYfjaoqizt
lPXyo71tHlIwvWXcLFDVlGEar2hxZJTQpRs04499u6sQyl2HVEzI4drdMmfjd0lZ
QQWrApj8rEH/9V06Y5NFEkoYGsUBeVXtBduLw1/1r9JNQG6EfGgvN/sRVk8uMZ6O
H3/gDCE8X0m+eoSUPDP+xlTVbyLaQ+UfTXf+XXj69PzAafBNi2FCGF5uLRtY+rH4
0qk9B/ffwoP0ptc4GVdC9ad7jJrOffIDgamgPByUo+Ku2+jvBALd4+mYPuhG91kk
UnzKCL1JoZkQFtoCrnbwn0+z7orKoFZ64D4aIZ7DPDK0nCEcE5CdvVhNtH47u2UA
L79l3uwP7w21LkBH2q7YJX/OwmbWDRVMsaQerVerJdagqBVdGyySxu6qyrKc6rux
yS2f7ugmMEUq7ASLrmob1KkT3pTeawmDw90RLTOkY+OjOhvmLXXyLtoFHiExcrbA
gYZhvbG+SylGj/A/pSw9+LqPxAMEClDMrj98wrwG/3z8aQD3VyNeLbgV6awWaP5C
wE7QMYkowNm4T45QaZmFIuAezEP3ZuabxOuoNKbB6NK+RuyN9Gz6Q1RQT9Dh/ENN
seKtN8RreA7ie9GWAEy93f5wrk0yz+BXLkjMX/Js2QN9O6CUpJVMHi0thprGLu4W
XSBV5MNhoIuEsdy3ox1OcUYPb2r1pUbkvymLy9jeODhs7svIrkpVDvZepIaSeRQ2
RKY+tkjeNdbwocH3l+vJXIZ6a5aW0ta5zbb00ko9bik29DobdofJp0W2Antkkex0
zAoGdD0ax8oM6y1idBFClo7jG+plW/TngCIr023TSoYW5KCuoq5jIkYdzr++cxFr
CGytcPBnH6DTe+mjpEuLjO8PT2onvL2YHJn2ljWjp1p0OIKD8wuUMVTNHCBdL7/t
nCw6ND1M44mG8T9vxgBjTVsswnsWe1zbOsxVsdJopXhF25h5yAsp8/bpGeQtbrsa
KPFSsvsPQfVH0msXGaVtxKjYsqrAOpLu/juCjS1s2JmVOtWRNwzGUZFeb8MqqUZh
MC9Te8G5Xo36zV5RhOIClPXheKCCAubvMyxwxGzcl6JEHQlG1Z34LRGL+kuDM5BI
bGBLJBU/PCIvwfp3gBqVMCQq5PPTlhvWXHIihV6Kt0O9/O9C7ksqaGVSDxlCfWfY
oFaPuE1gUP6rlBX5OM5huiFEeBw56MmLTZTv0+fHFv+2W32VLoip2on+O8j2WbKl
sik4XELkq/AreLHU5qoXj1UzcJ46459S+Leiqv7X3Nu1rI15sl8QofaLHARyfQjR
CSKtQAQ9amWKAeSTGxHjrrvfs7mvvUQ8AKsmARO7+uyTisqmtef9wGje1K1GpgNe
QrdVr9yLTLdw1LW+ds5XY6CnZ/0Nd1BJ2HHfEJ3HcM+dX8uyeDrZ32/AueOehJh6
jkMQmZyaZShI88OwsH2dIjaHNGruMr+PA50+HPw8nQGG7ZSiz4aQcujms8CRHdhl
P6t8wzxfM8wapVeIEXf1pjvRCsaTwghMKgKfajJO/Tcm3A0olEE0clJL/ZYn8jnP
8JTNpgn/8H+J69CyOJBtLRlsoQ1r9fNpDS6evjCrhpxwSxR7Q5oiHFK96POecQ+7
8twTYnacKkx0XarBI7floesMkW79rhD36KwtuuunmgIA/72oHetc2z6xyMUx+Yvr
Cu0qhYx+R5LQ1IaeGYi9ztA+Z/TobSIYdmqkq7NfCuWMv4ZDs8v9+zFVGCU4mPPv
XmIeCA2TTQ8w+obNs58vpn4603o2fnLdt5W0O2yXLDMTnymTV2B4zF+Su5QL1wXV
brNcNGvgq9l+RRjkAhFTSvT6Ge1cbb0jl9594SsF7Prf8Jq1Pm66hsCUWH/+YFRy
rq54MFUAtFdn2lfuMiIFBl6JqzqeiCMs2HadnTsr8ABQ7Wgehy6vdVDRJr9wM+Va
8ucDGA1pSDkVaUwqQYnOgh0RmdTtyAj968q350bXCGF13DyKTJSRNExn3iiO50N/
ieBprIjaOxBh2jkEqDrG4HGUBCjzhdNw/anQdu+kkvpibZ5rlvxoJj+UZQYBreIl
NUrCIDCzGH7eOIw7pC96LKl+J/gO9hx92ALdBdstmaDafXT1+Ui9wALtYyuO8SnY
2d1FDYfFTHwE8zU2DxgXnJArjdz9+axvIlO2jpupRczb4SaczEFQT50ESrBvgXG6
bX8Tt7046mLJ22yGkbyARyAXcS2sio9vvtmK9yd6aGwm0ir3y+AJmmW7tqcBkCr8
nZThb1erfaPsktF92mi9dYPUsRJecDaBzgXNlT0mIEqFpjZzwMTwJwjt6krh5G3p
+WrF8XJkfawdyxPKdhiRZxA9LFTZT97FUbRP/IGvr+PGWI3BlnP5aggXo3AdEWkE
ZZ5KVHSTcFgwttrwhhJnF2VgFdtgKQTVklt1SMoqy20fs+AXYyRW669EqpoEunWe
nKsMAZCs87NcynxsBrFzg30tZnJalQWTbcVQ1tLj47suqQmv8fAeVtXrcJudp/6k
aP6C+7UFn9MLFVroond091xUqYWdyl3f2vADy6OzsmDuIAVqF4iuvaON+XRurFF9
ukQOrrant/2fPqj0uFmyYYRVg4gMJ8+LUNrsF7KyEfxrAxM8DaVH2I7ROk/Rl2d8
YrbH3CWUdpkQyOoc3FeiXuHy2/JLM/o4w+3AnRVp7LnGtwKnIH03RR0exP5mgKQN
EVn4eG2HN4VjaYvAxd20bi4NZUrgvev17dZj7gwf6mOZB5B+selC+TzogqN+gK/W
kbwiD5UW+UPHhNGpWm8iEEtCJ6TXVpjs1GnHkY6NqfUBc8WWXbin0A6Y0jBcmisx
rv72QjqBQnXLI8ThlbaZ0rgr772nvxZunwmjwJGvm+HbHuJOHuRFU3yNRO4Pt5cJ
cQAxsEYu8oBVTTa48dtYoxvgI1gALq9xlyPT6LfPCOOhRFpph758qYa24y/4F2fq
s53+TUoaPw08CUfXtFlK7uPwJ6GMN4E7k4PKdz/H1FrR+a40vv3vGiBte1lIpVZr
UGTf0O7iTVaexJf6N94TZCvwv4LYKQolJEqVpXgJ33XhYnTq7nWkT+r4Qr9Rdqud
FMTgRkWuflHqnCdC+7UKB49fMi6trC26dzQEk7PiPPL4v1RAJFy/dbGUgci983PJ
pVqmUQSEzbhRgpdUndmtmqoQTpJGmnASvAB8ELAvBoWzfFqRS90aLvIJZmRfVq/r
iJY2q7qrzgQi0n4qPZpAQ4fjy8MrcL7zIUfKpeiSjYAMp7WUxmyhSFdF92L/84eM
GNG3987cBxQRAwp1QxRLvuYVvQNK8Lo8a++GS0kmIX66Zwsduk1LPNwQyBBMv/lF
FedMjvU9Il2xl9qjheBzqK3NJvYEY1wNcSu30tWcqyTbhHE4vZyQRxnev3H7P1ZF
nqTn4WR1+GTlgiNoLIi9/zsMcjvObDOSBI9bEjYyh/eagDfa7qgGtVGc9VYoV/ji
94EwsyY3ocCNYS00nQ/dtPvWCFbTuC7HqG6FsH4L4O+F8HKfYXcFtZBF3QLW53tg
vENYmUQguLAayOSNHYZuO5lOKgq2dwkmsmwzh2O6Uap89ljUZp5jqxDaM3HJLvtb
TqC5xPiFbQG7BxtQxZUWB0w6RvF+9vWDVv98GiwanWmIb1l0vSzkrPVGSagF0uum
clIteXZrbh7/81VdnuHTTGoE38ZhnkevKogLv5/bLgP1aF3VeBu5PpNDfWc1lomf
JCkZQXsyetsxb3clz6G/FcrGGkWK10n2jE1mw6hU/XaD3bSbvk8oOwjMqopzpX+e
FvWhaaL4v1kY4R7TB/ZrxoILnv1SxEMP6dyPwVhulygNneDSzJ0IyxlK2Y7JEHiR
b014TqAxmv82KqT8iGUSX8Is37ZKwOVmd3v8aeAaxxHCsKo10/TaifZS1z6ZBf4p
IsLwBtiR9Sw5CVTd0o4u1rv4PQytz+KyqEhBupfoZq5bb8LGt5wP/uobneAGfbb1
HQuTywbYfquzjzeIJvcrYGAR/6CSB4kBB5jdkR5A5XzI0Hw8zllLJ5cmqz024eb9
lIjvFIznL0ZEtEH8MmuDOP3RX+pBnXKfLihtPkCi/SrA8GqVVR5ONwtdE6tqJicD
73qUOOd7Y3wHKl+QbTXFf90f1yq6lfN52Q+clnUM15e9ptGxGyhzMfVrfoVu6UdD
1HWRWmtgQRZ04W8LhZ/drYsoGayYylwBKtT5pC8We4i5sRM9PEllN+N5WK17iatF
EbRHFRTYYui6cNlqwjAOAj2lOOVPw5S4IuvtQKHy6FoZ9g5RkmnQZxkYLDKkgL7F
hXeJdYk5FGL1s4pJFm9eNxArM5fO5L8pW8V4XL2oyr1rUfN5JAD6pHHkh9EwgYUA
SRBQoyPqOsqSNKT67NLG9It0QRiQGk65BMPALLguhvPFbrWdL65nIU5XoGjWgOu2
Ot6Iqn0UtMabPTPLDp21kP9M7tvnBK00d/a8sESwddZcAIcHCIzaRyGd4Gq7/IVO
tIgI35tsNC80gLzI2WMvC4iPJ4T00xTIhfPQIQiJLpc4r9heurJPUuh91rYPY6+L
XHzsEHwLwpfoCaMXHNKxOGUdje3cbJ0sqxUWOcC6nmbh2xJ4FUrZeH0CBE39uEd+
+mFUeTzb9fJ+3VPHA+fodJctoIkaa93LE+jc9pyvLxUGNC/hytCMkw0jORIP9YFf
ubr5xzlDaOw287oyF9Hqwq4ErqQOqhOGVYIDhL/8Et+JiZrr8Bz+1EX4fXqlnMuU
ov6mDVX78Pj2v6lpMP1U7tuqZ5sGIf8OvkRrRedO2DHyzSmInnsfPOVAFowvNgdO
F66tH40g7NCwmjelS0V+GaEgZ6J5TcAR1iArxYDtAeIb3e1JSTRpSI0rzcO9pc9I
wnIVmBKF+x+SxHsi3nTINplLBrzPAO4py7Dq0vSLcaNfrK2CDo1jFKfWOjVGE7Vw
nm157O123IJgP7t37WQdq0541EeUmQj79KWcYZ7VmTb+zUt/8H1v0Mjm14jAt0Ph
fKp6mrKWCdyCuBoPZimE/koOaciwuA2dzUBiZVHe3mDAuJo/9vqkGAxL8iFxjlom
hCSBAq9n8Evbw/t910DQR1biVmhMlUGjwZe1yX9NxdD8hDtRZ+6JPji+fWAoRveV
bW0VtUvGnA6u8yVRyhW7H58iTQ0rqDDVVGdMJU/4G10CqKTem1tXxcaCaZRIK3Ur
TFfB+SFFQOOIZDa0LiLxxhHRWASx+ZTtYmqqXAdlNX6Aq6yC2BZFtOM19AIUkjh9
IpA+wRDQoQDtbLtJQG3/vCytfI+sPmujKZ/L5X0ypuK8hJX2q8iThKq2Yvk6VMoe
viPeKj6cMANS7Av7+BxaRQNLMg0tUuBFbl2mB/8WEaSHfv1tR3X6F5oayCMdm6SE
AeuJA1RwA1vlB8e4e1dUuR6IztfHTyahDh5D9SjTqWKttFDUk2MJ2yQ0A5BmRhcP
S23LAiguHdr/qyxU7t5DnDiDqROjOXFbRGIwXAlas8XuevkzuDnAKM7kkH1Q3aXc
uMr4gLvQau9y/aRNr9vRrd8FvkVfbEBRoSrJ2S6hvOlUKF7hWRrrCkznyenBcwAt
VG62fHZF3wYb810ghQwNM0UUw+oncw/ws6P7gD772oNi7VXVpP0WJ15mfcqKOCnj
w6VG1g2uqoiQCa8ppP+SQ7bb/edQqSY3Rus8DAg7cNwPfOkQma8EbeU4vnfuwOPH
uRfC3ius/JeyQce1ZAzre/nH3J2idglErfTT7Zjf5FY/w8roPH9PxT067EagFv+p
De7554NPZqVadBMXPGTf7PNTs1vTqeFslpKJsj5niNg7B86pC/fMHcripjBKm3Io
uUhmUz8qzXDG8xQwfa8ubVcjbKvuPHckhWqLtGBSHBzp4zSCtZ7+mG41U1+bOpRs
pEsaT/PtRlI4cNJaDqrLK2JoOylyug7K1ER+s+Rdq3uFwqdpz+yzVRJ3EE9DLzRd
vnFwGu+QXwAAiDgHKZfZtQccIPice6nFhySsaVboUeEV17xOJq3dSmCqKt9GNesU
Kq5JeIBN3sikA8/a+Jg4QNQzOwwTRUb8ZsVJ1F5nIX48LtnhS7u4aubnxVlM0Sm5
3y/6KcBMUYxPrG2ITuPo5BnSdBtipivGzwgex4Qr9iA1nK3oj4L9BCtycJ+kexiL
rcWzvu+A0luCelxkESlAbvM0VjrpOxog4iARzh+VuH9jfZ97YBpoval22FBOXN1B
fz2IM0lipBoZGmgYcYMrxLtGAWG4ejKymNOVcCUJ89+xbtx6vgsrkIhKKBeD+Z53
2KonikFqET8OIe0J5ZsWoVu0ei4nGdVv+8O1/tB3Zfb8hinb2KkONov1MShacfef
zGvYyY3/evW1X6qYyq2C78esCDtMTtOzsYmuxWZW8S666v8LyMCx5hLxyfVKUul2
RgPgpnx+EOFO/pCmyRFWTEF2r2/cehy9VM2h6pz9cvWQ/hJuR9tJl7EzSQpm+4XU
BflHEJk2G8AgFYQINJuWcGNF9X+XjlU2rZvJlr2dZL/bqOA16avCWhGwBjPt8sdE
z8o4cX/vD+O86wY3ZKUbE8QpSUUekXg8bvnSjdAN2T2yeBmGBb1r91MHAno3jIap
n41y1HRzakT4JikLlyA6pcn9kZ+QWdC5yGzc7lloK3y15YmTXPGSYOHX72n/oMNN
pHVdP2u74ZcKbCCtet44EhDfd14tOMy0OwG3fHxqsCeI5NqTNXx6RCfRF5+U/Gnk
KBL4/iuupTBX2pWIkm3GwEMH34FknLj6KT3E9iRKLiQIkv66m1OfnguYBft438jB
XLsw6qh2lxN//yoP5l9jPsI6oXcaao4ncAXyrXxgIhu38LlrgprMWMMqMUoPw6ow
eoDigdlrwc3KpescfaaBkNB0hnCnluU5Je4DEOz5ESB/Lg73MLInhIkA9isjS4xK
sEP8N5gR26I4l9q79dOr274YSdoQCtHitWYwrZMm/9ic02l4dpTFIOsbA/3/Apps
cQVjP35W5Lu3oO+ggg7RFpXKVD6Q3+HwytBpd+zqyIPEPhMZ0p4pTsCa6Sv9huI9
SHVaK5BHmt0K4bjD1ToF4PgZNFWrLhXyN9x/SfP4+9JuedxNNZ9j+behLfILWz4r
yPkMYTyVgMVmvcsaoFDn+gOFteYmM2xuVrzX0zUNAUq2pDePOK9a5wigf6EgCvdf
Famy7pUWnQSJVWMuOw7/Xx+B4DHzVbJtuAr6IZKVLdC4FX27gen31I0EjO9mO5Zn
bj7hD50EvGvMw1g8Ph492LRmlHApMXQ03WdXfKdyR/KHOejh7c7pBOCXgnrSCIah
siHefG9OAFjz3qqjF3xbSQaUO+GHnHGgecRDBKjXsI/IGHN0gepxJ7N9zG+fuptZ
COCyCybv/e6hhfWSyW3fa70NaT219ytGge+9rEKYLqS4M509GaX6VHp4+lh24gJ4
FRmf+kh19mlg97hn2UoRatfMYpiJr6E6bg18Xi/leij88hpSCWqCASxs0M7sgb9O
1CzjUN00JfMYRRCcZpj15i8y6K3SBG5AZCOgCJulMynGa7VlFjLWwAKazzmNXNrf
lzDGVikvKetEvmLFG6rZCf4fvf6bp4F145NfNCUIpfeyTJYzLFvMd1xLiSSHLTtK
7I+KCKdGbYUZikiCfACdjnApLUFmi3WfU9j7MF2twEkpG5j2XbEktEn4IPOOxdU3
1UibX3cdYrVin6kh6oNS23Pbf9xnHB4odP64MvgxQeyGSA/D3moTd6CwSteDrlcL
n1XQ+WI/rhR+EiezJie4kfJFG8soMYjgLxjnu3Aa+0sCwslOngTzyjVJa0FBw1Ll
LSsdrjlwWQs6Q/Fqo6ROrrNMb4dlLYYUlx6OEK7xJQivQIDrB90i8HN6DnvaIh4I
HyvVoJ08xhxfmRoNgbMqiYALC9kY5xG/4eDYe57MUiuInbje4Cq7bDTYl6KybUQE
uF/3C5v5/U/iWIHDHM3Ll+1Av1Kdup+r3DdePzbj/72iOLVZrX/z3BTQRvG+tt6S
suVMC+3sOh5iY7DuS2bDxu9EG1hxCWuLq+ohcgPnOB/KIAk0IaKOMXmZXbxMC5Mj
/lZSXPwSvYOlxNmQhXWlxFoHto9RDvTPe47vu10+DP6skemEj9kP41fpRXvyzFrd
oiDVGA2Aqmh+FeElj8H0L29BhkhboGs/Mu1K22l1g+94m8LUJ/vTb8sgZ8k31VgM
OoTwNnCFGfdPrCUkdaI1Hg+RurjD5kjjj47sFMcp1Fa1iOt0+2TSYK68VCD00s+x
Ws8z00PvQ2oKZOCjdCNQoMLHDAZC5q3O2peBp9riQXcM2gwan+Cz5spbS2JquPKk
m5nz/xUPoCBlEn2+/3wB+a8SkEsgDI2Uc6ErPrEHqwT5zo89K7mXQ9/42r1rUMqD
r2kFJaKRJS/X8tsxpvsMWNtatARzZU1i91muZSgMz1UWe6To9O0Od+XZbTGdufJr
ADGcHVGtFCKKt/BPVHQ6vrQEk0yGwxsBLmwHcfeHg02hmi3gTkQZyiZe1SA/dxZB
AisJns2Vag9U75c9rm149MQV2G4bwNQw+/q3mO3hwfR0DHjOLsM+RWYnImeqWlN6
VaoUgUQzt4w2ThxA6q9zGmzJ8tlY4Q4m9O7UZcEKfcccbIOW1sfyJMIw8YE8K1k/
czBxQwrm6QJPLJSYWl7V6TNCGnj6If1AKXTbcAArdghbJT5uSv1pzcXiopS3/Zrn
g4pWJaId1mcG4q7mye/3FCU4+00riTS1y0iIhDEFKwBn6DFYKhNDvTMYng5Piau6
o+ySgol5tz8OFMeyFjk+QVcdDoB6+glMiMIq3a+Aa6faMee74dY83LHEG3dyUz5Q
D8fp2kHPtdXb9d7yBX/JntFhNZrI84T1VVak+6eF3FR4n5+luZsem6U+2Yl2vhAy
FCauJvwbyDIRlEqheoNk//CtKjYC3NGmTY1R8bSmOVlm88QwrwX1tySIBcgdjQae
op0EdXi2tp8Eoqn8ItI612XwKxqON7VO2PwSjnxZrflE5TUPSiQmwIGTG5gHU5+r
zFvZXkGr+YjyuHZaXtrcsz0zIQoRKoRYeMB8uFx+VPaHX3OnTvCXy/96g62MKPDK
a/+WO8X2b7266cbddIB0r+v2vA/D4YxrHRrNWt6ac5wHU9j4PyCYjSlmTVpwzw8r
S+V6llZZLzlumOwbx2e26uXO/1PVCSaLHthmUh6ydVZ37nWZq+Ix3jk7BNj/9OHn
SUN43K6e/0cymvotXVZJjPLZuDABffQQoVevT6t2/SJ+p3OVVFjHQ6zpp7oIcdlq
bsyitCMC3bJwKEi5bTosyJcElYn4Iti4hAcV1cpNsIwuHfoCQO3pCju0/fIXWaqn
zHhUnW4HU4uDZRpUpR0cLwJ7K2swITwo/z2jJj0DnTtLgvPHfqtb1S9VVgAcMk6u
knOS3/95SM0YA6xxEMJ01EeqVN+zk72ZjIQoLbMgoFu9l2T+TzVwzVnWhr4fwLaX
GJVQQ9krlDUdLfNVNwSulgG/9kojcLyI2ob+y4rWMRZFxJrlSMAmiQ3ODxSy7aBn
GZ6/1Ik5i/VGKF1jM6GXFxh6mAw9ztBPvlmUSJPeqgjxBUcQ8WiSRCWh3AlOhgyy
AILfCZsUJBW8PSj8PKrT2B3pYuDCAbDR4LtIJ8I3YzFWCzsTiimTqcKrKJef20nH
5xHd9bifgaCbojAywymEK4PAu+St5r4JEEUMnoWVB1ZT7voQ2OxmrMA8ZY+NyTuE
dy0/laPLbjYjVW6axga28cp0IIViPtBrSQXVmUDMyWm9j0/QEKH32RwqcpazDTFS
KDygnQ7UEkNmnJEOdNLGMD7YXhA1hIUJ4PaSlQb/olgLNA4Q3Giub/k1Zmm2xkpu
JCYuoKBdabjTmGjr3M7ylMX32asP2RqAa2L8KGF8jPR+DAyUP0G0Y72VSe4Wl4a4
Fkgdkqqn8HFME3XQ1koytH8p7wPJqEcqwwa6mp5c/NswBe5D+LBdh6pCuQ3y7aat
kxE+cQ47ABVzvgwWESNJCZrQ3byrBZLW9JzNo+PSmqryHGcNkZYLGxQYDpA+rtL6
iMl0ngxEP/ntVt6BubuZXaM98WCQnMHQfsI5WPAfsK+9Iz4in7YnKQJOl2harTT4
9VNwY13H/hzdydZKwjba+6429qkBE4BmuAGpfaGnhQ4Sn6kwvfHJTip2BmnpoSPI
Ayfq4EG6g5Ti6CLg2PclNL9SZ6NWf2EgxGCzVCN8k2/+MgOMy4IygrozakdNE85l
Con9PXYQzzEgd4erz3D3Sg7i1KgLt2hnw8d4C+c1RC5UELqhz6AjLttkZcslmU2r
USppNXc4pSUFaWP9IaGVzXcCHbRwM4DbMOhKBEWI0wmMw1HZUFLgi1sLLe5ZIp0A
F73UMlmWQs9GDNDhP2MMZMa811lXudPRoLITIQwoUpBPHx2M1pz6FpPldSr9rtTF
ViCeafSDVcFX/ZC9ZF5TaHYFmJcogBEn24bkHAoeVHPRCZsoxdJX/L0WeIbby212
0vr/tHZUUmC3x2Nw7Oj5cj1Z3R2Cxnfn0RNZ5YI52IKXCEUSYXGqVrwl5CJLu6OY
C7tt0BTMSlNO6ONQyJNBaBloQVQPC88wP9FN1bL3fwO5dlzrvWPls562PFWd+y12
WmxaTslHivPIVGprwg85jkg0woLW9xpbZSHbtMA4eYdGAlSDid4sAHMpo1wWcRcm
O9pBdPNOE8ReLGbMSnZbcaXyH8M8UDY4Rg166aFzy1fnkkjFMMA2lQMyZrwuRq+Y
D6DiAoAw3CFvnu5VKls3RMn+oLaMiux0sENh7NATQeuHgem6wy6Yn2DvhIQ4VQgZ
9LBhQ6gFB2q8J8SHFzn+d5IN7CFLg3I+SED8G2pMrwB3jk7cd5Rk95otPpRGQi0G
35jFNxMTgKd5qBtE28COzCg9FOgVKNsdeSawyXW7RfBtkOvgZ01D5PuIg4Y6Yygc
eXukssinnXTxeC+CPTj3mysMbaDCk/Rsq76MxIRCXT3vjZ5g+bdgZdzDRstKCbgY
EvxRpxVGrDBeIj9ZTr/2HmHyYqE7yO9vdRwkNfdb7XaR56rZkpQ/p3rwGcGdE9wP
wzxN5tvslFYah0zCR4Poh3U3xasaZ0YIHiYfzuK+Bzf58pL9ug3tqOdoatREL0r+
ZgfoEp+v0jM5HGWemtHbveH0K5wfDw7BrVyyt3dUTHo9JQkBbSsqD+lKpPvpmP3E
VY5ImRWgSMaghLvuBlhXbqCXWiOVSuYyGGWAibWIZ2XYHcHLP5BbZU086c1kTEcZ
KtKVpi47f6Y+dVAvDZjtwtm1pii5jg6GOoFIAdj8o7/8D7eOBG+cEJ5hlp0uCT2g
YAL5grf3iXFHItU9vlMFUHbJnOGAGVXhKZgXkeGkCQFMSqSJrh4vRUHjozJoV8qO
wPC44OCMrNnPDEz3xp2iH5RCm3EYfp5lbmYo3F0zVhZRHFipmvfDg6qqXOgcd0AX
pBcpppybPm0ePk/inrwHn//W7TxA0CWtyeIs547yU1luWznQ5A4Odf7CmjCpDbKh
SOJ5qAZtYOHunwwEp3p5ybCNKxLe9msjJ1EmluSRU993TaK3aJNCjZQnKky7Irhw
y0vltGfSTsdEavGndQIIAJWG8xEMFFrExw6W6DxUANn/iXNJaLhd+twlRvrGnICV
+PLOVS/8VbShOo3sv5LuVACW9JAoEt0CVaERAO/jxRIEThtLkE8cnG+KcUbvz5N0
I9WbKmcCHVUv5bBX5THx3kFF+LQtefWA/1Le85P9aL4/iLaFIhS39gYfn/eTe2YR
XBKD0TSqOMLZdljV+RDzUvF37OdtQ/soZXZtgRungjyU4pL5XDxIMAGscB9jEo00
7ZO5scwTGoALnJK60b8zNH0JX27QS2jp7BVkCRL/caPNWHJGFvzChimL+2Ch6hy7
y3HqCKaWOojC8tVQ4GI+4jfwtBuZStcU+nvUDd6bpb+ibEUpf5Cvv6NQt/yEj2m/
6dNwcnQqSyfwjOGL4modIPfvjeme5c5SlYeDzMOJMphBE06aKxLu6zpz3kcCWrYU
6ugaecUGPrRWX3zYVq6WvT589JI5fNIJWY3DPFv5Lo2SFUQOZ8J2ScmvbP0P71B+
BdmX8QLwCS1yeEs7eMim5ZIyUuZ5ohckjh4Af5oELUPUSBjMPalpcNo/nlyWWl7z
zI+VXQo9MBpOgzMrN/wveLnb1pw0EjDCi8obHkYVpnr4258tSp201L1EGAaqhN7m
rMTnlICGEh2LFm/d/DuLADPAX685FDTHrf3GphxKA5aSnfj0m6NhADCpnjcUggXP
5zuoa3BXrJw0fCC7x+0bPYxnEVxAJ1YNnGd9utetHy7+2bdt+hlvs7gAW/J9XD7l
2t+XElBK0FYZRz5w4p8gqSCnOTEHkkmpUfHMQl65MO7zfA8qvRX7v5lsxg1innFG
8arhKQ9K9p/mpqeTOW5xn3o5CI+mEXE4chDEadLeecKFrexwX1s1l029vKPA8X5u
X5hkgvbDZqvvNhfohAuBiHeUNro4cyRGfP1Pf1Kauh7qur23M99pf+oKQv97/jyT
mMJobc98ggLyHd6cf+Shux42PMdrDvKR9lihlVMHbjh/ntxx9IG+337W1hx4rbPC
3rnJyFF1xBZ4K3yQmoEBnxr9iXtT/6GZYv5HgoVvUVxGRDz71LOn3aE8CRNd93/9
6VmMF3FzLF1JyoYdcz1b3UDL6FXb8nDGsKU2FtA2QPIl08/K+m0oEZF+Uc+lyqka
ORmcQZdOTWhPuQzsAQtrdibB1RSvd/kBNq7Ep0+ict6q48FZsJyN88TcdSk2mP38
VrS5ctvB8bEZLDibSkrBN2IdOBnmjB7kMVsZsEq4nGztETApUiQBoExcolDNMtUD

`pragma protect end_protected
