// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZLkEKV8zSyE0jHKdPoB0FUZZHJ1K9MH5FvDMlySQsHzMFwzRaowbngytYwMG
e2tM2SU1Rtlya7jbaw9bxSHnevQec1MNkx388YkQcNuSzn8TFBmpTx2H6zEs
O+Iv+fozCIfAW0MjGK0s9qzLgirFgVF74LOrN/fSWanZMB3DIfY8EB59sXLr
uVnVk9WqaSKdRoAFElEKikIoDtl7NrUM4BAFUFycg+EX3L6bMQ0ozgs+dxd9
RAGE81Ah0kSyUZs+fiWFguDemP1TYHM6ctePW2Z25kyYwjEO+xwQQORecH+0
tzxJ8bsz5qXyJ0+8z/gjw4IG2TiYVliTR555qgJziQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mg3yZ67F6+inb1gM4gwM+4SlppT7fcoLetPeDOl6Nme5v3iyxHnjKqe05x7t
ApYTPLrkV5SO+7Fs5wcn74FkWiz/OM3/zSkZ7I8lNVsqiFteAuVFbDO61Pqc
R7os3cPdxSS/+fu5g9/0TH2tkRlV2p1ZwK8JdaJbvKF4jOD+tD+7kq+X4RMh
YCxoQ/nQxt3qLhlvouUH3q13eNxnEH0DXbbd2KwqX7AN7s/oUt7XlaUbrgVM
IHsQnmOgTKnEYnwEvHuDVC0F7djFYEQFrUohTw/kuGHdc6uMFYXfKOw/tWjI
77pEq1Y1HIQHN5yYEEq+0mF2T10ikaY3ZV2d79csMg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QJHLuuXfpBiX2X6zVXv3Giz9u5ypOwyspO42PgDmFrQCUCBCbg4mA/XA61PA
oFzNL0APUbrrbF5sjmUeaatMACZMQIiE8qmgZW8NpfTGsYFZhs1zf+FYtZkx
LrzE2HWKy9n3lk+cU/z2s9E4ntp7jh/6+07C5ar5LfVlyPCdxfve9i6PU+ha
7+MtY7aKlzv6Vt3yGnCvXo8UWVFzkPa7c32bGG7BXDR9m4IWhsz7QX03EgWO
8qkEZ8vU84UWmiWjf1lM0PIpGBBluiN9jhKpylpQGApThrtKT1kYUvWGj3DZ
jdUMb3vEoULsbLXjpsarn67It3coSXsWITC4ZzNeHw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PuEkaM+5woXuqJK0Bo0zJk3yfD0p0riTXeF/lO+WYd+Ur5Hz76GsovvWPLNn
5AZdn32EaPFlVapfdSlTtClpAYqkkxq8VktNiM/hV0ruqsED4XwRSLOt4w2m
B+8tGpSo34xiIX8d8Qtzrulm19aQQQTvG2Uak3e+CAOok7XNhxk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pJotaof0jKihEQuheYRxZy584w93iBe8D6LfeYCHClk6JWAYNgk/rPJjCQAU
JSfkxkTa/lHDUkoC2uzJnKJWp44s8hUboQ/7CjFhSX5S+azYb8ZBY6X51jpc
Se45eeO8Xb/6fPv+WhRMiWmGgEvYA8YTDFrakbts/5B61XwG3aLU0zvfJGM7
0fHj6NZuIvzjiYKYJsBcZ9FW7MthBuem7bhFVjNUIAMcVxRMLZE6vbw99XEh
lHWVk4FOt2fXFmiwl8sCCb192wSwccmINtFP0m57QPIpE+5AF6FH9FPWHw27
nYNoAB5rUeXIE/6AaKNFQxm2FefihA4+/fjvQ+BkUNNciwBAo5o9PyZQFOYH
PKthBkZmisQ8T1WZpMOlv0I/5B34wVA1cxiWsJa12dBNUkpgrOfPzToaqY/i
7W31fsSZKfMjOjIGz4FrLCPdU4CaMR3weQY/1mdetCYJXZgo9Zjfcc6jsDSu
OOIJQCoWKG7omRpzxK921Ki+7xrsuBZt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
O8ynp2MxYdZ7FAp4HuKy0sdfDBJ0mwgUXS0xiaPwN3VJwCgyVuBD05/YIkNO
XotAISheNJAUEky8Li+QSQvhu32d0JLTAy8uoPlguswEg9LrtsZ2osRo0hJ1
msWWz3lrRn1CIGH3LySpwkr/V6ueO4X8raA9YpDIX4lXpwDLIqA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hjeZm9l8Ic1TUTWDHrgf8+NS43yIqG0vzEoJmxp6EtzxBmNz29We2utQK27R
gQIl+1DL1TDzv41Pzt3pqyu5Ds8Qyfsqcsy3LZwOodU1skkB5pX2+48AhjAd
GYQhWeR6oAUe4Zu3i61CGlqPHVeotv55phnnksXJjwAgKtV9REs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1120)
`pragma protect data_block
OcjwhSdtphKV6ZFFsc5w7DCu2pqu7h+ClfZeFki+4I2jTn4NPraXmMVVLMeu
cGJ9hbRnXIKRaOMIGFVzX7kT0n7HIgT10GQyEbcse9ZNxxHgVexcn/FMU1h2
WZ29QNaeOVX0WcYW4c401gD55WgzwF/7DEaC1xs5EGZEe29awsKB0+YQ4AZb
5VrBHna3CGaBVUEXPb7GcJiFYKSLitJwPmq6o0aFwHS8KMT4Rjb3qW8ck8kK
V5lU4EN1Y/yCX4H6LdsyOosW/yKLqqCFZS0N1Dw20P7ZVyVNJP+EMRW3gcPa
RTDwpLgcz8en8+oJChykAZoYpBYHS2lDR5IoAUJwSxuae0goo3Q4Wzbymta8
yL/gXPr/uYGHgJQGZXyLuhwz2dpSpmCqNJ5mEw8FRj0ITkCkH0vYt7+29UYA
59j024Cxwk9in98bp+7NVcgYjCjFGhGTONlhfoxwhwAlrDg3F88IidPkZDsS
msoPhFIRmsOfM0AAsfu5n57WlQOUDwf1V+ikYgaA2sJorqrnQh+t3M5YmxbN
jd0rP+yNWFWJT/Wmur8DOPa7/MERH05s0uCWCfQCJkmFspS9NdNApb6AEy/C
K3AenfxcFdsRrMXxIraCwPZFYSR2eQYTLHdKDg5N0anirprYg7OeEHxHc3LN
QrQ7Upl3p+tv8xFD2ZIL0mJDOvUtUBYSThtxz9kuo3xgx2b0cZ4mjpelDHhB
DH7ZTmHI1Torw2RwNJxHU+933ONBHNLXx9ltLEK/EEXQwQOD3ex9UV62vRNa
UCcTnQosYHrZWSbU+hoIr39a+eGARFEW65RPTLxcpTaXewKQge0uXF4qp7xh
0pHPrAUiE3VmZ5aEwd6UxfRknQHq2jRpAy/Gi5GtCqN48/74Ry6VXArAC2cj
51+if4TXqf1qh+M+VwNxwNfMFVGR7uo8vLZUWMMnlbGqoq+pgSujqllLIuy9
2xl/vyCaRGcK9slWSGincrZsCsMo9M/clrU2JkaeiFrbQ4a6hVwTFJ1SFDai
ZR+rjguftJnsVzzfDeaKmjdI7ZKSX6VnwEjZWjeNdoY5C8ZcZ4x8D8dHFQ6i
zzdbty8vOE2LLSBerHYdt/3O7hfZs+e4sql1Kl00anzIoFouqKXuMPGduncq
NnEXz6o7h1lTlnN5nM2CdTuL4d29KlJDg2otbST7MJfOAxNwxRzrFLzp1pCZ
rXiLghv/kQIL+H0dxd8esrvtps/9KSE/6TXSNwz+WN73W7v/M6tlboW9ob1t
ywfkzFPdGfDTMXBQ9Dr7MyPU2UlIGgcaOiOroQuDIDR3AUBMdEHeNhmxFsY5
By5DuLcYwjkiXyr7U1KTspLFg038xbR1Hhf93J6OPZ15QKzZYzZIZLu9dWdJ
6l9h/sx08UA9W2nk2zdZ/5YfHWR5VO0zrAQ5YU8oOewmU3dxMqUZy3yW5jwG
lQ8GU0MEfUoI57NRpnKm0u9qqLSu7EKKj8YKrsqtcuH4HgSyusi3XA==

`pragma protect end_protected
