`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
EPI9UYGt/KEorOT7LwpjKEbB5tnaQ1wS64IiTyMNMPbFVjgGxOv7STCjQb6ObpKS
Cz2pKZgs05yX6Y8ChngCTlrmoyaXz8U5Mv9Z7HSeLqpE4lQTAhSCC3rzFieZBes2
UAKk+cLQ/NOwtSQYAOAaB13wwuf0eBjwcn5CCoIEADU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 29440), data_block
vHYiY2I9ZEPcwnoTLTdETPJbLf7B+jJqpubHnLr08xKwzqPQxEr3VsB5o6ce5wNp
6fDWMHF3/UTIBvJBo5l8N3RZ/jKq0l8MWmNgaNRt3koPQczWEKoWYMQ500BoDElS
X9nSh8RYEiRawfV2sXeU1sbrd6rAR7vGUlooACXeDvDIyOAiZa0wxa8q8iWTRJ7E
R7+POTdv7pqGFGDgYW6JFPg5xvq1h2ZS9zi0sh9ifXW9LimLa1Z/BnbPdwaNr+Hr
XSzUXU52oU6/K+iWuv3aFJkSUldWdySxZ0s7Wlx52BxzFjz6Y2xC7FAX5SRIrfz2
4Rx1svha6OEjbI686KJ3t01NBzDmMdthnlAnb2Lu7pTUDcIdfQhLFaJJAAlN96W1
obG1ePRDlWCCQREKB4yaOnaE4Wf1yn+Lvug4YsFR+yQ8apYsXqcp0S6pY3I8G1cz
bqCCKWpYOEADRDEMTVv6JCNPVnVg7AWgBO8aTOHnHwkmyUc3QmUWs0TPCbZMOzZJ
e7cp6nJpn2vxXrVURAJxx2GTVIitFgsojjmfLdQE2jSwevAVR7yT8e06EyytvmLB
zZl6bXp/9ewx2HmlqEkm1WWC2LZrVUIlNlplHMQ8NEqOlirosflT7BwQESn/n2Av
CYAShXVaAwFOAlV4TlapvgpmNBhN496imDx+TKfgftA5v+DLb3ql+TrdL2aDNe4a
MhxKDNIA5cEuAdEBuAyBmCtP1KXT6yfuntZSEpmhDvqag6x8CdlryRP2rY1XAiNk
R0RkHXyj7iLyu2p71129SzKEHY/HtjuFwi5T/r5GUNicw7KixoRl7snUjxyzD8QR
hDbdye91UZY9jYO++DVQV3c/wXFyzK37RIdyoWpQVt9v6BOEoKP+5rMP+LRaXqGN
5LNjmf3hWfXatr0pxMZmsq7HvLCdTA854eVAP077lWvfVHoJNto9uPkJ7KGvoCHz
NfCAz2htspsiOb+QT/fI4X1bbP9FUBnTfrNROzwd+706wsmw5CVdhlXKjTr6wevQ
+iM5s4lSB4jhMUVvFhIWEae9G75xBKALl37I+ywXgLf0jnbIQkIY9QACzf50VzbI
4TYUzWxj1UMqwYSlTu787QW10I2Xy8FhlL+ZFqoQqMZ51oTKUxbbpR89ftdZpqQ+
cZfZibUy79/TvQPOkWMonmnRT9uB9lFxn2AUhsn/tsQafZ/YvM4UEJGj2iVhk8Vz
A578iUMxcMTN7z466gQDc1VJD0Stk85uxCBwdrDfoC+DEuzqJaS2iiuy2QtPR4zG
08Xi8DuiT+W1En5G+P24ixpeThIy0et01wNjrBI8zu/Y7cUjJRZnMJCbxtSwbN3I
EbrKmrlM3I/RzRxNIoImbqmuSSA89X6hGXXUHl/+3xx488yWrqqHgtJJN9bAdjOB
D9pOBTA2QmihRaH/52hs8iWoh9d23Ojz9pkIVbwzCmkPEExXU2BKLhctaASawx16
Ayw/mW9qhjYDSDoLH9mLQkg9486ruHX8cT6Ksu64H4ndpZCLCWhr33iVFA3TBt6q
z8skrLnUcJmNLDQge0sWRp2oLlOpaM+/3vLu/4DQrei9nwfJaNACnab7SwNS4rnj
3VZ8Ve49f8yJgAp/9v15bISrxjAiR5lVlZMqsqmuafFCLBbkVvgurxeY6ZLHNYLg
h6X/rAzOY6+p5Xb6yq3tYLqMPiBM+pg3NjEdS1oXE0lRusgf66DhOHApaHOMVTtM
0umD/0nrcCM+MUICGu09/vWQ7cJVpQhfOkVhvcCdWh1QlpujZwnbIklPtzujrx2A
NuN9nzsBfGWl+W1LLo0NJ5buATwhhfrMWhHIGRXayGL5pYHyBr6yoY7uZJy1xlyA
ACNZsl0TmViAMIh22pKzzlvwgGFaQqxhFCjldfkGznN0PZxUnQWjAUK7baJIo6ai
ro/qvSLg2x/RktS+j2ppokXIJFOTnFlxiS6AbSqA9iu2AmG/bsPQ8T8KNZhJILv3
WFaRm8kVnAStki30ERI/9LTiG9fizJq0n6PX/MeJ/AcQFxN0GyOiUYuA/TAKklVp
18nBWOdsmK26fd72uTTp+CMY7BXw6QluzTWWJV4OLYGBt8nWyCEnAr7xv+iWIGBe
UWjY47XARhWoKr5/rHojfuvMFpgxsamwCa9AlllJd7ZgFkrN28663kxAA56DsDvd
ZPa/iIl9IXoeOAs2qPZXF1zS/c3j71dn+lK8Pr9Hfg7gl3igQT3Y2GXdAa1agF/v
TSwMCc65Gy2PhVC4Lrc6zAI7T372jjCrlCPOsxqeaHeGiDeS5lDd64MwRFO0HnkF
aDad90jYYiu6pPa/1RqbyG0JQ2UWzp6hcwZgLazhhXn3yyeumo5uRwumDdKwNgfg
5s01P0HEDPCTNd6cOq+cP4jAKon1Vsn3CBxCGe1dbtWN+JbHlhVPRucZ2jhcm+5E
t9TEu5QVQKvAlb6k2jZ3WKOlRvXgQ1WwUHK0fL0GbPBvuB2vdyACfl0rUVTA5nUv
nHqNhIx3DypnLlXsqZ1T/k/K4mI7Ecn6cwFWNWvjFkxXCliQxYVEgKq2fLnmTRNA
cbFL9VabzB5syZZ1yx0JLIjc3HmK+mWkXHhMAzxSVKvMZbXHMtTipTNkmBBwzG+V
9dnEyZ9FVjQiQZnF+zcsLi7jHvf2UwDDGsHp0rEpNt45liHhd2jaBzsEoAf0/N40
XCM5AuYsM7Xl/CFld9rS055BwXt4pZZ/2OjkLlfKM8PyTy9m/OPzMrrqVFS916k8
8EBudBaaJ0Hvxt25tvhBxEa8aIxoprS20Ret78J8WoGf6iQjZMInQsyG2LTWAcRk
LvENvZBgaUXAabXpIJJs0fbfAzauegGVWB6Htb20cCKAPe5nNdf79nkW3fr6Z7SC
i3D79XHJfg/G5+HgsXrROm0RvTym0Elk8dBXASpWc+p8P3wgJ22ZHwA36wAyEnro
T9AyXJxDroFcNel16rcYXXWdjbkuXJuXf8pu7JJnb7J1kRPro+Kc3xyLU3n3DA4+
gCPTk1JXoZ71zQd6zgUN4QdC28svdupXAe8LmZBVrO6Uu42kPuDV/nXPZVWa/66l
Sc4GsfofRhLWBRSIqou4FOZakW87uU8uIyYy8BggxfuRZssqovIkPfdND0l8xB6C
gk0Dv6OXPF2+lsLNGhrZbkDnmKJ/WwIoToleadwSNfljtWOYsJw19Dd9qrVz3emV
8n1aBJnKCyCeJsVC1Zd0/SrMgxVRQgvLDUwvZ3Pm008K4nQZGKDEY4KZiVVevdgo
kKhcBBN7z705otTEjn61HvBlTsNFpXtXagzFHbmrmX1zbZrl64Fba2BH1c6ZoblB
IinvDBKPDd0QaBEkjdkyFkIxVOy8D/86UCRA35L5OTr2/QRQJibXGRSljlkleanP
e4Eq7pD5Q1dRgxXKEuQGwanpTwgrAhiYha2u1Vf72DlKIfHgLvS9IG4AHorlYi0J
fBZxBwXGTnws7PMU/sXe/+X1bImTOgGy+QbK0/KnfGeujrRGJKQFqEl8L8fEmV/f
CF2XDZCA6A2XvMMwcXjZKsSQwuA55Ooy+/f7GAyO4m1qRbDqnZGUYXneLyV/8nM3
A5OWd5bbC4nO8QNHG6t3ClTHMESrKFjLB1wZnsXIZJskxE0L1KjAqRHwTdD20rtD
6L2UPuqyFVnC8BmQ3fIBoXgsUQcQFveWlN8FDRhpuPbVBl8zLPRfYLJpVpIYKl8c
+xu5gdITphnvG2DjroEZt8hspRoLFbCqA4ExtQlvqnEEQ2N1pzQp6STPiAl01l7k
7kzx1rXogDgpGydkoncivCKFU5wuBTl6fvqdSEXLIZu7xkLfHLoG8mSbQwRm2CUS
8jk/wIxQQoH11tLdhAEKQC7HilimcS2+UOLQpjgXPJj75YKkAE0uKv7GDuVeHMU7
jehrWB7JYVyvkc60Poi2zCf17ZOi9LlMHGSbmSzmqZ95QbnyLJ8Lu61NUTCDAEmH
zspp7SkXQhSrzNwhuMW7QNEDA5XKfqNh1ygeVW3KFk0gHyR5x51djQUeYn4AG+Jp
JLW3p3MgtwzgW0TS0FWFz3qW2+O5EkrIf/63NfrDM5WzBaN8KcqgQ51bJkqsxS5T
1TJ5msNP+tYdu1ueY2Kc5/22rBJbJ4BnybDxrQz2LYLxJqVQzW0XmfYQdRA7oriR
BN1SbOfMiWdFV46gIZIATwSfX3lSKntwxb7EvZSvdOK5Hpjw+ClWx2y1HM554hek
9MEhqWfcXN4a4jljjuBeaW13lGgFiTnG3c/GkxtMuMo2qwO/+rILoXvSRCfPWbQF
3C0c7QsbPUHSaSq3gLN+oYPQNRap4f0aT8k8UVJ5rGJhGtWD+J/fiEe3dOfwuvWH
wvyKA7Eoo5JIcQxILxBlU2iAtrc1eYXC1fe9DVu5LmeLm7bSLyUOZGGoNiTd3B56
0xNUBFSuFveOUlWJALyCGbPjP3Lh0aLeOm39lfNZ9ipwf9PgQO4Ssbh8O2QVzJb5
UkLf7YbJzsPE6syFXDNVf5NfYCI3eQLtLyFyTv9T+0iy9+Y4CxTYyz861CN7b99E
eA+laAAdQhJTDmeaN3Br8cnijeiUY533Pk+5r0FurXkGQvYizVvk2p8kM+Xo+KyS
WwsudzmKLKr8FkUaIsJGoV1lX9bIcZHhmYgDnIoVZnQCe17ikGMlxYjWOrEeFxrP
AQxu7kbyfxiBQVIZipFiuayVOAdhNfotRzyyfn+MFzrmNy3FQJuPFy6URQjAsdxQ
dGhn5Xo0V2prnElJp0Rtgm7YivC4S19I1RJJLYjNlFE8JwYzOtCj9GYaHnOgaCIM
M7C9wyeEnxWKhlbTrv39+2Yz0f1JhivCsEtIzzWSmUenCwFxZs9pnIB/0tRFa9ye
ibQ3kMkAc9FHIXQQVv/4cCGQuzrG9rmz/GiGkNqu+Ga0185sfSxHXPolWyv0mgpO
QQYB1Wl1Dgds2KeNf8ARc1lZ6BjJCWX+hc6Fv7rAGyW4p3JunQburlW8xMPsLf0E
jCh7If98c9u7YR5cChWFTJk/oxIg1Mo6dfpz7HQ1pItykqQFgc/E10O9+IIGAutZ
wjq4VWkaESUDoHvOpX2sO3KY3ULfx01unZ/tn3XebozPaRXtTbtsxX9C8juJGkNg
SRQ/WjJAXQLT1xa2RVQsWpB9iFdIUzGcUiJp5D/IkVwe4w3ImjbhJyrkyn4cslks
fzF9bSGi4BiIABlUgWIgoEpQ6CQnj5tDZ3/z1OEVLiJz23Sl9S09Eba7hTfw1dZz
EZ/vrsuHyLvkUczIVM0QW/Kc436P0BEBxdR3jBi67hSJn6lP6S2Nsrsy8XjTb20A
qo7y7g9Io9ocNDiB6feAWxxGXnfZcsli46NxrvhfAOaU5t/gKPr3Vqnvm8hbu/rn
ppfB7J4xPs9D4uuA8PJH4Kmyta5oYs0S2R7Ke14d5V8Q5tpA5rxs6OlktBG1FADt
KmE7CXS9u05uFsOcps1JyoClTyUlMH0pZsGSooIcaBqWRWYoDa8aO9hlzLRgqTq2
swOyPj98Laqfejz976JUegFMGNx1xR4LwMRQSFRdNzrei92ipk6MPFE0gRZxxE0o
MKACjQ0v2YC3EzHLEg3PvWc1plNH9wFDgi4QsW5BUINa6MshlGmpEYhcq6EwA3xQ
eqqJeNGNTNMmXT3v9Hun9FZbkaCTqxtt4A2Ze7g42yieRKiv10aNs8h31zA5jU3O
owEAq2vt+f51KC17hhSg3TdSSfkqnHxj8/3gy07ssGt0lhQ9uij9Mk0+Zcus7XTF
/c3a4/aIE4D1ImlYwodF8SwHgA3n9GZlfh881kyV4UzzcTShY6A6A588KuSXf38f
J9L1GFtdSlADqgBoCKK9q2wv+nwMpPxnf6zedpDc3gllXtiMYestIG9uE5gh1o37
TDEkE5dnM9KBxa1yBmvl/sNe5Ymz8TK/pS+PWBIvC0Ip6DiB7Ie5UeZPDjHcgS4e
TZMBMowiNqxKCoLHgnc+PTo04BYmePl5WngEC5FikjJazg/IPjESnWSbgwaiKUDj
WI3BK1D/WSIpTDvRF+XK8oqk3vU1qC8SywArtZQQOZcleGyMWeLue5RtWoFqecUd
vbv1SEXgkydVBQy1IbSoI1ORpkCkfw34OIQ7YIfS9ZmEfCke5hVrkHQILu7AcdSB
Oz+FOqzjKXKk7B320lO+Pl3YTiITehnl1E61uV3Sdyee4QUF3/mYfd70e9n8/InH
AaryiJeKDyHJyZIkmE9C4zgpaSvZER6aS8kLD+NCqHw5l12DvlKX08LWNgUDMIRE
rrWWMPo82DjUzo8sjuoPzawYyC67RxkBbF/d7qY/G7d95ESDfz9YJkYFPaWBZ7uQ
RrqBXEymHyrdyvUfmpVM7fdqEdPCrfCP3mgv6+JAi+8jfWzB/A4yLL+NSD++a6xA
hiN8LW6D3437bqlkFXDIN2HP3vguGhQO5W1g8M9JG4GCPH/ZqUxw05qPkPL37cgm
Bn4OYMpoArliq0t0aTdTGvTrO+rL+8zf2rxd6nlvyhQWw5y45dkOfwEGqQsqJZpK
KJrUWtSsZuBSXiVoHry3Tjwc40AFiDy+1RnJxzx+8AWGjvbvKd8oTumJn5GYu3P5
Rbq1J/89DBfjBZxZPonB9jpSSYyjO87dK8M/g69DDflnnggpbgOklqforjL00L0p
5LlnoBTzBRq8Z69UqQ8QeGlqZipim3WOK0BzQDjk1ikk/RcEVdLNA6OY5rvFYbRN
sk6YtkpulB/+D/NNxmx+IEYwEGEA9F9N0/WjBvZI6v9AXGyixb04keudrtpOs/kd
26GuHp4EIv4IhbcoSO9Pw2iUbOxI03CgjddecfMFp/Zgl0R0O7TdqRs9r6Sudf3U
LW7qCjAWtvnMZpwEis2TM3YImG+b+7DIpF9M6sayPWNQUF4MGfnB0FLXOBJ92hhZ
krsKB8yAFybJpLteFpR6u/v/e/Kthxrq6aSwDO+zjJxx4M/qTM1DM553+IKU1wIX
T+tFetNK1+B42ea5FE+1A6SFbmGdE4kakqJCfxiEP/b6c9Frp/Oklb0JUPVwArQM
iSs8HjU57ee4g84jTyeOgIRHMB/HzkCkVRiMPFPHUtju1C94Xvwv0aDQ5nh9/9lB
GWNMREoYBQSPP+iIfXe5z4qHwxK+RX4+2zLygDiB3VFuPaqSn54+nfAaTDW3//Eq
wUfSByatqqN3k/JuNlqOIIIwHlm6e+t4aW5WIphTiiXYbjbp9YduYXbqjAYABI4U
hBHIAUFE7PH+aHK6taiE93F9rLb9Wn4VQgJBF85vvLs0SuxjiY1Zvz/kg4PzIStE
B7Bu1MZB/UuWVDYdOsa/Yg5rX9pEN/kRf6jiqzE9pbqEKcB6Q5+OydriB6asLfm3
+VQDouAG7w7Ktxs4wOboT7Uuq/KWSlPu0oEjd0pPwg2tR379LHmyp06mU74JOs8a
EO/x43tR85Q3nC5qfcUyRtyZ+y5P9cRRBljy1Z0uH5MVHYsStgS2WZpSlDps8Ifp
0aGO+7urLOHEo1rKX/AEf3nl54A0JwB8UsoH+R2VAhtHvgGzJUvr0/MP/8M0iC9H
L2lkgZqYeO8B0lh8XkJi+LUyc8aGJI5AmiBZB0fqkcq94OZ5MqnMPm8ryYJ+eSWe
G4/bxrQxnn9kEoKLghaIchUo82TiBtg9RomABL9GG6u0pG0QQeebIbSv3wZJvmrv
e+D6A3DUf/wZfP2Z3eTDUMX/ODKbQck2x8KyEG6lsmTBl4tlYubc0/vm6/3Cd3df
+dH18RGbZU0Kqr1hyI0Nl1xcm/8FAGLwpikDu537itTdgC3hN2TYkpmKKoib0yeK
9VkDLbx87HBrIiO1X27FHjd4GuGUkgXiQq4yWjd5HdAvl43M9oUds8r3D9bEvuw8
m6gAcMDQLLEqfSyaAxluyKO+75LWsk5w/q1kCHdybnj5FwRk43g4NYcBFGvmGYYZ
AV9z3BWuxWnwDu0/ePjPsKMoGJG4fiYI96EdN7Pn/LIqSETVLip/9UcL9VO7FGTq
hnXHbFdx4P00FjaiHRDAOy89ZiGDOIzvTmSYP14sxcdjvOLYQmVKlUeU9K3tjH1q
oGfU5DAKAkn9/P+S3KWOikes/MIQkzM7FPo7wNgPdHib14sadoW0X0SKMcb8Yd5l
Xo3eZQCEpnfBoFsNo3IxGljulOvtSSZujKfch2C3/7Va//yoSZGP6NLnMHXUDru9
9rsHgKSruiEBGND/qCDcRThsAN9+uXmRQjujSjobOxJpoQERYEUduyxYFIml9K9z
6iyQ/p6NFW41nogwil4hy9MnRbj6ncVg9JA/V/FO0szQkB+mX/OdO81O1NJ7Rhwj
2/Nb/sAJ204hAh8IhrIBZIDeGAH840WDzA9YzMcYHY8xSS5kI0QMagzJk5DfDRGW
Gv6NdcM6PeVMdYjMnTKoe3dpgZgpozuVtxTQMxdQFok6hiO3m356em6NopShGZ9o
ngsBbKRc6qVUZQFUiTRrnpNblq6ZeOKC0vGrmZKWaSJmwPe/+U9laXWaSM2jvX5o
CNnPI+H+jRxN9phbptSZ87Nyx/RXP8YPnVM+knxwSTeG0SWAmkK/3Xuc6uAe1i7B
av3oqEu9FdGNixyRQSHe3zBlYehnHTqDVZglCPzq2Ao3LIayLLy7ji7zn8rfD0Pu
s4NN+pG0/sZH+mKo+zuQtmzqm9rkSXloTJkyKouZW9GhEJ5wmNiC7oVt73NkEqAD
I4KcaDxMbLWLbBzIgd2jzK6Zn3j8dY3F7DpJd66/aSW5tTSEaz79dvUgSTCv8eSG
5cQPv43RGXxOEIRYUZYvwsIwbklC5onesTckNIX6SFmHb1lrMWWSDmnfQ9G+6Pcd
zVdaIrrgw75acBiCVsT1nvH8ViuoqhNoxlsztxhjWCXzm2UJ7sNyjk2CqTgpvj+l
pwXyNV18j7+cvaH2pbebLtticpOM2GIXMnLUUzoAKQXHfQkX+n6rHADRWj5jHUuq
7pDB+v2VN2ipHKYiUQ013fzuiToVDW5Ym/3nr7hzSjMyFkSLHplpPa20ODGo9Qif
upq18D1njjoSochO1QKnpU2Fldpt3EiSLbNUsS0U4olU9KwBgdKohlLVQWKKgH4r
+fQReIjiXjOvXK9BmBYqPFBAilMvRYbunnDig0NbKi5CbjAdHXdmFNhFzUOH1Er9
0eeH6vsB3zTa7sJNJNCns6KKY5bryCMwK4iaU6xuLVWKJdtIODPvdIlto2guHZGV
SZX9OqwO4B1HbrjkZA9AQntr2CmYXfW5gZf+PJadw0tiQEZRoh1NfEZxzO7xKzvi
S8oAqXNzZKLyDNnTNUzP6VUnun7745Kw2+wpPv58THQScbfJ/s0GAdnrQOE3zg/y
cKuZaraXH1Oo+xsm97GVZBg63MvtUzWsw9sJXPs8ZteOs3FVuqMj8wX5Zrxm+xyc
5mBrMqA65xKFWHxIx+90Y4di0TJjfeQCBF3UYG0s5PcWq/s1k6U9Wzsk2pjsMl3E
6xjQIeEL2NJqgAx3Y1ML97Lwa3AQj56v25bRG1HiOCY+v8v1I2AWiYQGsuTcq+fU
FPStqsdiz2Rx0plAbhJllOuCs2loTucfKBDdvK+CMHkZ/Kok2/Oarm5LFomtUG08
1QMMsQ15eSZeoA4g+c1wBmNfEJsv96ruNozybhzHZDvfRRScla1rUFPRHWW9MwfX
SmUj0Miiq6Mt20gda/gpqouDZJjIIK05j6CeBv0usyhQpdve6NLVxJElSNiJksbE
1wvBo49Z2Vyl2jbf4qCdPtajeuum12r0g6roSjXUuRK1DsT3hhpIsKfklwgQDdTp
nDx4OL2WRREpNp0d/7mpnZwVr0xQBw7EIwJcooc5vJGf8y/Fq+PWOBq/Hh7XS6eH
hUIS+vXXZCMl2qD8CcBRBwbFAeQZkmz4HKKFwU/ubG5uoxoCUvWD16CYurvS0bhj
6uuHulFZhreNnjrnzxaKc5boFjcOqHotf+uT6j+NfWvUUD4HfmrjyTnkwEp3YFl5
VX1Ya1nOFLAUFZs+kQjqfFhtYT4GHN3xgh/zKw+J7ZOvD3JK8OqI4xGmrQ9zhETL
FX9HS0/8w4pRGRyDFZE87+ZVSxgfdORfGNqI46zjO+UwA4Zi9vKfKiLE+Jxwt0L7
HkK33/RceWhXgukOVEQMfh7m24dv3UiCoVMrazaUQahzrNul/0x/mzS5oS+d6/Sr
6nsQKs9e7Ldrwtnedwszj4toYah7LaZXycuqFb7rHpcJBtLlVnHVrJ2HtUfOvyWp
swu4KRrxEL76i3jsnp7WLBVaVMkqhn6EyIhx1dFFNwIHN+8FTXUJXk7cQ92chM5U
e49hlMEFprYNUdQK6l+YGWWeX8lr8eWzPRJOIcdOMYpkEjc/H1sl5vOiOQzLEZP6
JrKpXejb7EyqLYnBjpTD9u3puyeRsqCgAIvkA1bzj+wMWxoPOfOI02qX7G4+kLZp
lE3/alzfgqDe0t5xdnu5Q2Q0Xow1liQRQLl1/yK0ZdUHpLBciqpHclW2TL9WpEQy
ZYydpYshcETAEuEndv5nFhV9Vkut9qtd9cQ7WWUOUAmGJyZ5ogW//xZrg8p5DNMn
fj3pBMjoAJs9G/MxoXsjcOb6wDA/3o3HLfXr71CmBExJSWQvJ3oRoCl6HKTvdJ77
a8kOyJsG48VXrB9pkpb9z9dHsMptql7i9+DObjIXqlrxnCjBOhDaX/ezwi5QCDwt
FlggRLoFO9GbhBUCQd8VxwsAoDOwRQ2a4n29bqoLDwtU8NaR/SEGDvl3+bFWck/a
67ivQOCEVC7woVz4zojoB7iUyK4+xH4blOTqIQXOVjoPUSlOgOd1IaIG+wyKDtrT
Liyu9nhii1nQcbhwWQH14HzTTwKiPfiuYG1x0TTkoxzC7Rq6EEqUmgdcuBXZCTM9
zGLmwfWqhUNJ5hZHPOqdUI9RybLsASwArZN1+HlhkgghXKdGh/eqpPP2bPGC7zgh
z3twmA8vTRiq9bxhNb4AfnqSNB++GQBf5XZ8Fxn2qym755PWFt+jHZERYfoOeFJP
JmlOVdaZx9etKGXQK5dwEmbG06AQwfm3sn5qHWRDf2YwtlhHKTm4F6sFhN5kUKtn
G1PElHVHYZ1A0xwes44qkSwx1yNx1hyNoCbyvZlYNY/TmETdTSzgvg6CWP3dr2K6
1RygzQOEh74/MZUsIhgP4VX+0/8zt8y4lt05Mj9VJ6Kg2H3lDUOr+GT015tVd6iF
DI4/d27gN4vsX7/Jiat7eRIRQdCGC1rZ7iko+fPRQ0VR7efxHd5N2M6iWJVh5kjy
IswFl3yc2oh6WlICij8KzrgNyLVUN1tcDimQzZyraQp4nfQ0uP2/coFq6ner6QrI
gBatFHUjbzibwg1+aQWsn0eN2zXysw0efXI1z7KWEX0uQ+Yel9oTpgmrUfH7OoGT
usnt6aUepTMCEBFHhMFjgU7QL/tcDG2EFOzHv0Sia9aofnuXyiUx+Yojqhn+qLFo
SvjBZ+BzBmHWnEPV/zT+SypuPbF6BrYFQ2JGE8hUTqr3+ndBRsE0OR6ZEaXyPaAe
qereV1OHG7e4QXmM1C+a18Wy+CoxXZDEM+pq4c4dgWaMk1qwjpDAw7NKNtNpLmrc
aqpXf6O78VoTCaIoVY0jWWMMjxDweBZPv1UbB86BsBSlZrYV2RN0QdEB8vBSszke
qUNqps4kq0Cua66eAvI8TqO4DDkv5MQNMY1HdT02wjVnZEg+TpysPutFMocQA0ey
YVlOVW9tPCj1Zzxy6SuwOAtCjxDyNBd95svSGvvEb5YM2gtnRTEMTvW3UsxGp11z
U5gusfnvELx+z2rwckfRZNKHh2TCBeMP9ArXDMOAVfy6vWH8/A1dLYCZ86ShbHAr
n9rFAhnSYPEmqc53fso3xEbHVz91lhkFusudPTKyfUYwUcSXMJnN1CA6PdfrR0to
BlT+KGkFU5RVQp7LVcI2P8Gbrr5SW0CciLOo/1TWe4tZWD2aeqgJkiQ2vdlj+7h5
oFMA0sqyJX/uZPGU9ImYdemcxY64dRAI7mF9TVvJivFyPT5On6WvLmMzYk2IEvCz
E3LGv95WOlf7F7Oisdmx2jEGzQ5hbZngFCj08PnZU+GfcHxsAAYw6zcHD34HDChm
UhT5zLz5LZmMbyoZLdFImCfXEDZ5TO9jBKP8b0E/S7Qt+Jq4M63/qsnPnXNr2uPH
kp3pQj4USYGLSw9d5SZcPUg88Nl/5cUaguyo4cUcDZR1P54yxIOyB6yx/5ulNX8U
rFAP/OS36EgpqALIS0s7xKHVifoGxo3tUzch8/S01N8gXXIHMtwjhpHlf3GHRh8n
kZgMIKfDrCDOxWvFynmglclQZDv68l1F2YE0mqVmMjrX76jP5xpo42uF6XkGDJyv
Gg5Qfz4MDwzeMS03CqAO+7ww/QGTbImovceXjCwIMHu4Efz1W0x0iKIDBP7shY/x
W+9h668tLRTKvAcdlMJAaXXzFZrtfZGMovnUlMJjtN0flkGgosdeQjE3tEmlv4pg
aHjZWwtpOYovHwvQxn7IWNGiKEJ1p+Vi+tLebY0PrDSHhkmH8LAU2TRH4OyFngtx
+gmfX14TxSAR6p0+hCEpf5DmP96OBBltPR2CZhuV326T+NQQviqYLyua5TZ6VnRa
OU9Ctxqr7g2+L9hiKjXl1PWS/d8AQ2ntSsrGC1i4hrcjbVdMo+yWKyRA91Zu3yV5
TbWsq8Cf4Nm/hg5szcFUrHoWv8uW7IfX4W8rrparrXxbn+GAvaxlv3PiLzFkZlnq
gq30l0d7E/8bkPFDZHTN7ivrGGVGj9wSYzNLHweEgU9GZRyKhB3sKLRS/cT7Vd0J
zW0lMSUZigE+Dx0e1lAUMh6lxfUUnKsFDSEQYNaq3bfTVtje6/ssKfKx2iednd64
dmm7A4/EDvYHgpype/JHFWAZ3Ui1AJUnR2QT4pqe5pDFpGLTCktnhvovRkCLgA+m
H2PEtEmOnEUAjK+bJMKwBgAKFmV307l+G0T6OsvIbTbi23w7xpbmFIZGQPBMh8yG
LFSJX2LuO0d50kuQg/QrM7CXB72yBPGn07uxv8UUqQgqTB3BQSO0x9OJUxIE9sK4
I2QAiRphy/mjSVGUdY57ZgJ5/u4YXBuyuGAv70cGBJT6lBgiGwkC3TY+ZwYnEyOR
FFef5rJd5waO6w4bkNQuSliftt7ekR5Mf3xTQ40xu85RHbm0/GgEoEw+R81vxosJ
TvxIcTJPSmwxMFXMUa+0VvxcxFx+Znkx1bYgUF0cmLWV+m9NSpqwfFEUZd4EBr9N
hUNjT8zo5/WSM+Gppp9rweAIdHRuZ+YLBMkgfLSvtebgmUwfP0iw4cY+AySzbhvj
95N9sHOPXziH3cJQ6JyhJpx+E799HoC0EAdZQmt4ciJqT66q5U7GAOT8wgD/wX3F
ErIAY64gXK/WxOfAnHIwm4wevr5B1NZMw/T6PRYB6MfewbQyUcRrjV/aLSlRnPv6
12k5hQ4fBNwmw3UoS9kCDC6YKHo36s11/pqy7l7umD01ZVp3OfHJhPaLxIauMDNq
17/WCrjQ8+LP+3mokP3O7PpOo0iecd8HJ/5g9e0Z3lnARFwVjSfmCXKXQkIbm+o4
xYE9mRW51A6Gpl/Y6eeiqZsxDQCkSt/Ble2mhuNAVec7BH3Pn95Hcy9IcyarcFAm
GrxCbAsI6f7rbcbqkmB3st7C5cCePggr0yseRYOFsTKNHtngdgyGnvnpBGUrNzFw
rLLGXrOedGVuljVVYiPkR8kCNSMVq6G0NoTb/U72AWFFX/5ZD63YvPc4K/SYNF4j
FJFCb/hvJVrDrWitFTJY7ulpahi6YQEZJB4JwY20CWr7BsIGaW5Om/i5UqvdRRln
v3rrBqoim+UiZjHV0trkqhhqFWsp1Bi8rdPW+1VKqV8l6A5FMXmr+zDSHQHIoEGn
vP0wgMARpxp6IhXA6qxkVLvXJcsYKcr4mIjp/RlgnfTuJG7GdikYUHjNzfp/f8n+
6VYV3PO1yVyR1yhroKpYd6k/6bGGE4QArcMR7bjxSXYx7NvLV8alqMHJrg7oQhNv
GGdZuTYIx5trM2DUNv7M7HOwh0RK69A8RzOAdHHVa8IJXp9LIDzJ9YmWfUTa8tvN
8TXcmsn2eQpLbxF7PDJrgWjAd3qaKQAn8vp7rbisizJk7XsdNeJFLHQO2AZsX/XG
z6a0gtcGyYsHZ2ITBboRfNBnxKh0wEsX3GNWNOTYV7MXL9upkmR2DOE6Ku9vRhhP
JJyOg/XgAulhKWwkfFLqQm8He5RK4n0a4xACR5KbDNrsSviq1R92+iWRgb06HsFp
9r2cFiC3fQR0vO25dhrVQo2NeEnt2SCAeB3c7HmOkfG7fRDfp6ZfZKwLLreiEmC8
ptLian8jvklzefu+MvfjwfmzGlANqa47hwirJfl8w+TRV96Hh7/GNL6diXyGD4pg
AerDkemtwylImW0N0sgmaSfczWxdtkB7CxSvBvsaENL9twdeesAMzXzUEI92Mqd4
5msQV3McX7IoK3vl8LXk/LyZ5XmykJPAo/10wYh8066lur7WfludLE81is3QsurS
T43lAT/ymeSbJ/z0S4H3NpBEpEpIUVoiJjIGqpCZlGCwhK/iX/C55iVoKNOKnJ2k
dxx9aY/mDe12mwhgw7ulab0fBE/DkkvrVc57JHsKIEEq7CZieV08w1kJ/5A4n0nt
QPhT3E0tKlMzNP9kkGKosM096QVvvAL2c7UM+Qz66+f4GfoUtG1u/NjyeQA18ZDm
I06sOAIlOpUOyH3NPwl9VYtuk/NdeEVbQx4e8BlFmFnO0EHVfuRl1WbY2fzoQkGY
mGy1iW1WEvS/MA0AuT8HrO8h/6BZd+2uTEPBnUIBXO71Xah2GlF5R+LYaGgO6w+6
Tebc95BBy2f1bf6IQXOPMhkn3WePX1ranlFcO+W4zsjBS8jvbnZqdIbozfu5HhCX
4zc3mIRAgA9+/Ulov+Biq65o1iWRUPNGnkjIrnQCalBin4sExPKpIvpJXzXQs0jc
zCIjl1Eob9tH0hYqyKq9evg7XgFeLEW7tMfoj6GzqzzlNY8kVn8zCEUDUlFCw6yR
zy7ENMKJ2mGiGSSyiZwByfqDDGGRX7a9tCQeJL2Gmgdg5WNLLh6qaWAS7sreHWAr
t4BJgwtcKI4eG6aSAseXP7ui4mvY+huF5/fWFb46y/mtBk2iMG2/uAw8sz08P8Rq
K/66iKPLe8DoSEYMaxlp0u09VBStDEL5c6E9oWtbyxLb0DZ8y6IngikqkJN8rBYi
9pr+w33/xV2KHQ4PuRL+kejDOz1XZ923PN/ZTGVuVhv6PULzQBIwwzYUKa/CBOSz
vHlbuCBRmhtEAKB1C7yITnRnve3zM+VkEXWMpLOYLZOoIhJqrqUd09RcWnqzWjdL
tN8HJraDYaNb5Crq0HXqfHKBTQ0NJx38/yL6mlFnIqvXEAVn+p1RKSkyzGtd/B+H
OJRq+AwU7+XShbDaxZRXNAFJ8Yn+pPXCTqXqLzs0TJwqjMyarl+JdxA8DiNYMhds
mJ64bx0YGdQqXDfeYI3zmOQa+PvjSHO/TJ8RubSPjyQn88xdngRLBUr9DW+Kh4Bc
sasdrX2N/Wv7XCZwK4wTKB7bv0S6FoKwbjYRBRKxof+/VDPk5bViZrvvyw6nSNXE
tzCguEbHr4LI4yifQRQAVERSh8dbpbWaH37Ptp/cXD9//7c6zhEqf8wDJtoTuMkR
Prp8JEHgDmS+DZC1lW5jbmcZlMnqECgk7HHphgN1IkGvhwCBn9QLgYICAaue2iW4
fq91n1ChRWPgbwplJrlaVpwn8+uNM7tDWuXZX3mCFijyu4RWEV7zxx6IcxFaDhT9
U+HmWRgQPzKX2LQ0VqoUkVZXUu749MYd7wkeWcS9ZouK8IGNRpr01+BSmcMpCkIc
jqGH99bxJOsxxmgWVNt+MWkiMTGLnpEaRfXB0LKiE4VOLb2o7BLSSuEk9BEp2rfr
PvWwj+/SlhS1sUPUjbkTPqxiI31HZUQZ7mrpuliu3TaiTg0tPFcu9FaMcr95sRl9
8eHjBvP7d86vzu9w18UDY44Qu/EeEqwBWI2RQQgR6GZYartwtLlKfe4hA6lZKb8z
TrckQuPhC3y8pqRzql0fGQf0v9MXx27++HYgyagYD9vIzOGCDHTOPCV5pp8jEGdL
ep5GYwOEAwH7tK77POdkp+rIirfc3G4ZiZoeeuK12yPg9zIsgIuPr5Md3A4+q8ok
Mh2MD/ICkSZfI5tMXu6ydCj184bwnF2pl6Lqv90xBsmsnZCQFzHyOKP2trIkfwzM
zFIMI1U8ZfeW+oqYBsKOie7KgLmhZl9bWZPcLZsFLE31mBBbERTO+WEKBwEiLX5C
LkcgIZ0LtAGvQJnZsjwtfAYrNy/K06FW5dzcsrcB1mM0UJYn1t1TRw+fQu4J3eav
RR/ruwO+ezH/Fn8wDGPMD2D++NMjA4do4ASgVQxcEaBSyVyUAogfX40yHRUsw5Lq
WUH0cpGPF6lt4tJsN3vZSQYXeKtkFVhbqX8vP+NWmC9HsFypJzf9hngwojC166nC
ZK0CbjrzEeXEqED+0DJfNiUDuQXqiEyJqJI9RX9N2lUBeqesBXau6OnB5Vo+SolX
L2fQT4GV+02z0Qc0rTIuzAjzbXfbtz3EIpg8d8KVulSBKw3sQ+pXjQf4XOdO8Pzd
Cy4bK8NPEpboh4xZaBtxTu1VaFwgPiw6k667ZRD1L5cONg89NBTGhtc3vH6si2kQ
RNnHsyQIxDtYm+g5DEmJ5FPjW4/7cj52ZAxhJtKAPdsF0DtLR+eDPXzhB6pECh7e
5jWr6MNBfScbj2TzZccqzpjZqSMtM9VPq7YEdiDkqg/bYssIiJoseRWDCAk8tK/Q
pbCnr+8udLy5EY+G5PpM+l2sdPOKOO40o1BdjDpWPouRtJLWP3aG89MWkHpVX2V9
eLTPV1Ku9ua27LtOq+6anbyloG4lABJBdzF/Wx1HjuU04OhEri25mlt2DwqkpFzX
RM4fHBbGQlg1Yx0LQkkev0SqGTTgxQBdAHy8inqHz8HLSeC8FsK0ZHJ+E8axkCyZ
CSmFWTQX70iPn34GMGJbGydtKFhcm1SZc0zBCEbC1viLnY3tQ7bpSfxM9MdPUssj
r716RCN9wP0xzBk7sX/UbdaPs0VmWMKARl3olGcdIYRLD49ZRKOnG81czNoyhHrk
5tDw1AhJHYzuZcvS1UTUZtBO37pSiR+w1WrhPdDGSA3dgBWgRQyqQt9j/85a/FCM
dP2XY+2Zhl2DKIGCHbRqWfVF0q/8087iMp2WxajL3/YqHsVhrMqYEPDZ9wuawP2b
bzBaN6e+aejH9yG1XN+HOJUKrnLW5YXQDhxaoJmTMViDRTdh64J/fibW4g1h7Pq0
lMqn4R0/I26gXDvYLFycgRN/KLCkDZHTEkipPGadRLrbWa+ZYMl50t5Mm9ZOoHV+
iAiCjBXipthBelAPWgNGgA9oPUMwfhfHuHDZOD8n8HUtUPUK3lT4cuTfu1A9WQWX
BL/vqsU/R72/vbb7ig99sO6tJml9n4dV6bJl/IRRpRx3/ZcBH0rh/Ypna5jMZSeS
ae3YBh7zuJnsCqCa5aWsHpICyX43bNXMD/TfPrXKsFUW8wLj43cgjLlB7Ci77VOO
/URY8AIpYGdtXYGsXsGw93rVwcaHBwsv+FWYU2ku64o9FWj/kWDhkInBn7giG5sF
hZzsB2uHnOjU/KuApDq+UpBbNTMwXXgEakCQBiCSLI3dAzvAfquDJUHEdYIiPZaQ
MWndfs34NmzqOzAJBhI8lxkukAJBsDvWf6lOVoy/zchrRhNPLAwU4VlzzyQWH88R
qCQAjN7UlNtnmTLJHQq7HmrpDDSqhB9h/4FoJM1yW9Pb/YVulPqp8QhkKop0coNu
cn2sZBzobmTD2sLYAfAB4+yz4PymO8GYGLoz9gkX8pLQRiClT4uzC1Xb4eaW+PDy
vi7IYC6qDAF9CSZZ9rKgVhhogRzKpyzB0ftGatJpinlTp3jVL/hq+c2EG/nH1KqU
0/ZLaT2swJQ7At8tE8rN0kRmHoDpiytCp5CGz3cZdV0GN2sQR6Nc8yTeuvfPM8/w
bbcINPjFa++99TvNgTPXCAgdYvRBMY+ntXtQZRIv8lrJesaTrPOQu/R5slzacBJx
PU0mAlSO9v2y7fDimvnrW56eWhQPw6A/ulFBZBZzOcjpjJQQytSN+ibT/zalS5YI
+CuzUZOZIvdFbrKtgpTbMs3+mDuwKk1sY5Oxc8qj1dwiWAbKEIu8ikoauEXEY5hr
GmZ/eRahF3hHnrB3fGn7PRHoMWEWWN/IExz+fquCDwkPgtK+W7VwAJtmBcUEJKvq
0OIISuYG7Q+434Zts9+cZgJAFmLcg6itwIAGtboH1GGOydUyU0vVfmTJ6R39CEim
GU8FyWEluGZQUvqRMn7r8C0Css4R/gK/Aumez7d5LdjqkvhbyAZIrzV9bRorK6nR
wkqmJ2RWpO5lZ+Cw51mlVD+fqgddKzbgq/tfoBNHvQQWH3FH4Ghwrg3wlRwEz0uK
xRYQC/A6Z5oRwunSe+nvce6hhZWCDSJSGj9/K+i2AdC1O1Yk8DVLM6Dw9TLw8GSS
QycItrrtYT+lAHt63xU+WTKqAO3a3M/YAwa+BAySyFrM51T+y7XZznNip2wCjp0B
NU9r70htpXIoxO5obyHVFlfhE8MOoj1DEMlMKq/9BnYU9rZq/IXFJz2/S2gSBBCg
oVYnBYE+aKwwyidnDsbeZI4EUTtgjRcdhe5eQL2bAmJ7NKwEsbtEbHml736rCsSY
iGb4n8xlq6s78i5exHdO7K5ucw5YDdLW8Sz6SrZ2WEbvdXglD29cnsJGdygM4teT
NyIRmUQSd6qGo9nnC76vUhB+5aaotyWeY2QqmzzXR+D9jJsAYXR6pq06LrF6HA//
TnkF3uWugYUfggyHsZv9uNupk4M55Lyz3NtNBpdDhPQ0SDT4/GbpL1lUkTJCtsj4
gJbhtHhSo0hbIZ/f7VmjXcvabX2Y3MkmiglKx7pJ5ei/zH3BZoWmD4pYrSrle3hs
9LRGuXmosr17dmqe9PPWRzCpUWkt9byDQOTMQTU/0dQfE1khN2GzvngdslqXcoAP
x7xopGB8K9RB3I55EJIUmwdHYQhCLui/5CD24/BiqanemPoym6VUbz1bTWf1eF3d
CGoi2rpGVLxDFDLpRpYVABXKIRroeljevhqlYApPERkwBbNxM4rH2my7nnQBXp/N
xHdGzJTihXYz2zclNtELFdv3RLeKfz1Iog73+BaXz76tD7BFo3pY5vX+r/4gVJFV
3DxjwoApJyzMD7X0pl3I4w4cqfAFu1+2gPc4+1qxjRR+9S8Gihh2nidaSywvKxGq
qS8xVZpawAIFrccgLhQNhV2kGrV8MJn4N/vV27ercIWx/X8euiVZtVHQLDK39rg/
QbW86eOsKGObCWordX+SJQAg8JXrOaE4iilWtPiXm5yuRQ7XRxe9PABAppjMMFnO
BnY2N2+S/t11BJOOx7tsMJUAPIoPZJyqiKwjI3rqJFzua1zyGzT2nRlHtuImoJiK
Dv9gSEs5j1J1uRz4Thl5chHX0SakORTiNX9FjUr4euN4Hd7/9PVzoUtN+cQg9gDg
YfmPz7T4veNnFUhALoVL2yjaplXySZU+6zx/68hNX+AII465/4c9g2jjfoP1NYZA
f/oKSE4GLeHzBS9sREheAStwwWGLJyLY/ZBKNgcyTUctxoTa/OTfO4Xnon96lNxk
sMOfkixmN8D3JGW38Cou2rLCGFUAPetmEgSBXwDzIPrPOJr+skcJg73nmBUdnwfy
njuvm5ZvZBOQeagU/xv0nekFBYVoXp7z7iADnYYkmM5Hcsuq1U8F/uF6QE944NFt
+DvznggBMJuR4olut42yvt23DG41mfGH5cZF4Tu/weGPWqOnCEtG8AkR5qO5T+dX
onBLDjPxsBHb3YyCkgWqADSqrg/vEtB7NZFy8AFz4f3QHF68Qtx7aGPFpNcVS4yW
BUqMxW0/K9DEe4+ip0vc0WjpMCfitRGhzsQL6CUAuYiFqbic3syGOeNNehwD7gkH
NZ12wgRBaVe6ZWhH6QO8NKjeyibDq20RmZs/CG3qzLz3EAVRYoQUSt4UYnhVNAA3
dC5syOUgH2QpABTriTgul7tISBPAbMssauAposSsrD5ngEG9o7YkZqpiyyuJOGd/
l5UAXynA2R7DHd2zOv8GlVFuAGzoKRC9NJ2Ph1NkDByW5CivnXU78LTybabhX69Z
jPLUHJ1h7iGGyO1Q6PlzxBv+daCWSlRRwLHG4XJ2n2Svwa/CKSHr7qonUb9dn1iq
tehHaCv7oX9CZUt8c7w9+v3hfobAj5/DcBydGolMnFgK2ZmKhJ/pEetejKO8Wp9h
TRlDE0jri/HAKAIbf8+SCUHurH1vhPknvW+L354GGuAfrGhqq/Hw9s3nLQeO9j/1
4jrKwj06uHH4pQHRVhM3kzrZuMKPKsHYraEWuDshOvgyozGV3hGR4JPEl3xqbavZ
BSRU74oyOHCkQZW8cBvXJt7+rlZKjXgVBg59PnR54wh9UVfGzF9rW0k2b0mh0F+7
uHG+WwfPuHwwRDgal8hmzUkY4MP+LPiINgSQ6Gv7vd38t4ihkPL+cvc2ru+w5+jH
X6uM4oym9mfqbatU+e6ynsqnfY1tqJ6fzqxZoeeNGsSzFsYOGgCiFZ8rhp9+x9U5
ea3gaQTb0HblZDG8UT1nmxEOjHW325ki2INJ6jWVepkcq7PKJSUhovE25h+UH4w0
zaojT39LIGC8S2UPgO9uUM3+g8LF5f94ihUhmp4s4DKnQKBgkguRE9dTMhlfTfQV
hMS+NkifJ0AZXXWax4a2wVLQXAPKmFHFCGMr/WWov9GK/5wZHlEFoCNLAqLdbxJ5
f6zkuoje6o1UpDc6VFdgpu7HBSNN82U+LnxBx/wzKLWYK3NRl9d3dQVGq8I5fYJ9
op6VvDBa7LbExbdR8sgZ4G63NxW5b9Vyzz/0AlEGwSgyv9rSfCydA9XKkMKephXU
3ppQUrHE0Pj7155XO5QlpU6dDzefdYjZr6XKcSy123rqCI1qvO8IjjfYYgx1RfAU
dhihjKbyY5nN1C57H6xvtPv0j9lMhi7dPXzf5fvc/XnMVNxSWf5u/2E9gVuqNhJN
KVibCs4wdAOvKiasMqTrlgPm7sfrI7YCwfsUbx8g292FhTMHTWd1JwtHAWNuBQu9
FZU7NBvAT7ITtNGE+3NaJbY0yVIc9XGEBy7bHdg4sE9Jx7YWwrda4+1WUwF6qdH1
eW1CvMUc/9LQJ2Z5GsW/pb5mw2bvuKd5wXweBXxNyiKR9pivfPqX1nRh+MYF9243
GaN0bYKDlA1oqPIEZnRkwluqd/gNH/Tcdgz2NiLyQtvEEPXAvsDQmNcckciVa1FD
iOnAk/FviDa4jlf/KnY6/siM1vkkplln5mQ5R1u2K0/8K3kYXrxFC549l6a+x0TG
AyKmfxLqIZqJtYWBAwYgq7RpngnDjaouId4FV9S2j+RkGXnwu9lzBxUDo6bKWd/K
8GIakGjEH0VIKUrgRy07osr1hIQVb1GROhBNUQ8byqNDLTH4T1ES0rhJmLtnXgE5
nxx/viE6bEwrsEMdMD89RmYTrI5Ac9rr0fMe8oOniiEZi5PwxIevPQCm1zBWvUJV
KZxw6t9ic70gaGuBGEjrAl9OLPEEYbmhffOrRRno4q1IO4+nrUM969a5bImvJaf3
RY035yu+9enbmwyTaIcONC/Lt/f0Sr4Na6gCMPSgxfXLfqnC+NnIVHkv7okK3Qoo
YY1JegQCYHvvUGXAmE6ROV8q99gEQUJrXS8RSwBESjLuLGYIFMZ4NQtBhq/sDssF
EEHyd7FIo8wPuyE4Glyvz6rPLgSUeQTQ9ezgUN5A7ORzCQdKeWPl5ZGcX26OZnXQ
adnHkUGjljrOOjX1Uw0GweUwpH7ey3MPl0GFE3CT6Iz/+IdIIllLeVWvvWr4R2aE
qKrXz5i785oC3NJK6d3L3Aom4cdYg7ZZcVNoykdsLFTuIM+PDE/zncln1+VWQHRA
tuDZeKYQKQEdin/h903tPEm7orOmETSR3Y8Gt54qFqp1eowY7RA/F0TvX56FuJ7e
wlhugYHw0RmTMMRCXEtBK5YrLP1rEzun/hgZq2sT+kfYfwAMR+xOhDkkNAZ9RlFN
iPSs7qgtf1yBiKmp2F8MS2MvzCH7ac1r/42y/xUpU8L3/5lSdsQmZC4K+/8Z6b2k
OssTn9uU6pN3vaKvn4nDkdD58HdFekckGL6H8b8Vb+x+m/xvyXOs7pDNuH0vyXUZ
XLq0Wlmm+BsRwHlPwZEHTL6A4jbCi8M91MlpkpfQPbFTRW9393jVZ0AbsKSYGuz4
xVD1HptS7XSWmSYmv4GDPibXp36QvpJAaBww1tgvyumM50NH0VdCTlB5Vs/QUTj7
XxBari2BgzNBL93x7yWRFk4599tHlTxg/9C7Amf7XrafIaEchEovy53KJ2laSfSJ
lBcAz7rGoQc0CaQiLyqdJlMyq1yrp2ZyFJd0eLVY9bszbV0JIlPKd9k4bADTAaUu
+7Ap/UDRp4S/+Z13IqUUrgrThEXM9TEUORxbYd9k5Pn6N3OifSO0mVos0CxdqNFo
EjR0C4lHCRAzqT2ECNkAiDuptbv1zQBhsdKPP6hJO+au9NHnQv6n4uTurwo5AHoT
ZRGCH27aRPQmHAkyrwsgWfgiiiCREI4nNcf8kTEWU2h+mKklgGdoX8SubSGQRrpg
6kN6fsELPupy991FOnK/Io0r86pLQyLXwIpfipAvDPKAiyPFGTGlMV6BchzeHqcx
kPyAZpzPuIsgzUai2BHDhN57mZW9DFkMs+2Kf/37YF9luViKWu3EB8qkTsFEjGCd
iRFONLFEbaHpfjyiJ5WlYpcgkG083gDvZYjVrXr8/0ybM5hrTzmItsrO02aXYUam
86QO4gRiqtgmghc3PGcPE0lZIGinq1Tu5zCPyFppEvlWJ/aJnDpOekiQO3MF1PPq
FDI4XRH7dCC6rYUu9P2DOZeH6voQbydlThtVIottyfJBUOWIjeUb2X42zPHVVwQ+
KpSep06da6N4c/P+GFmFDzoTTQXcty28gVCw7M4ksBRBnBlIQwUWCWjZVkRIYPym
MxSlD4twPY17GCnuEt/eLNKKgHhTaL/JCec1nP5eqYH57T2cmMPa5Qtza0geqwqz
8abSvx3M3pFIiZj4qan2hJXhN7WROVYL+1Sh8ZiWEv+XvB9I9ug9U0I9vnK5FC6K
v7FRCo2EOhUUqo3H8uIST2cAndRM+fU48FlsTujDIgZSmrHWYmKsjlbdHjeB43d4
+JBbx4QoMsRXXs8c/9C3f/N+Xv1h2C4x3pgWfHTnadaf60N65JsmCMjyKzTZoVbN
/deQdFTKKgX0o25Ey24Wui0FfP7yfCel6mxW03OBnHPQfF58eu759JMB+hGE8NLV
cOSavNclp4j3exj7EtV0ShKqWIxGY23r9a59IlaiHcDDHsp9Zr1oFmUopEjMgt5U
oJ13JhvxHFKXpVyQJbirAGUbIfSaIhxJqoDR3POH4JoI0tFVJ8lW45aDx/tLE8KP
ygyE60c8seSn+jvA7ud1o39sSrZJ3CG9CKY336CHC6vb4xdjdRaUxwd8H0SQAEdN
SN620Ckox7iYE34JE0m49Oe5NBafzzkYDsmg0G8LIo4n3NhSkfE8v0pRkYsgIYOY
7JWJl/ckqW1eS6DCAjJ4RK1fTbk2taqQFx0XXdn5KEAfgsbDInpcgE2MW2dqWSb6
IGjHiMZ5Irj10oYB8fkOhdzDrGF2hPzc8MahJPjV60QveIcjNDXuuAcegia0RJ6Z
oyulji06/RFTBzAl0MFxsM6httqu9K92M1e41a0iA+zYLScAjVq6bkf2oaNI5ust
gSdrR6r75eSFK1uBjcp2n+5RRRjblgEwbrXWUr46h8Fk0QIt0Tr2EUUCa+FUszgQ
ld4sZcnHcskewLsg6oDNwg59gBaw0b6zYKtEV/h2PnahbUZAbWZIpfLcHTve+CFS
Z2xUqEyQPAGacu6n/ypW8ZKYIBBEvWijo5eoxbSRGlqqm/gvW1lePVl/NoP5rxam
OQBaZUTItC7Rp3xB2xIcODES2py3YvqTDrUT4Z+6wCFWe2Mc3M2F7sp0YscKBLvr
1sQSol3TBI+gjjW8FYGSz8aJgyH0wS8buHRMibRxgbXHmWaw86lcRyNrzVOGpJzZ
fVye0omrDKZtvbuzDHFx9SAGavo0Tt35sGiOp4zl7bxwjRVcNmIo8hmixkQR806s
FwWrEoYDTOB1e59J8pfVSkF7CywGOZm7TLhvH5CH99HYoEATg4xw6JOU8Edvw9+e
rRxnQrVyZpwTrIIosBIHpjZ5hfzRANwTepGauOZEvgXYWjPa2QK/IdPg+H4+Kw3x
4LZUNiJSSVnu6Ejt8criPHxeTBgk3Whekx0TGwx83t88wgzOYePotInxqhei1XHx
s+I8T+aKbJETMgXj8BzOVQlDm3YWTQo5xOMlYoTsIFXhPH/uWxxPWEZI2gle+DBC
KIk+48Q09b1WOsiJYMcxcShsibhPg5y0FzPElVHPLFi8zwAkcu9UQIDY++Emidyd
vRvfpgnM9nePqqvX3MNMm5MKSIfxZEKCLoOLxD6OnfnTVqR4QXAhjdf0w7se4vrr
0F1i3VpuYNv6Qj0JtpP2LAco7Moce6FwY9B5LaNraQ0iX8BAvv/PIFcmv2+Nygcw
GwTQI+WrBYNtIxA2SQlyRDKFBBiSskG90+RzMRMdzNzfFj0XZzVGHabC0lMUR0xC
kdo59km26onIgEufLxhN5lFT4ymqprpsmgZh2CJMLZFOGKKPp3O+r8M1wEN4vMLq
ggjT51u5RC2nutGHDJfSVcUzkmtFlJmlWGCJf4eOc3Xmqt3300h6n4iyEpZvguuB
kOLXZ0R577NM/grJOvrfkeSVwflCEvMZrOK35RaLuzMs4NleiqJ6stFtAJbU3cuX
Mt88DlwkZeT/hqui76Dx8hU+nqQ5wARpHirb0WUgiIU0Em74vuS8Lnn1oR0dEA1q
kYlxApwJ5JBpdfS2S7B+1dki02mUlmmzxEJcZb4vfmAJNLtFVAO+qfnhFlRkBCHY
ECTP3Us+yHbbz5z7+Q0zv61sIIQQ0gyOvBvBFJ49mEuLteNYljfQ9xaZ3OWPuf1O
LmVFxKSkNLPkYFahiwbr4u+icA5CWOqRFlLoQue5lvXWl+lx9106A/nkUOpKTwXC
GgfTB86tnJUq4Rbf2/jvEvvZRNverDguu8/VUpDSGPj21LCVqQfo6JFl15AuAFsw
zBeNSd6Fq2uK4lLlyflTPI8MiLoFNLcLgnWNGaggIkTRQhnFmgiG9pKOFroTKQF3
WRNWETK78ypWkpUMau69Z1pScGM/8NfZ20BBdr3Tocra2VJwJZuj44pImrV/zpGK
tJDLPBjTQFYMiLrUI+zNFKvuo2rDNuv+jsnzIOWccrakyuDi0sF1qmfSv4KewG0R
ZD9fIOfLU5oQYOvJZfbKVrXR1pXufTPyO/8gWMiR4YFd8F5psAonLv2D6xM0Y/Sj
TdDwLSeeSPmNr3/M3acRZCtVuYKU8QpHinJhgPYrJLfXcoksqGScwHwZOfedXrr4
2QhHq7mxuVar9rflBz12CazallzqfZquj7tS5kOy4GGyriJi1YzNkM2cVc8Ns7Jo
MQnjC0flr/op/bvSFoR03ey0gz3oZdEaD4TJ8Kd6SlaskorfllQlvAvDMd8R8Mww
2mVNVgOll/JrSrm8Ypbj70vmMBryKgTRntreOGEZglUgMzD2nFd+LTTl0gSuWFuB
cqus/8AcNkULSxVdT71ZX6QEt0MTZ4EwC/VGCUaQqNJ5GrcmFib5vZiQ7XtIlvjh
1XJ7yH5XxjExFIfp0P0sSREVYYMIiB3fSrr1r56kh2crqToOvRak2Pp+ZIqakQqZ
z1yqn8m7vUWuX1ZSR+awNYTJm7tHLdrv+Tdd5MMotx/vp23j1w6LlvBba89UlyOJ
zyUs/XizGs7Hlm8R4sGQxZkVpJ/3ev+TsOLepQLgWOQoE1IXKN18t1+OME4C4Uu3
9lPWKvBSk7QH8vHBtvMO3IMO6gZTRrUSb8XMEiHAiaihTTX7kh5UHktPcLxBziPA
mwftDYuO1Q/eAz3OzQ2xz/HkVvcT8SCAiLacOX1uSgDNmcujRD6OfQfKNPwvdxOt
MqtRhcjgBucPAHzmygHcP1f8l/i4eLC4+SfZ790e3rR8GEuYQCtOoElPerhHozZ/
pVHq4fZXlTNFRL7i/+/s7TFLPxie2ZrzKxnGkZlUAo8lBHIJ6F+RoigQndRix8f1
u2VSUCiuwXT5CJoJPNO9Vy91aAlMvx6oGF9CRlsDKvDWrP0sNF9LpdZZPK+16xfk
aHCg/QR4AdKg143dIs9MP0EeP1zCQZFprRfPyzJJyCK3x53z5+TFxXabZD3uMIOK
B7H9NMnSSpQRpsMeBBkCo7MGEKzvBB4eY81So34sdqY9R8IFS8FTIvxtWjUG48aM
tvT8Kng6SrTPH52ma8Nlqrl3V/KantGBOzmdiPPJPBl6Qkrtgjt3yln1L8Y3NAkT
/4FqXy5BfUfCxF8+BgUoZZlUwnRRsWNxOcZK0W9enrDdoFXG3fbabwPO6BYxpCGO
NMRtsr1zujl7yXMOdkU1ybT+YVYQ3mVCytS2zcrV0fUD8G0fZ2u+OEyu4a51gd//
Nf1PC51krBvkHyOoSTkpZaYFBk2Zn//Dxx5eRs8W5qYGNROX/mMfFrc3Ahdlrg0G
i7vAE74FKzfadR4nTGFC8No0uOm3mqehl0RX3PdvFwZHEnG4WQzdUz+ygTq0FiFK
PN+kctxLzfFFssrYDtZsS5G82xMYco0/WOlxCkkWkjIUy9AXlS+gRfJC5QeOulC2
ifLi6L1vlgcUseRyN11Zf4SVor1s5fbXwk9ZnP3anatr7QVfnh/ZjKwCcRzaUqPU
02wBnmiEhk9XgUQtOgOMdd+G0NQRXpWKeO2PnF9otUyANETJMCx/ep7V5PMd4jO8
i9fmOzwh0HbV7Sd81xoHzct76nEZGQumxzxoxe7lQ+blH+vt67l8k/9fPB3O0Ajx
1c2qUb1LGQDppw2Zg5TG56Tk/Ib2qLikRMutjNSkMrrJwFhStzJ2js1LGbg+BCdE
NpDvnrloL96qq7MfCnClVLp9smQKjkVlD3+0ME1GrZLH3v6GOvsipHvuBpeUf6zD
fudrh71QY82ExPfOfinbG5DLhXtUC4qG9jkcBcAZPDa/8rgt0XlI1JroJG5D5wCl
Wpx0txymwxoT5uUgSya+iw80ICveePtdozx0L+nn1xcUYAjIU8gN/ShR6PZTA9U2
GKyqESttIQYvhedj9+NFJUDqJsXNybam6jYJqN8gZm5xR4gRERnGCl65B7YVza0L
tWb6a1RtRkY4PioqtvAwGAbB5ozK1zzlK+6dgh/Hkq6xniwpxTS/vRVF3o87WfrG
iLBD8Klvhb1PUT4nGXhqHTahapjSPCItnkJAhCi0aJf6i7OF3yZp3HqW38hj6fkN
GP7cR8KrRFarbynHoZwb4qCk3puRPBcQcrPJ10qfa7bZx8o1NHDDPwKC6/9BSWHk
/K/gut5KK/QNDFQTNeYrLv8BA/s9hEhC0Gf3EhMsGZUrQwEkFiXt9n0l9xk3hPb3
FdjHE0MpUOT8I3+12Iqx0edEpcSJtlKL+rdkqBhqW8TPOeBvQ3DHuZwMr3bz8RSH
cy9yoIQH+kk8VIMSovH6jAy2rfahuayFbiej5+0k+tWI9AD5H82RzNVVCetUiUHX
GcwcKa60BMsKc0j0lYHvmWatoo2eWde+4ud9DWf8StZMAFEA0UBD/Gn/gLhEUNyr
b4XHPb4evtOQdDui0BKw0lyuLLgVMqH77KC2iiz7M8i5m3Ym+8cgJoxM7xPv8brw
TikunBjLcwZML08SMjJs/hrYwvDnSS+s1i3REIBYVVgScZzzbbcYvefoFZf+b7pa
ThnZOPCcDW46uBgskpJXkXcihvlRrqXEgOXTS+vWNIzFNypbE1WVxD+EiQ4kwfti
Xolx44DEYiPrnzGP5TE3k8DErs+iEsktKI6hEW1kMdJkg0jjkWgFb9apDrUu34AI
vwDfy7RXTR/JL0opdqhl38WHCB3tG6vblYFAYdCSUNpWOOlOoUZ/q9Dd5KAsVqg3
M1XY0606MWs+RY0vcUmN1QqSSLc2JtNlpCBZ6K4Ten5AUiEdpARFuSm/LY9Fhn1x
MJiQFhPeV8wcMIGk0SvdiyPjv6XGpJ8OdFRH7DeC78AzHLSHeFcxp+fhQVl9iTmO
KMcmQZnaimYJT5cwng83h98GO3XqVo/efTA/RltYy8XZhI8vntOBvCeU0gb1GboR
6sPodXqbRi/Fs9X+iRzUi76M71FD+q7c3piYH8jYGYO3q21UAqC7Mem4xVzqwXpz
AyB3nIY/5cxC9PWOKbFWKUGA1EcRYEFHCaNOzec94lWf3pOgVXowDyROeiwRUNeL
Wutl48ZI71DDzO3+rIAaXKy/5AvvDa7vy7+ix3wIRAXqqcUtgibBMujpk+1sMcpz
ZePPUtOTzAfg0S6c5nrRMSOL5RstF+YuFr3TKBvyjxBaRtWn0UVkWVKEj/+25Tps
IXpFLI2GyLBzTtBK7lhDKePaH+/K1EnobhDis1XIdYG3XEoxceL8UqCFlfpmaJCW
7bPql9KvATpW8kiRexYA9t2t8zjgV/I7jHGphe0ONWJTtEkx4eaZZV+lgrqno/tQ
uebzIwYlyCou2DmYPx3xCAGMZxjRZAb9wzOpnqJzpbrkIm7mxBgqKI3562pISXE8
q77LYHP2wuSTwBLMLsHHpCkPc+iRfvcRP4zTraU0r6rYMl1Iz+qgvmLJcdW2Dnz4
skExBXM5smSVlc7OKfB5vQ+GY4e8CvCHWSmXfXtPQo53v60xpZp/qVsGSHB0dbKr
bK+WvZAEF0SGV5vkLxE4C8mPJ2kKRVzGtoZ8Qvea9zXlY0VlXpvpaezlxZbgJF+Q
FsQmhQ/SB7ddG40RioyG5Ke5WV0LmLuhM/d+fXGtw2EaGEgi8WEF/pVSc659FnJw
WykPLIce9Iiq2PaKGMUujkf+xRQduqHnDPrYEcrvjD/aol+QxggM2tdtwX85YeeZ
+BPVDEkFIIHvvCHinkcRz2YupbwW98Rl5C6eowKUqa8uMej7O6khS1u0/oBiAqfF
bHD7O8834cAVCauNZMIJB6COMEYDsyMl7Bu4PJAtH9UqVoifP/pOX8/DkTSB3NJZ
2FSWMgVtLmREX1bt3bFZWnRznJwWI/KAo3Ifh+/UAYcSGheVaM15I7Kqy+1wmEQ6
yiPHVQX2nkg0Ctv6huzbvhyO3OSQWFReYtZTFhqQNphXUO0ZSx9M4efkMtohFZYB
LfepojD8tz6z32BdINZyRVvloKaxa3Q8JTY1CcZv/kqLicMQbqmuutIk/h7DWO8e
4t98930RWcrVH+SDGsgXSM/bMk5NMpqrrn3mINXmx/pDhX6RNmocXzB/xNPDyOvy
mODc6+TeBVIg84eDeqxA7fPpbnsKHLEByzMhp8tO+BQNUzKKtz5Jt5MyWy8WdQ7Q
Cb0xX/QbDuV3lKuwpX1EbbmTgCfTBQw/JIyCbv0NKdZCuaagIKQioN142TVXPdg2
ndyk2LXwgGsvfMew1+Pmo83XHSG7q8dMFz5zebGFl8O5Baed5o+QzlMoXhABVXhO
F39CwMKyDzVVtHnrgD6r7XvkIIfkFsErFr60vfjdke+HHJErfbkPpfwkPMPFTvRZ
gewruevzxPfntdVDyWmFqGC26cGm07GwmTjU54HyfROW2E/Ik8JPpZ8xKF0CAfzS
T8DqNVbYq0M+Ttq8g31C7X05kdgzZd7QAHyHfIo0iJSDJ+7EsGXJfXhDkm/8cFQ9
8H8pmw/fGfwbF3h/i2YX8sGm8+PCRxPiSnOVy+xSoKgay5/twVPGz099pmxhrRkm
aUENetfsmjnmouBPlDzPUtnadGmqDvwjjecZ96iZk4R5rXHeXPr2vUIBk+vFB7pS
3kl6o9gX1ylBfvS1qFAYBWxk5O9BZVi60oeqSjRQCWtzrPhvpfgm4MPlBwq26+tJ
CGbMhDd31btp7IfgpNFnoXMxylYw094F1eLigPMEQz4vLIRTADeXEGrTWjqnc80S
+lxHF80sKHNYnzDFmpkQC5ZJGm+NSEVSnTOj8105ExlVmRjZ195/9UhJM1cm2Mlv
xsS5v48v57EI8dYuEXiJJtWvbBm8O5iVyMt4dABcOf9p1Gj1FLNSOIire626xRrG
edEZy3Wn7o1O09znYh7dEWNkkNVA7oUWDIFPfs7T6ZwKyK65p8fPuJ/Jd9CafcjE
OtSBeMvejRoFIpJYo4jeEGsTsh1vsp5DYLj6J5eNS+md7Ac764Y0W0YL0rs/ZO/8
uw5Wsk9yBMZGYzK2B7jAw/0LzG61xAe3HPBRT4W8kkGHpGSpmrqmGMDgreW5kO+R
Hcf4LsoQVxxtfyiHDUQYTWF/2qZoKT8ogtpoF1HB7NzoYuFXB77JRGq0FwD5C9PT
iwDIz8bQEOmcLAEPRgRF5u2h9oExPqrH9ZGaPNL/bBlG2InvdLAvO+1DWzw20Qjd
NERMkMC2lz+FFPOCrdt7e3uqWhh3mqVOM+9EId08MDRVCiCiTk5U3laR/3G1uFUU
lbiHRd166uMYl2TKOX8+dQKrpxhcso4/c8svdglbCX9FNIUAsKwaZiS9we4GuG9z
1Ee0irxSRx7rIhKMVNIoN8EkIqp5BTPV48lgVYB/1wKHqyXvU9eyfHMFec6M5zRj
fYek3N7cuM9TMXqhrkdGBXuZTdU/Xglwif848zgGrrhNavfTPYNIl49HyYNDsVoy
i/8DASfsxKkdrCZktsIZQwZwZ+/BggYCC8SktGk3XnaE90BvONZMXyzE6OjGITVH
97SjVP79Jw9x3ayZRlyKhGNRolmDjNBk31vFROHsTfBE4FNGi8Dsf/zANmS2+8Q3
sJVYlzj7+n0cVTB1B7nMbAWeTxNJibSRxepGNkWSEQyePGnD6/UowTUAxiKu/nYO
ASyHNUc5Nj6G/FDwlbmhPcRO0itReyRUM8J0gn1pFHb313XrXgy42PuBSL9+Kxft
iK4B3TRoHePR9+KghVpqVx3h9ZusxevUGHDkr+xvJWJwhhD66bLX8uQFj4lqubNr
2lorjpAxtUgFNb03PEvDWLkE8GB4IvMTFdsUL7mWwPtmwOupck2Pz8iZWKA+/1C1
UHlfBwX5Fm3KYhEcD1/0QYpIhywgEPnyRiO4cZH7B3mceIHNdmD5a7NuwdDH6viY
caxga1YseIf0cbE+BVhM5XrWQc+8NjsB1F6EXHGCnsSu+n2fdXUveKvsyJGjtnig
RXkn13XnPug0Au9NPDCHcY+ShrmlfJP7YfDrGMD/fq9aKSUO/Vgld2llUbiXzprz
wV/91acRlJdXbe77bQ/iWJ3M+3oAFYH+kFTR1GkXkZD6GMdQBGDzs76hr2c1pnwR
axuc7Yrl/WFhM1wSLR2Zex1rfC4SvjYw7CxhJJ2bm5iJqtUwQ8gF9qNIQkGkcVKw
aRIGD4AOjCrg5GFrv1ZMrCDYCnlmPayQypt8AKldDPIknQfrFmpwxikn04ZK0Y5U
/UTL2txBHtjhQ5elO0zjE90T9ePhh4QAZ5X+I0o5JbqA8Kb5DrzR+/7OzG4FY8RQ
3ahoe+MhQHhfzWfKynLSkFAvLgmBViwaexTn558OMl494dRXuk5TuNuyH1dFRrD9
zQYA4OCwqJxlf+K4Krt+hBU9Y5hStLwTcl0USS6Fukn3eXYxDnQ7F9IQUWAZm2qY
WFKXx0N4LHLvVdH2HgT1m1avrilYwANMQ8ISO2I/dIbg/iHGL9I9XHk55ocWkf99
Yqay6EkvT05Px4F8k25RkfiaYjLJJZjQR6P21xUuOy29RfzW1ZyfLym2Ee5L5U6N
x7v9j0UNeVR3e9EIPpcV4YzMj7sncmwIdob6gQKVezwjQ751LLQVZd1ymLJtLQzg
sY6kGRbOwHjb4mwEt1AY4Vs1hjdnLsG24jQcy5Be0e3aoEJRzuQ22SZQgeTlu/6z
ZFJRxKw+Vvz5QmEatBT56mfilDwVB46t1tvdhkISIHV54AsUCiIlO5uG8MOkj13n
gi5iSeP2qLnqz4k1aJpgWiw/MVmLFSlH4FUi1Hq3s5qjoxyPi39c1E9Xrx8E0WDG
XfPLOKx5AVR5mZyN3jwqM/tjZxzQBNDKz1J766IOpTbwvJlWnO5M6P6S8imYJ8Dc
P3BWKhliJ6BUyQUHr8cHw15+DyINAS4V2tElRF1so9jGkdFM5K64++YFYy4hOzXe
atmo/eC8a8TXc5R6NiTlKr8VJKWsa3pSOl2Tib0o9KzBbIv74UbPnSAau24cRwtD
+R93nMLuFB7DLyoy81dPalD2Cb9IkbLPwh7quDbpPN/YUKwzKZXFvCuatQ6trzh4
SgqhmUyH7r/NWZI2b0NL9jn5Qj2xFRM2pAfhzbPP7RKOt8IkdhovI4PHPG9jPo6I
uMw2bEv0OSX07M4HATA05fTItiWIxDp/mmbGoHTSt1UeOhTW3N8WvbDMAgwi3XOV
g6qeLWN6qTPI6MjTRn7nb78m5hyTwncYm5IEYzaVfXU2RAedysY1mOkXUaRjtWdL
IL9knKdpCbIzAYXO/hZIrBGY48kd1QLeuojv0R1cjS6YaOIGyM7+0Ap3F5/miTNp
sHpjt9RcIwfVETcQcxe2W6q7f8dbFcZtss88nPVHf007U9Damb+tIPe793KdtbhW
qGZK+/Af0xYLA3s1vJnog4jMZnYBeRWKnf5Jt6qrcSS+1mZBScfFpxC2sJ6/LdW/
Y3m69B8hCzD+lOLAE99PIoQmJ9aR5N4wnU9vH4Kcm98+z82t1pFQ+qfYdITGf2Ow
ax76eoxvgq8947/sT77R+lySAm2T2jXdKZS/SAKLMLSE+qvoHubQN1+PsBv9/YE3
WZZzoMKaeZxreSse8UT8BE9gauKFdAy9s8m0f7/2SgOv0v0VBtFF1DImyD5sAjMw
ulC54h6iLvmuoFtB75FX/znpnMPKrDh3YPAWDNmm3uN4tlA0zvpPLAQKSw9lZhia
VMT8c+jzb9xohmBnl/WCOsGI9j7kuGJePhH0hRm69EovZEPX52TmEUqX0lNEkk2Z
ZwDFcNRV4Xqsig9PX0GhXwCbnO8fG8PJ8CQc10nXWVO8SI1JxkkFJF4uzinDffN2
XbmxdrC/YdHqn5Ln/A5q6BaC4gJ2N2yTxrYTf5pvAQvATAb4SXmxtogZN5j0h09S
8LjTJjrORjWoz3B/BnKABXBv/AY5QMtn2CGWCDF9KR8VqoW6xg/xRzE/CLu1U4Mj
TjXOri8VmJglr9l4u/Y9gDOOqqFkePQq1xB1mcfc+/kgyOFdlg5EZXAFpF+0cK4g
Xbi6RgX7oMxMTO+a4miGkA6qgF9rHHo8Gd2NAkoCXvfR9haJqaDvrDbvB6CcLRjv
XInRlNSCHRzJdSzIp/YDllB7PYP9Ih3ARla9j0Zt2W1jIxg7jRd9JOVH+d5rOOgW
b39K8d+aH8cOmnBmXS49649ARPnN14wtsGwbn695xQQrUR5ZobayQMrKD+Ywn6Sm
W6V/Vstu332Gqr9oerq1PAEgycAeFnTyRCouBPL/y5BjPZeKZqsXhBafutg9y0W8
eFJTQtnDR7sKisaSMfPckeRw8SjfM/3zLcPNeQLmRLUpM8Umnw+ugt5oxfMHvGIh
0ZHUvw9a9TyQbJT4QBQFqXsxqduAW1Rx2hGNbU5wGmdcg2eYd7H17R02AjLmJHo6
mkH+H4NLrnl1GEe1aoE16QuDz6gIUKyAmbMIRSAPTNVVyibx0jE4dr2GgwGNUCfk
Sm41TVlRdxFZOi8jxPUnXma5SbNT/PyEUx7iIDOEhQ+QSLfPlPh3jA+RWzHsvAW7
ea28QDlDGq+cRaDMZml4njaP6OFT3WXD8xG2/g08HOfZMoDiaVtcfKTR4PS11rTn
mcOoNIxXHyyJodTN7/dJf6htcD7ruuHhmznDnZn1mpZT0V+9zZT0NrP5eVqJS5Di
IbC8+X683Ci4CI51ld4Lo5VUSbb2K9V8HklpPe4a07TC0Wx4T9pqb4HvtUHe6gyi
BLa+JLF3lwAPujrDXHbMXRLopCPDkxUalkww3hPBYHMmWXXRmi4mTOTeamq5AFBI
2GvWdQaBNavgs0cvxMFHxh3rB5kywGLca/yl9LJPdgZnhWLw11s6HXntVuKX+9zk
DrNII2FZDzp9UZJihD0xsgX6ts8MAGycuGYtl8N2fltFL/2OaEZQIqgzF50tS7yR
ivuDUoxbQHeK6TZmp6soGpysuPFzipN+ynui40Rhip02MW/5Lk00Prudzc+AtzA9
FwQq3jeuoBZW24k9FsyOyTQdSHRgg54W8REJ1TIkU6ErTHxsBLZXiD1zWlK/Olu6
PjJcnzUp4zJPmtPVxAfIH+N06Gb5NiL7OacsKlXzy7OyqVf0kwbSjwYtm7Vy96Ri
/0bjMNVaojHUjcvw2jjnAjlw/fRssJn+UyzI+y2GMNI85cg4EySZUmAJf65Yehqj
V1NitYvkEY5nMuHn2XqwSQipIAe2x98T+NdRgUz4rBuDbMRI8o7DoEpUMixBsF8K
EfuM3dOaN/xUPmbjdtTtbW0lYIutxlP5RjPbdLD370srnyxItMbnYcSwmTwq66zF
+p9E1LXxYMQPc0vwlWFLk7tZnytZKSRLIWlnd/CzMdDN+U9TxsvMh0Y7M5dXA0ng
y0GhUvZJl8AgHR6+R1txcqjkSvPWKs6aPWXRK/w0ZrJGd7TgCPRLegdjthB/b7i8
yZB4Xp0AET+Z+Fq/Yi79HI3UAlhSJiEa/m72dpOZ35sIAw9OOPITOygEKkeOFmTg
X6oz3qQSdkl/qSUts0fwUr+M4Rrh6cG+f+f8MVEE1m618yRk8+netY6uWKOJZ+6W
6iWTeo4Qmiif1XeOXs+rXZ67dJ1JW7eVgl6Tz3lKoIXVWztHVbnNrWEGEpqeT+0b
XW+Xwhk+IJkaXNEW9m4lAXR2YJpuYD8pnoocDcBiW5pJw5TBrC/5b0WHfUituRHo
R3Kh4mVL+89iToEzrkYF0bTYv6Ps54x6+w57i/RfB+kKMlXFhQaIHgk0E1xo6nVF
VNBVfjQ5AnFBlSMTetFrt8MBzifNzmoz2h1rfeM2/PzzPMZRSTNQ+wTDQrcHJI5h
2V+d8d7No8sG0a+i27Ai5oZqt4OwiTScTg8VTwG+bqU5a3K67wC/m7WDkz6ojn2Z
m6dXuQnpLzh/Gkeb+UeT5N6RzPtugEXVyQbu3exJImZGH87dSrcMQoujYOO/Dc7J
9qd83RISAlq53aKdcFbEB6z1jYG6JoIFsuiUdKM4UmXuD5aaUqxgDIEafo0bqtMp
ygTfZ7tJbFfF81eyrLE9PbKSRsY7bIrqZdtNGJSEgPw237mWMwJkL6iNIDPBwhyQ
5T2mMLw2e00nIoisqsvS3PRDchc7ZA1JAGNYVz7gPuIiorHo+ln+otUx5sN1JgCz
8o+iPj9MUvb/+luLZ2QqTo2oPgQONYMBGDHd63WeWKKsyCeznIB1f/mg/adrhXlA
kbKJHb4C7nVk7VQxsZaqg10CzshLE1ardNyQJS5hQbwSK+b37TcaBNRNxCq93oWX
Z1hyUZh0uu0KL2OJaUi4MRtrsHPbh+Oqq6MYgk0GCaeTFHGJmRVh+xcXfSFbqm0n
wg3x3CdtNSyuVLQbpVYbh6uXlSw4dHNdF7/7Gqd4OqP1SPEyNilQzHdnnfGjZlPF
s1694E6F/qVmaNTvgg/M7ZcrCIYeWpxQOxws7DF7bFQ9k7WL5+IhDMax/Flj/ilp
64KkQ2YH9VGraybqf69Sj/NQetQZ4QN7YLWd4/+VBmyWeT8igRViZiVvUMBiXq4S
O+Tg5RxMuNmt1edGShqTrJsMCSPb7DkbwE1Bqg6pAQCrL4Fko6wWJCXybVnhIGWD
Dz+3K9mVUK9DAf4sHglblMLBBCuUFyG+NRYKIk8fFwtMpoM6rDqk/ogJB4/v+ExV
NQzbLPOcXY2YjhwoTqHUAVw5SbzFN1ahZBKUr6v/VoN59Ppd+rXRpAan39DC0zlP
/HENwiuNjo5zjgkoPe3qEw5vME+NA45klvSy30sTE0IRld0eOnIwR6ChGCnJniQA
yWgGq1+9wpO1aDqViJ5uf/14udyhujX2gX7g22ag7u7VEJ1c6Ysz+z//FnN8f91n
9ldrY0r3eCkCMQu6mhmHIf4UFrbZLOn8Y43/tX0cy6DjeDnrWfVzpVuXBE2xTxx1
Pv3Z1TLy1bZPmhPkqARJcWES5m+9DHkDt18oxurh2Az7NyaNkIbatzOcrwD5lLIh
bqvTF6cJuZG80ltOxfrhivXtQHFBzyNixpdKXNXc/qjlDmdBW5aRUJqJpj5qAZfZ
rXi2NSDeVTZHnr39/PoKndohjVpiYIMblN6dRYUo23yfv2qNs2T6m8OjvntSmkFv
XxTVVXx2soAK1aNA1qixdPDHij3g6KpZRcCbzxhuwyJsTqolCc6hkQDobr5vK5Dh
9a1e73au9ddPagG9ncKpLQRzQto63WjQ+1GQVjVcox+zrbI8Tmml/+R47q8jOXvL
bvUJMBT55lm88xgZ1QkptYqjq3/9h+puHTnkto6WOJimaSY2sON6IF6ol+RtEvqs
hweSImqB0aZK69h2NWHOjDvkhe914yYjRTccYgXrbh20dUZBwrUf7rDEK6PpaISz
JrTVvXWkLryUNpFnGZPgEA9FU4W+Egk+0JiSCgbbxuWW7OTbLJHI/5VFrfHmR6oL
YVIZuBQUxTAz5MSseDW+qLZsE0AyuhZNhPLxa2h1C7pdvyX9UtgcLKU6Y9fNYjJ0
2rePNiwylWce/5zHInEu1M56EDKn9r2K4sr+pj/8rKQwYBR2kwP/2S2juALiyOU3
ijrqtSE7beDJfe3VAtKFzK2DyBg9WVw6cB8AY2bQcOT36BAR3JOccHqvMG2g3jZu
hc4B+3RcRUOXpC7gAoVGpQdoijdd+i5gl/FmYyS/Dsyvbe9OmLVIVNl9nXhAihEL
AoWKJfJzi0QxmIOwDyEbaZDQ3EitsTu0FbSJxswnWSeFdM0aWZ6HYf5Nrzm2qF4r
9732JUGUytQyBoH4b9UAeGPOPZv+5bM9lXWjp++tznFk6mDpxd1+92fmoNVrz5po
A6BNdbj2npsWYgkOKtbi6IV45NMJMpfEGriJ4dfoeH2x71GX5Rpx2J1OUieWxK4e
QqKuJdl0JjhCTQguC32tHOczwqXxCHvLotvF9aiVJap/Rj4tc8noPCMUxI/zoXMt
Ydt9ZoDKwQUZ0qxUE1Stge53ADKZonX5pKRxtFzAi1ahRaw/XGHeL+jHiYGGADmH
PDRjXUVQqgv1xomcZP6+MthVTILAU29XK9MVOrh++CvFX4RBFKlnnuB2vtL7AluT
FYpBFGlrhNk/QpQpJZO2QqEG+SrGFMOI4MK5zSym9F2AILRxzkfQbhadGtKbrCrk
+uvAY3EsSKVFXVHsWK9gsA8Y+BIu5A/ltQUsvkFyDYel0Rdfknw8+92qf2hp3/Pu
ZxFwNPXfBs4fa9XQ58+8ZQT5vlXfC/PhdnlkY+FZ+PArkTqzsqsH51zLaxJueEmu
yd9oLvmPGL+PHd0m1NZlMvaxEXifFn8z4ePC2lIt20ofTADj2A6qm+ECTVNhjQ7o
n4O9zXV5xiCP0Z6IVEw/LLMz38ODPnJoDq8k9ye9cqfeC+8HcDpBQrNkAiexySUI
mrVJb2Dou9WU+l5jSXnFYQrJqrPDQvjnE7z5JXag/HCLS1OiYERcB1CsbiOxhVA7
jAraO9gpVNLu4D7hdSYbEqNfKXWJ8rTgUBfzSIFLxFCociFdKERnHSeR+GT7Bgnw
rqGhZzyVXPMy93JIahUYJZLOFL1GJemRRFhqBAUtYjr95v0I4ABBc4f6b0OjFnH6
Ve/eqUiOt0M3JejKvLaLBNiGf32ZOa0uhT+OZIROsI2PYCm/WLIeorvLWEegDcMy
QlKhcO8PXyE7Tmxz5ECb9ToQ0X8Eaq3CADcBuBaFZCZ41GqnARenUptEDzWrAhnI
PlZpLIH5KmrH3P1Kdk6+UlGhSrkwy2PEZV/X1u8wQDsn/dO6jUwupiV0yf8jfbH5
1bhZfePGs8aHNfvp/6SktnBDhFMYL3n/nSc28+f9UbNlDGaJGGL3qvacocDRryDB
hvk0vdQv1yy2wKzOtAbp/9Tic/w+LukTAGdrT81aCc+h+uBnXmahSZOKxU9Xxdzw
k887HMFFBSjMCGoh27/dKZ0h61pgk2emRf2S9D2RkWbQd9yb35xeAikEDNcuwHKg
iFcolY22bm69bDeVRbr7wK07XlGkjluC/UvlsWKnFnAZsfmFwkd9uX4nrdsEyqvb
TlxftDSqwwoRNbpSiEf2X1At+Q1E7bQvzHqq/H1QteWoUuqrDmsj5LLNE20tKTUw
VLOzFPmCwVCFkI7yHWTVfQzOwLPOpa3Jl2APNPVgQCiqm9jajmMnfp9vJwI3fs9Q
TGNkAE7cyd1fkD+2D7YmMUlzfXH5V0YTa4976FjxqMVhsUrCnDXbjT0LbmuGxwPL
/2C/W+f7ftgIDu/gVQwSrb3otRT9ZwOnmfEMR4wjS3Ixr/XtBJTf5xzvP9NxnCcj
pR2zCyd/AWvIn/ztCbc/NbwM4eFkLlnonE8PU4TB47/caNzJUYL1/EnHrjDq98R4
gy62UEDa30/sSL7jxkYFcDucEdj/7gTP69nNPkSiYmPQW9YdQqp+tkIlow0pFi1R
Iz23BhEU0pQ33Y330TrHVMKyz58AhEuAiC/bA5QGF70Qyt4B/1h2avj9KIIF2ip1
J90c8P3S1jw4QwZ5z+WdR+fY+pM9iNNv//ra9A1h0c587Lb9FEVJpbmdXsREiskx
h9Q1D6MAwXxCRwM1+wDsXDKMYEsWuw/J2Ws6tzbcrfB3bIOnPj4/f6cJZOad/9UK
11Pcjci2CnkZ4IcUt8xdd1yP4u0UT1+SjR5PJuUhM2PG43zeh9pxbeqqOh7h06PP
PW4qSktL9KDTOGXOnptsozU7DIOP6TmfMR662uG1lrcGpRdIVfup4n5xRTSaYS44
yKpJipQ2i5mM7jZ3ekNaEMPh1f047DwGhfo/K34DLNeJMN0hNt/mERtz1qrRaUSS
ViYEpu3LOMGn/HEQltTE8gBpWuHNhJ2dqk/PKU52qwAchb3V14d6GHGQczxPI7W6
CJuDhz2FQXQ9hB3jrqPBDA==
`pragma protect end_protected
