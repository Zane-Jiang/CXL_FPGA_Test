`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
MU4NBFmTmSoioQLoHNz58VkN9UnFKL3hUP4q1jb3FAr4n25EOWW+aojoH/oayLPT
Qfffsrgc/lL6TCBxKwlJwRQm4Wyffme6lGuiczH6vbNJatGyo4YdTUlxUBmbEI+7
buUQ0xatqFRrmzjN118lhp5layilB07b6J71N295NCE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2240), data_block
fTEqPlcdnGeL8fnq0mmJs7ufrBE6MSbvg5ntJhDfHFSv7Qo+A01uoTIRdKneTQlD
ZA0tiCg39anFJCPPkhanQkhX8kLY55hxMiTw082KfC5aF+Dlj4ZuRFm7YpIhtDHy
Gx9OlF4tr+95InAogroM/l3JDmauzzIZqixVrawyjv5h1fvh5bo0IJafFrvaE6W5
UEGGrU0/RwYBJdfxDSfqpDui3kJFFPrvFOpJfaEJho/mdXY1gJzutTmdFSy0nN1K
6vto/JwJcyJjoOupr6iQpinwm5ymqa2onV5omRclV6i9Bjiq22/nN/iIalXb1XHL
Z8EFUQwC3xkfU2v8xr6CQqdKfPEWDsQyTMjL/Hp5o65/oWR1R16iJqjimiQtMKCJ
V/8sazmjlnEUltC1RvRZZoCb0S+dvE8wgVufjlK7Sf9DVYT7dKsOTqroRjPyjJoS
kAA/7YcEMi0V4lDov2d2s2K0RroGS33vwVFt4W798a9rUiOgTqXU7pow3iP87rQY
tl/lej3CrpQlUGIghTDFcAkGvC2QfMTHXJjB7tGmJJNI75DcAhKpqek0hL8DW+GZ
vUuDi9X1iGc6dJAcj2fOAerppKzuEGUa3rgUfhsEBtLWdbu44abvu3xZa+k0tXmz
B8VRxhFO/SyQkFzWryCNdlgZRklHrIYzhW5YICyh0cMdFN4yVHBDmXwHyne/VPaS
24vEkVy7xWpmeqD4AOefk8CdeV82e4o78bsR+jR9vd074g2EVX0wtihSxCeG4DoM
z9afDYvMnPIx5rAhxYy7K+bhzg9K2axNUVy91ZTJPst38TZvOoeFttugGPl0fPOU
b2oju0C/1Im0x+UuXGK+OAvHs60yLDm1MSSBsd2bYxhejzBczxzfYteURNynx2C/
wrAbkgRQb6eWZ86bNGGyfvwDySv+Cpx0XMN6+uKrblY2u/UN8Mw7uANIOBZkvs+6
s/+eEdsQeUDiL1jDw/aZcU5+eBSpe1OTvqH32/zeuYSzXxPtUAGbm0tqY6+j9qUx
2KVgpejNrJ6K4LYaTdbX58uC+qzDPHY6yrx685/Yd3BA/P4VCzI8CNQgdoIr94JJ
ytywXaSqRjNPptX3OO3Z+Bgqi69P+qjTogYS6o981hBrjFeCBJz7eU4asB1LVFTq
QrKnNxPUZSfm7nz2b54wVXdoXGiJCrY+xgpVHNX9RzImjyFiG+U+DqANcO1tKRDY
SNsYQUskO97DEMVT9L13s6dmzMq3B/gY+YmkeufELaOVGKZ29mmDpZqfBT4/XQbA
EcPGUHLfIEzuhxbGOB/cVyXk0GCsUsZiVGX5Vhvd9YGnONr763vpW54QqkEKjCP7
/VKpCPKL6shY1615k/81FjCGj1n41bfkbpXjU6EK+tN5sMO/SUlTLfW+3cEBCi7f
teBWrNMjBnvU2T424LE1UcYWzUAUluKwqCg8KkFeVa/s1LyfrUGuwuCanj8PQglw
AGF/G0+m8Va8RZTXwqj2lWMFNXTgucpWdWEwsjBh3cZL5t5UBEvKSHfbBJ2pkree
K7Y3atyJd9bhC8M9PcomwMpw/0X2nMlR5JMPWa1w41o1Z4GigLC8VlInCW5zprku
I6QTKOAV78Vf6YJ1Im9M2kDrm1sqxJS7bFB8WA9rIvdSmqzN6hJSxmAaQJaGFUlY
jgzjH+39XWSc0Yb+J2jf71c53RTZbEOurNkFKczRVdK+1pC51WAxKUE4zZAHX0vt
+Wnrdax9JgyTmY2Q9kcMmLY5bPXuSjCClCPKw4fO5m4Qg+xfGE/y4QlGdiBuI9jl
5qnHz1skRlPVdBTcr8kioReSg9ybGF58XrvJZnCA8M4JcSZ19yJX3h10kO7jm6TX
pyTYDHaLYwzWExMYsKqoHfpPZCUDYAc/O5CneBPDg65BcjzjA1wlMH2PMYfaCgFh
z9jqRC2bb+RvpaYBhEEyzKxhOSNQ0CaaWG7bHgDhZ2ildYiWYpWxNDNhar0OYyyQ
IDb+0I4xQ3JHIE6Di4cqQrpfIDUFMOLEu5xIQeZpbhU1eEqv9xE/dzP1YADLrUjU
w+W1XUdApnerzGima5F/WdEXmg6ffAWAiA7OfOZ3ngknMlw83p1Y+e6BnuSLxZTg
ZafqLmjCfAnC7iJUuAKFo96wDcLwiqfupnfjEKFLs3k4Yi8pKdR9AGEmUZ1G8Qck
y4md+VrfuXJAnGUGagJUBvLdYMyryJzWb0gQetEfud3Fm15xtxjlSctlUurc5JUB
Jna7uw/YRdw+swFW4dfYGvjtq845mHCESLhS+DITJJOK01o+NQ9egfXEUObvV6Pd
CSvn2UUe+3x7uaVaxD9MsNeMz+E71uBLk7Oc9GOH9nIp46XZdzrAx9RSoUgZVPdU
YxrzZYvQjv8pJMnlmaSBD1DjRkxHklzEhn6JHD+M2sD+61JAwaQfroWMxfkJkzJN
6N3FQMCsotqF2GDJjvaV+mS2vYJ9MbTmUL+UX99Bkkv79D+6KsbjSkCdaMWFnhag
9rHV5WcOjh+yFi4UNk+KQA5QfAu8HSIEG5vlThBe4x3dx1f6RQzLCdW9hwHfc1/4
9zZTxMZe6ImfIrc5E7SJPw5Z+S4FJ8ZEG0Y6PjPQ61wEctljPHRFhouOX3VHHH5V
dLW9RiWldfC8heJ5PUVuYiLREk/sEV/QklvDn1kBdGCblHH5ZQg4H+SWu9HBDlgd
U1SxVEtf6qlDvgHr1tjBD5DOuIUT+itGLgK3B8KnPLkPlrmzT9Ndd6saPDF6sEcT
v827uqOmD20pqogEfLCEWXkgam+EIO7zonCVLUuU8p6YUZfD9h3Mn5eIFdYlXRjE
0ljEzdh3AbL8o2EdPhARO67x/mXmlYrSghFZpo+zSHKwxuV3F45+ExBESACFnPK9
sEaYedCLuS3/t8wICvwrkf18+e77KmN5sQKqC9ky6q1/CzjqEGr+ZVh3J8lctelY
6WKYWhmO9myQHkM/oajiCfD32a2x4MWK5Ct3K60vHaE=
`pragma protect end_protected
