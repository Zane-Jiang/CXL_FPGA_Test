// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
zWBIud7htTB7soRui7kZ5Sf4CXEPL7jYOKIfrg1UC+rpZhkT14mkFsS/6lmf
rpHCCH7wrPxJYbncIDn69nPxwG6Nw/dPAJskb+BqYOpzvGyip2MVWcrKLmIZ
arjHOIuQ2byApiv/JNg6yHxkk18xyqxoORRwMNcFnvRwkD8dA8ehAhfP2YQ7
A37N/m/VSZHb49Pc3ZVtZOCdIS5ZPhcL4Zvhm4g47SK6sror74IVgoSdQ+Xf
ZqqH+xIurMMu0y/7K2I1toRyOMT1CqpY1yMx5PuMhB2Le4IbbCef8LtMXEK3
ajMXjSeMTjfa/B2YvJjHRQEBvh2+1em/IJxClcXh+Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
P6yMv87kgMnXFghBujTnIGKHcAMC1FZ33g9Zjdiki5K5iis+OQiubykDUyGD
Gxo9IxsebSPxjHr1UI7/jt/q09kJ8Z5RBzlhF5nL/uaHbV1K3K+87GSVFG+5
7qmJaovXZp5Z5I1JLM5FcQG3XeLzuL1IqmvgVyLIqoEhcu9mh6xJM0YvbxGJ
ts02AQAgC7obPFuSM3w/Y3M2wGHwLPqfnVMlpYwKJA/qU6VeDM+2qDPSHDQS
WZBecyBJR0P+gqDJYL26ZKeXHqjd3dcH5qZKwSHs73hS+kfD6PO/RiwC8//E
Lm86dVtKudqQ0vatYWvnMTGmNhzMtw9Ca68oKCLgyw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pN0MKZfMYGYXVjYmqkZ2hafIB/YdmF0Sv4W4siHKtu5jbj+G4gRYjJzlIQ3/
SXrWeEm4royJ6+AN57Au0VfU32O39is7muCZjZeB2FdKfLP2hPGsq0woLVmO
ObCQfUKDduaWEh1AufHZwh+ZGQB7o4W77U63RAgkzl7Au6UfCGWbOOqX66tD
M+mcBjEp8R7xYdWG5Cl3mf8GZ9IUjnoxL3KYn8oMKiejCYyVdRlM0hcGUK4n
51aESLn2iBGPU9XTk2nTchlTmOKGbTB1HAtlus7lr/YRps3NZJgyIechhK7t
lVh3ECV80bBgVZZiYJn0DljXjTHmhV4Pdwm1ORGeGg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
f7IfFso19Kma+jmTMyJa3E94grAywCIyILo5vdG/O+dUUSo+8WME3HVmzu+f
fHusFiEQ/YyLTc1sCC973OQT2LKu0MoRRANoWTPqM0sSkdBbNc8QGUeY9W05
luAdlz0D4EdqJvAGwy8AocQ6YhxmCv7ILASSPp7GGuCcGSehtho=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sWqQLgJUjWL5YxGQZnx+H16fIvFea5aiFBfbU7+PtWz2WoKhLjQiUKXsRZWY
BYsW/wwhoF94DSLKJj2b8moL1cm2ClfIJNVwnSHYFxnJKsEf/Rh5p8sKJO8d
5MphfwvXU4qZFJRSIyLJiJT/dtgeKXZrKq455PRebmrKxDoGmI8lrxmKZ1Hd
hjDlKgYvSW8VPFSA3hFsHefiPT1EBoCEff5BHYajPE7nkMer6i0HaGysn4lr
sIFv0LPlP2+cyWavZpNyu1YxRM1KUErVeUd7DVXVO/QzqDaUiPKmjE5pU1x+
zzr/kcPCMqxt9T5o3C0BZJdGesd96/OXV1uACPhzhEBMWsVYt+dynjSO9vXr
vMCdSNY3tjUWxlRyuLN/JcUnjuJcffAR3ooOUkHJBOOJ+UMHBway/9ZXCGLp
C+PtGJ/LTRX396Umvl00CEDtY6wwjO2FXZ3l1W+EioYBd3JenySrVOkbrsSt
PG+I+VOUJ6F7oeY+JU/Gdi6c3EHFW/hd


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FK+sXQYh5xGFxIWZXAKhEGNTkGn6clhAQCG+ClWJ4hZfdvi32mVTnYY6oDb2
Y3DIlSpMMOEZibNYk1Z8dD/eoQmQ16H8ZqyrP7/InNSRybpCwEmH8Sqh3rZz
qBbmC7ml41PGwZYwq2jvokDtxIsJeiSeAWp5JvYWi9Huy30OpAI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iDloywNjroVd527zxHb4ZWOrXTN1CQi7eVhNdBaR5VdldmTTWjbFgd3fbhyw
AARHAeGIOsHxF5XxXoEIa6aekfKWgEHO4Rj66i6UvPlQU1Vaqw/Cu20atTRj
i2Cf/y/7YODTYepLElFZ1HasqcFwnKxmHm3HMpP3iz/jOLV/Onk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
HSRTwC39kzyjTdM89ClwiBN9O71gVAUKlNHBBxyVGnjkwNKxMQKLm5ngnG3m
gJE7EpXVtWWzq63Pvv6KMgnOai44llLsjrOEFYRJu58qNojHaGTtbaVBmuvp
zp0q+finTh49jIhqq4QDi9L1YikIwp3yl6zMIBxFVfVcOm3tfJxwhUZCmDGY
S/Otcc+/KXwRUsKfEXL0bIpoEFdtK7/sov/noeCKfo+8UYMvXbPUDA9tj4pA
b+YVjmHHGU/4ZnuyRWlYFr+uM5tXSbdLqPUBPBTlEGAoV8Q833OzwO1SpFbL
PqeVgMX1Y0zlzrn1mYZdUtuz5urDzGK84kGKproepbdCL+ARWgdEk2stDMxC
XvxfunSVlmdHGc9N+Ms4qHSdo90w8UsBdyzQRHP8k6OGgz2m1Uh9/2LcCsZq
5QuQup8MW3IOcoCccJyCC2CYFAeFHTS30Hnz/+obsd9YvvBuulnbTSDta3Wo
yMiRt5Se7woE7Hld+cKSghvmuS2kKPHTUahzOLAV8/MMaHt813RINVrZa/2k
sgIHrDIfMPBTspTzEHscrgkkkVPjABOpl6Qrl9hrm0zqAiizvDRTsAbTZ+sN
cYnnbPwH3xEGhLfjzykhyzeT2TsgeCSiYRANY50nN37ktyVOQXPlmkgNWQF6
0QdtwpcsB/FZuN6r8sJOjoQgflXDM8ayPzJY4XAi17ZqIeN0/WNDUAz0XIvC
TdXzeSkoCyjQZ16OGva9+coJCc6tSpXdw+anZk0E1V8AF5ZugCT+gdzzTUMR
w7Tj8bkCEFTUyLlwr4E/ykQ3AHVneiZxT+qM6U+A0gmAc0CT+ArMq76a6ZH3
1sWD0ks6ekO7AM2rqFYuh/Pq+pzDeX036tFzf6RochmtELZ1s1AmlcmbAtbc
5U2YfHUFjBsGZbMUgUrz1TlwWb2oE0RP5VQfXwPi3i2f0QI6v4ptSXg/Oiuq
/OkEG//X59fVQW3f1giyH2jbVhcw8w/HN/XT0mLEYxRiOmIEBTGVxVQlL8Ak
eaPLZcbnYc3p22MI17UdentVVUtFq4YReLYvWunI48RnOYfuYPH9zbB/Cx1v
zylLUypUOU5xIuhUrE/ElNWFbw9CGT7lZOXajxj3aqCQFkvAybCgmSyCFWRz
yHWbDpb8+k83kvO2LRCU74VViTb7+5RD0Dxee3IPsCBIigRFlfh5i0F83e14
05H0rek9NyDelozyXgwoHpjG9VSv63FCz0wqRwVv2ZfCYb3EhO1DKXKkBhKh
OOi6CvzTlu+59Z3QjB4ZfzBuIsbImBiTkYYsvJSXX/fkCHynL1lUfd/QCFDm
FWRFLljhpCaI9PJmVXn7Mm9+n6eLY9DdHoYe/1tbi0CTG68oW2WHQ7PTye4Z
hW01q4M=

`pragma protect end_protected
