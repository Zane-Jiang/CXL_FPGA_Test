// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
59WvmPj4SCA06vtwBwg04M530n6QS0gsGoLZAxPfhFZRAxfFyp+5apPdGO/0KlMZ
YOTSn2P3wyUenLGBgJrCLnne4Fdys/Bd5JWrXS76o3s6AAHY2VVGQIIlYZllPcDC
NEIy6mgQuD5/ABo/S6SUnCxNZPRE9yomuDP16L7GA6jT/MjVnEFeMQ==
//pragma protect end_key_block
//pragma protect digest_block
PEWD4tBJhUqkrR8JGHh9teP7knU=
//pragma protect end_digest_block
//pragma protect data_block
gS94yx0MeIpXXfRphiadGHV32OThrRWbNjLQIlEQwF/qlE6Fh20hsc+q3hWImgMb
EPrEgbii5vrJYCgOPUg9oFCGsq0rdaRCp+JDxsaZh8jHKRoNAH9pfF66UIFG+e9k
0mcC5tmQj68E380jtYpQD+vVZP2H2uMXBnKRhnIVik3IdSqROV7z3rhSyaUZhSez
RTStUSqfWrkgiRIS8VVo4l2eiDt0VJSN+wnpYXJv7YPtm8bxNaHPs0yWNs7p3W2d
shE7udz/96c0Jfv66+vGQCY18/yVPJgK3/a5YzLxeSTK6m3pkBk3cjKmWBN+UYFg
VhxeNpB8vr11iUHf4SFkJG2aNqQH73uRJGXBybwQK8Hw25kKJtJeain4hc5EGO5K
zm4aM19zJazQaJXHtdwBNUm1h69QB17YDpcTV+O6HPIPKeZ4KwEtoHLvmbKE4vs1
1iInMej1pQCrLucvN/2gGeXPGBWExcLrpxXQrj9eZivMslf/PDITKlLj76Zi1dm8
2JtHeBkTydk7H/uhVAgJ9rEcfQN9GnyulMQnCjY4lTjoqqYTbIpObL+TTH04JoaZ
OZzLMaGEkYalEhiuofgFIlASdvInd/u0Ga4uj5obFWb6m3ABtMB8Eul0kzpT2kTz
0HQ4zMBTfVR4Jlc2JfWLHi+eWrN6knmi/8Il+pxOXwzh8qLmJPmH6d0OcTRQyNAa
UbDLunvPYBOvUL4kvl3CyDmV2YfrFAk+7/rSVDBtv7mCVEXCFrtQ4pjZKvC2lTdD
X9cgImqQYZkqSX4DD3o2O6Krjnf5OPubUHvcUkZoL9bm+mfDc1LYOAZrNJN604nf
0hY4iwVHlxzHUJCvUwlEey8Id2q6pD8N5Zu37uM86nyHutfZ+8OpehxGZW7MNBIa
Di/+73NLuwkPQjdKqYbGe1IE0mMc9wRJa4MNBi3u2TyRI1UVe0FLWt8TxiDa7pg8
TQEwdkPK6Lc53M2/TdU/zZD8ZHlJGijT+jUtcY/3h75AVPya7wHEfKmCbHaOPCqx
BmtXzdIDbVsClBpsjtY+cwmLaMjyQJErxZDv+qLb3yFCYr+f61NGo6zkytCpOx1M
gx1WPu/YGu7OKb8uUqSw9Xt49MlEAIg67PEFNd0JWnH3lAwdSeKg90PF25RZW8q5
G11nzx9BCr4ol045fz0Y9f+bz+kZP139sBG5qv1HC456H8EV1mso0rGYLirBnGut
4XAsfnw/Fc/2m0d7uQZ7Bhu3xBsZAEiLnX7SYFgdZFHEkJguLn+iLDU/T5N1uITa
gcMh4hwZboWPn/L/Fc4AUiGeZESSuCoHaDs8YV1zILHoO77MWVH7O1Lwm7aM1PGn
mIg49Oo6sBCeQKdn5Vc2faxc+vtSn2QRdPqo8p5jZY/Bicxw/p0qQVhuNN7RFxna
8W93EsMyDIIWxGxkjLXKjJQOAQjxnsiJFM6R7HNvwZPLfnFE4khYZmU095MlSkMC
aSF8+V5SfK3/fQlN2scBTQ5bEQeWpYwQJrEMCiW+XT385+tJpfXk1SUGkDIT95Th
yiso77EwwV+lyYsK5OENBx/225sKb7FPRIn4AQqqKWHT3+jc7tp30kjGVrYOdizk
qj/HLqXbRTi6E0RRS07F4oU/WvIpCZ++HKzFD2Y9M/4jzYWvANYmQexyfZXjfhYX
PvElhoYtaRstcek5i38FSjyczo4MuH61ZNdMKpF5/4hgvPkwSG8Y4NY5vPVvTfK6
wqQNwdW0pUXa2PWdi1ejcKVT2c1e43cR9thnkrCo/g665qNp0Ef1hi8JbMflaQ8R
XWKDWf94552XhEoCP4y2Y5dnIQWyE/aGKEr5LvUGaGNSmpqxlOjTyULF4wVt1RRQ
L36qVgOexAmE8QmIGfWx6L1T4BQTbi44WAnrWi86hnF669vZlBs6HW8ReguQM9Pu
EB38Dt2wL1kpWJJBwxPYA8bqoyhQU4aqWrrPYpJHn19+2q9R15L5TRYq0NYVAuJY
WxGgDDPdgrM0IKqVfzoeHvZ/QS6X4MHnUQxS/O0sPW5j01YirVEleTslUVaW9e60
Pfcoda6Z4KEzJaifq9q1N+Df0cYfM12ozQUebepsxxgjmgx1U/ZAfJbXzNYsCECc
iq11qZwOIm3puPSaBkPi6FPdOhh5jPyBNVNz8Hbk5yMHfRJ9/XtmnPajzm+ooOAK
1q0PyRZsGHige+56G6j5hkuu1hBS5cg4JAF8Wb6ioCSqFWSKFLwNZjUdcsBQh3Vy
T7mHr6UeW0so9XsS9/jChNfdH0CiGVl+36SQyOY92Jm1Spv2WAO1TO7wadKmLtPE
fOo8CJWF40/i8QF4SA81jenWApEKla9wJjTyoJpXZXEH+VbvY2vvX85mVPNlym+e
aHlZlVVp6ZCGk66Jhdt8Q/mIZ9ciCmBMCAYiFHj/HuQWeSFYNmsHVA5+tKKg72BM
BNl5oN+m/GCzqYWyYU5WJ+mKQi57O1USd4WNOXZFKoanoSWylzF9EHhmBjDmaapk
a1lb15gYwcqv3lcQK/gwW1t3XqNHpiM7enj8wBa8Z55/3HbbQUsG6B4+h/0Wpx1s
FWiEdqbH+kdrptmIzghPGWCcljrWnPHWicC1GuWYAqPEi9wbKbK60e2CGSyMbxAl
AXDuFhD+usLioBFZE/o3RhAQOeoTqPWfnB1kS6JCaNL56agBgfP0qtN8GcrQtMuN
4r3P0GX8ikfCjrcLCEE2+d5NcknX2FHxLlLPAVMHA/LQJe1WuzCQvX3dQWSg87nJ
asabLYjKJKZjaMaFjIQUXND0dzeiQc9VcOkzlsH6AnTsZvFikkigMuc2N5VIZ75a
BPF6NV3ENMzRhvEjEngiz7+FgvjZOxnit6Xgv74IcIPZ1feo2ul/BirK/jrpwMfL
Y0vvSX/L2T7IFibPB/Pr16oLrsBeQObYyP/8iumlqLTDMMH2l6PBr/fLcqx38E3W
p77c6HqukLZnotnze5+Zd0jQcDQ+441qM3FPXTMAMP/MccWg5wf2OY5gNW8/ADov
BoJ5MUc3UL6penlAf7HokAY7muLUba8X5qihkZOOjC5LYOjeaaxChie2CKzQ3Fma
m2z96homaePk9MgVvqIHKR1a5LquffSv8zdtMMSmzMcwWuqossH13Jg49OwYCbo8
05WSRtsyHkjKGo1+kC35KR9OtxetV3TUKGNXxHKElk6ln31wFOE+colsqh1IIbbq
EMhv27JtbVM/Cb2QAWejLDvggiUsZtem0PmZP6JxwiKnAmeuycX3an41blMH/P8T
A8oggJgCqYB4JU4QiDmp7+9i/kZ+xOgxUhHsaZtQetA9Y1gxwYrXaMKZa18S1fk8
GUQ4myScbvImMsSzGL7MZPvARdCd3KqvT2T2x4pQiCkyfKs+QZV7n8rX0fPAWzNd
MymrUj1TWn0YncYEPYX8j79tuWgNTcj2iSgC8TLMATARtg+C6WPV5IMVbst0P4fR
ZZLEsANm2hnO1hT/W0fyXGbLY1IG8UQkwV+RJCNXxtphQYmz3I/vhAiD1gyZlkQr
o1kXx6mwtMaT7/mQjJTrgPoCskzgAwYejV8C3D0++67PcPY6D9HEu3b4XXcMc4Ap
XqhmYOx08BJXNb+qm6TcLZvHLeYqt1NL6UlnF06bGpsrVJghCdMlkUHUStWt7YdA
09yTUd3d2+FAjhQ7gMXc2E7FW6RTgbnB1yrpyTWnS8YYGiKGMm1VDe9jElzu69Dj
Ho/3g2AamLycPdLeGrpa/3FfQI5TlUp4cv5gQDgJ0enS4qKOd8BFVgFtZsVUNKJn
HqKpGyW85LR1DBiScU9xV60lGeJEHBEwbID6hxcac/3MPXTWXczTcDZDNllH+DR5
0Bf6Ru7wwrVHo290WYdE0nw8I2TT2P7m5Zx29ljtbu7slRl0wYbW0c5hbn3lRcLr
SP28H19/Ujo90w6uD7EThnEwXxlnlGQDQ8gmofAof0m9licobqA7Hy+LlfDiu4lC
h45Qgbq3MkRaMFReowidHK1WlRNzI3X7SZpCzBZ/EdTl5ObJqy2aYban724JZe8N
6Qx0UKAzVANH9iaVxyFLBGxYq3qvxV+qqMAvwVg+rTnFdFDCXPKDTLftaYkaj/O8
+7x9Zn4ISivi+bVptvB+C47l0Ccx64hdFJ9aTj+ehGylDnuiND/8ODUZHnpIgaQT
pSN5MhcxtBBhpoc0+YLH2mwsOuhf65BO/ioMnpUSsFnahHPyyIUIcG3lrn/MB6sm
EdiJeZQAdZL+OO5mpSr/vrIeFaqfIeY8uppHCiRLgW3KMqTwu7/hQhQCNxcLW+fc
79zynKVr+Da9xuVXdbbwWVDFO2OO5Ccg10vKoZuNoD24hAS3xQSkDnoxnHYHegWI
YcggpG8b8BeUzCSFgv3uTf8N7FaWjpp+GLyMHwTWiJFKPyR7+sL7E1RXUtdOdpXu
yFvqcO9bz4/6TacyJcYFTLDei2CzD2q1vqjOqc1Uw6mMQx+e1/PYuUDDdQDJcuv/
50q4qdf0XRxxAYxB8oZQ9uN3VzuS0pQXJdBPrX6dVwHVFUfHIpfcSEdwCjhr9EJh
XSDny3sI34WUg9VNV2aNprnjg94R+/CZQ63NwyV5buKoJeHcrCds0sGqbLnClNfO
LCAKuRZrMONNIABVeWg8S6jNrru/FD8Cl4lunkk2lR9w+DY6Gg2D7djlj7rMxGq+
s9gcQEdrKmFANW3Yqnw9FHX/GDrvwSAguE1npm/4O9MbyXyWJDmJDPZ0pmJ7y1fG
GT6xPT2fyMFTXrsoCNC2f2jGRfMH8pHF+DapBp+u5Lue6Hu0OeIbwESCU1Jw/Uai
1VLaeRMewLaiUF1p9nMpp8NsuU8iik+aJWwoZgHN7zwJPapQRdktw1j+Nbojgh4n
7GLcxpKhL8UjTzINjG3CmTojYLH2FGFdRR9AoOcifwpALYeVlyz1lEq4n7IR4B7T
x3vUknweIABwXiebEkrXjOv8jdDvPTHx/d7IPxiNkgr13PH11T2lt9ZSwN1T8eum
/oos8di3EZnD+W70pu/Yt2vhy3whopSOyt3TmvtB+uJ3CUDsnh+zEfxpaW1SFbFg
hMhPF7mGmO33rmvdNVpUNdasdbcrMQyC8YHic55MqXP3lZjzZqEvrJIKEJNn3Dft
OkZCeZocEIHFxbmMLGq70GaPOFyyr8Dlk9K1XWo24hCusL46NB6bqb1gl7w7jvhp
yHBJ3jq2pBfIOS3n1tkT2QJYjnRVoTNk/l6SJpFvts4KL1Y4hAMCqdc0d25c632K
KdGSnTXJaTJsxiSMQf67cTa7LoBrigdODykWT5xsu2QSR79pq45i4ftpepn3Pq5J
L/32PEUNG8nPYwiovfOFXLXpSWT3kHqndtGJRJLOaxFCdmZGnFfltz2nt6xDKCJM
DfCJaV9qOnJrE0jrJki6U6DndR/bk01dP+YqqJ1WHT1F8zuikz3kbe72jXRod+6d
trsFzaTHk9hWHs6uZ7eh9mlAj0r0RIa2s6AM5AiUKJrMTmGlpGeqd4MwzzChXEjh
3g6CgXY83eO2WVa6UYz289KFQwzQ2xqn50+EcAfAtVRCjVaEX7DFBec1w+fYQQmB
tLhaceZ6UeEEUhIM40XTbvEs7NCwqErqtGi2j3ZA8J/vCnC6XhtfUU+MttVVkB8o
6TxKiqaP2GJk+SPO5oLB4AfuCMPjwaiCQ1ICdlH1DD11OZMKzSizt9tdKaNnZ+AV
e7pkUexqQcoKxue8TxBKHbCQ40dBEwrB7cvqT68u81ybJbO+vjabJ0eAK6At2cpa
Bjc412p9hBLu92BkW1YGNGb0mmhMOUGcyyYbfLPb+LWVX8sL2cUTTKRIt7Jk4jQQ
QvER5ypphKd4SM8BnLoM95lnT3h5PIjjHYne7lBmPneR0OPciVDzmy0nUPPire1O
rN/chT77CpUyo9lnJEgR6EF0yQz3eIUXIGi9FS1Z0y+OuhA2jtJG9c78P6YINvik
NYBlcSBPmWccp+s7IsX4Bo2ymn8HLWLnQGNv1iLjlQ6KL+pMhBUqdANaxrYfkxMV
I362znPzlc3So1Z8lqnWhEu2r/iiL8HjfPlddqb4YHhvBfG7TovAGB1LYfJyYcnR
8o6g1bumqKQOwPdptS028zdvf8Opcx750MGm2/cQHDZK33P64cjVTgVBAsDnYrxg
j/s0h0ywaX5UbJEkDLqaLGj34qHp6tOzRB0Fz8man1zVDjtbgBHhDPPAMgPPEvZu
vQ4MUKTpsEe7MjzCjhVd6Qu7ul+nVpFqnlKtF8dI+5oqZWLbqmwNKw8Hyoif4BQW
uatkI5NQWXRsTCn8AE9270Jj18mfV1izQSRDOZsxiAMRAuwMokAsCwB6BK0kRB2j
1GE00AT79nTM/o2oHhTRIOtBvZZ2hKcrWkgV3tqpYGGuAJwp6MtoJegVtmSDtMfW
3oCK1i8hR8nocqPdokiTffHLmm4c4OsAhnWlaNyeJrkWfR0DcxfV+tBq7Qi8WWmu
1tLQBbpD7jIujeRjEpBXnm4KFgsWveOjR3V7rrI6OBcGcpC3XT9eRxK0ngi/jVy1
fEbpZL+1+UvAZpCJ7wDUunUxYSxYM12sybXwEuYXqGjaaXTl9jFehhcvVLKFdDOj
PB2Ekkg7+xkKqLQ9xi39STsjX6olDgCNVOUydZ4F8sdoWEwB1CcGL6caKYYXcbhw
CRPpQTQPioQZ3dokP2N6Sl1HT8jqeRHbGe/LuAoH4tsay8WuJAUkg2NPzOCV33Su
Es+qlwxXRhLwZNZBJKOBXXXBiDlmJ+OJYTItjxCmtQt0BLS13VRxWWXZ3fFJ2aH5
ztlLinUaODVfhOOWoeOZM0xCAFRa9u1SLAAnIRgDEjEerp0z89aEOjf7qDW7/OU6
hJ4HOQ4IM7Xy2WVBHV21HUI1MZZYX4BV6wqPPs1Hh5aPi06wu23Q6VIrY1VrX0vu
fLeZlGL5leNNAYsgwvjLKqSvadKft0vXYEw74qJhh1sUrQ8f5chZfbLRzu/xV30z
0FBu4s1cmhrMmQRR2iLPaK/8zPUcjyo3ZHtYbzilpK+SgcmOU0Y9T7PEaQowNgyF
9Ng4/G2Tov3aNeHc/N2x/Lq4jFJ5QLj5TETIc+g7bsH8ndp1/fZ0lTtRuOOKM429
lqzZNsEJZneHp7SqBQ+svjcsggnUkkYm8rKLzQtxUKTQtCwnkY6VYH9zuZwqWN1Y
kdBwsDXhkcHs1Xr2TkL/xYuwcCSgJEr57yh80Wtnwjj5oAtHLIR6l8y1WkKQJons
nvoKIAP0Fo7MHVAQ84VhLPJATt4w7PkA6ZjLTrkLZn5xC8rUyCJojkzzQvGbHp4K
6JlpAcbkr6C88BRYo60/VRXgEQ2e4lu8wMF5OHQuPLa4gv0zMZNSgJjBFYCZ84Wh
z4zf8E26aAeVLZWon2wpxFTWTNpf1qkQurtq4K7nY0PEs6nwIGt5v3C+on/WlvoV
P5RzoBr/ldz8wwsydIp+75dWDy98rMtxtcDKJ94DQo0C1rIojKEBnijwfMBf9BuF
24Hjwdfa6Gf/BMZMOwCMnnriNXFJlaYxRRqQn3UGGJvaGsquqO0Wvk1yULifGpu7
KC2VgZYeMrnZIn4J5h3oyyekBrUjgiKqRkG32i18J6yo/H2tBaToq6myR1L67Yhy
qBAv9Zc0k+o1kPEbf1o6hKhTNmTYQ/ePiY1skaO4VmCOT9Ee53fs3bPlCgq/eKqy
XkELw1M8OM8Jbjfwc/wBsXqe97qpOlqgvf8NfO3Bvh6G02FS/9aYU1ekQ7o4fhuE
imBUcTz2/AELjIsI8KBMc+NTdUaC30v+Qyt3lHaapLr8zxOKdQV/BQXwReF45WWb
WvP5I0KnZu5xa/RgviXlY2umCzdrDkIXu1jaCBAxRPPBjEtvJ84k998YOfBEf0hX
jqA/uBr6Qj6vQVD5YaIvLKreCH4/i6fEzxdA7TQZHcoQZDWMKICyXSbXBz2LlK2o
u75gerId7Ws+yxu9nluxZrksYepBVmGCfvV0cXZ3D2XA0hl8uE/YlZA7Hke6ip79
Z7hvjdtoXcFJfAReDeQ2ah+d0kzi6qS6beQvAf3HxBwh0qrwxUrjUdz/hEmrn3si
BFWaigZeVqloonHyLXwn5scKI42aJTXMsJTI+r9nLTm+M7+kCRPt9ng/KioxnoGt
cTPDaltx5RsWWzk4ZoC7sY1rYdH18Za7btcBTTgpKt3JVxMxJg98eTI10LOBQLkn
nu0gGMHXb9PquxxiMWKpoMm+Q2nr3XDCNYRm72aXyoRZL9gRBfDnJo4zwu3JJ7dK
xrGuAYvvtMCklzmjZcVFdgMKU5oYLu8k7o/oHzIbZAuobT7k9dxn5BQdfPPfntI4
VqmEl/nhx26fFkcGM5YX+l5xn4knttWvhM0823gceNvjax6UmX+gSzfmshkn+oiE
Z+2TyUPYZYgFLSiObuWk8J4j3D4zTDQmIqUG9VAwzhiGqUc8r/nQUpNIPgJQMkJm
PYv+uG0KgiVlqcGet0FaM1YjkLtwtAMVxDQwMaiw3IMg0RrQ+8LkIDuKWRlnvRBL
DLPZ4C4BvMv+E+sO20v0bsNLW49CshXkj2lBrg77Dudv3Lz2j98PvP41IAGZO5xW
gDXbz1gIz7uinXDoiiW+N8vBvqnRJ1j1NgMkhYNJfghxOFAs0rF2s2er5TYtjICS
SdAaTwaSESwFcH8QdMUHLw+uL3wHHjDmNck6Pqr+6GZ8Eq5omtj+2B59lSnAhrMz
+AkKI78QhktfUsvOh+FgY+Ih2C3njMFoaKEUR01XxV/ABgpXGSjctLV5ZyROEaD7
R+XMHUiyXANkICu5FN0g3exkRnMOwZmsmdB1MCAHgCpA7A4aG9GuYK6cuiAiQ+eI
OJxb4S+R6ASr5V+/IklSsfRvUC5IcNViaxF/ZyFXI8tsTamDHgwfgehyKsRaoLIW
xSMiwm8/ub5gfzM48UbZWFCIdTS9jlHRxRZNR7Xiuc2rNku0a4RmzIQ3tPIsE5iM
jWbVuAxGkZe7nrUTlipOyDdM5uE66DLuFKWup06bfxDY0N2zmH0iMBzUGsykAFRx
RVlopV5REDdSIgu9Sg/Fe6jgDpVaxdRVWGHAFPX52dvgUu0f9VHAyr6iBeJew2KF
a+IlJPMF3wj0c3Lz3JfnjHA7+EwNifo31MzcdWfRzp5NBfaKcdaFRqgC6DMuR/eA
8HfiWQg4+jtEsX6rINhw6+9vEwHMjU+OAO9qO+cSOXjskIjSkxGHwnwxoB2nguyh
1RkEAfvPKGqALPtCMR9RUAk8qB0QZn+Of9Ntl2mXVL7bkURK7hXhB82SaqlUx8nF
wBfxt1oYI9zms4KUSsA8xK/wyquWN38tD9fZzRvBgiZPq6CqFCTVN7S7LSYe1XTw
iQ4hjndH5p4TrEojq22VkVPPJC2o0DEQdZj+rPwNc90JdN5Lj2QQX3LBUun5VYuF
zAQCDgsM+pHl2GVaQ9836lvIscMDFmCFPtFJFgXSC9GzKx6Fku6rYIHqDwrXiiLS
TOMbkj88eK74v3vUJDxTGT6HbSqJwb84omwClQjAYchyPR3rEhQoTAvxoFmynqH5
M6gdLWD4TxIm2cskvG4TAFpNUgoOEldYw/r4zVY7vr7IzCriyXJ0A2VXeDfVIe7i
YubyZM4RXwWYQ6aG81jhYqSM+pjHmL4Gf2f5j4MZ3MNfPej4UGVYUCtNzOB1VhNm
Jj2KZ0A09kjSAkRWqcOlU8LxfAlMdNbY/T0aO5X5og+j2+i5FZsKcLx5tkscOyQs
4OQQ6RiNf7FsbmijNMDAwFkXXuHZCD1p2y+8QdzwQsD0AO/tggsavG6j6T3FTbOj
u029RSHl6fR2L8ptMs5KVM59wv/BZX9M7M4rcDLn9KOUscuhFwMyAPi1dT/CI0pJ
IhNURoqKwgrLzeq8ojfbKR2eW6o+2h2lKQDBwZZuSM3Wz5zFngeE66ZL49oxopUA
bA+/MUnDOkeOpLdb093XyjxfTgbgvNWOMrj5vbrRb2zyri9q+wKmIXgTGqXZm8fo
IMQvhJFAlgvjV8EfgkDuB+st/gtNksdJrNKsZU5RO6rKSsyzrqzzLk2LbOn1cg8r
SiAqZUazcIHvMC3XWujJ1EdXR8BR49BYrodUmMwVRvJsaUIXMi1boqPKiHxPgliJ
b3SL6qYMrj8sLwm+rEo0TLvnxfxl1KBvx1IfDx0cgCHMa/Rslvvr9AF2bJBvqiqt
A8Q/wfdW5j3D8RJntge3kQiVfO9H41g1lU32cjbXUOkCcjnOe6DkqTdKdwyuMOpp
PsyYcs2Ve8sT15gFhL9KQ7AfOJZEJLZKmxsz1pumrRthTS2CCwo/qx38GAC0LYbP
ltQIRuDWF4NsOtgsACcQnrF8b5eLBAtypaxJ+pRPKhxiaXwWjJ0KRpnb19Rlt3lZ
YZXcAV1zQ1Cc42nxl7+FqcJS6Y1qAwmz+CYUyK96+A4oHNk0DqIWx2C+8Lv+52F0
0lUsOwBfeBWn5GjGWPEakFNw+m70ilueJYBVwhT2eF7dhSg0ucHUa7aoIrbbWaDb
RdTmQx7BcORUm6iSQRGXnWdaOZeOgyhWhGTzQWJ8vnGWsy2OhBDuIULkDAx+mDN2
0oCN8ydTjRy23AS441xXPvNNJsOpAFCUGnptfvd4gpul3Mxqr3CwGuAnDDVwoQp2
sbumAQ/GoxGlSmobU4G8fiWk30AC60k3K7Zf0rjzAC5SBaVoQ6ti/l5+EthLihLA
BvQQ4btkYoG5xbrcHpKTbo4LYce1A089maPWvN4jTHNefse8bPd36CeKuOUlBFyx
uSQCzGClXnMe6lP3tXZpZ0B1skzKOwiW09Tx2ClI6mGdUozhoRo+UJGmHm4KRXDG
0bwJyYCbZ1CiYHsLTD8GkJ20g1dwjbzbBs2T3MtBMksPpjHGj61Y8jlAKhVquHud
2UKLo5xpZSlyi3YBHSFJZCrPzilQK7IDIeeSHW52TgvbriRwIPCYai7NPKxvvo1B
l+T3TOHhv4DY9hwMx98uqjvRjEXPrbLvid8Doi6AQf8ryfMyBYPL586aPm5tk86A
ZyMeG3qPJyfP4KP6yZZxCIXT4UkKbqHsKZxFMwT9pvZXi+oCwBNZRS4+BqCiZXlz
TGxgRIx1xQVQdn42yOl75faizu0xHGJBjjcpGlkKXshGCjLScAkmwKKuDaWvDeLo
PPsN4zNKEkH/cqr5loXVVKxRTNMiVhqE57jrbK4reSHCgCkGQBJNk3+Rk17cUlkF
+IKXWnlnNlcp3TiTH+zrwMdfVKroGUTIh6jIZgmhBfnLPXUc/HMLVCxw8Y/9Fnbr
gGlaz6pJPrC31w3PQRPTcJmRtvipD8eg1uCU/dieGCaxQCjfvr0t86xU2z8q9ypf
InsHUAF9g/Nud0aBko/dV3mqBGDEhcKVidSFdQIWA5AzXjx2yqecyCFNrmSrnq/1
RJuEsvY14tSnhm8xbrEqplri1PionLCfVvCuhzkfZlRfKuegCDFvk89zCPgAxb0O
HGY3Luiu49e0eLPrEe8O85hDz7FdYWz/NDi/VX2a5XiKnr7HpUwe3Ek/f/GsUk8a
w9gGXvX8Y0QCLM0wszGHrScCBQ5FOnuCNuu6IXEQQd1NlBsDs2QoZYG4mz3e6onJ
rVxKbVW5TBI+5L0EsyN8q5hi8/RVIj6pt6mKwYnRmbmfuwdd10Woc68IZx44hpi8
N7BFcXn9PJxRPQouYCNXaIzOyP+wUg1kGGwHidVwRfWCebRe4Q4K2EJhzG5ltAw+
rY6LpiXc6hfZgbplt/YC7Ri3m0twuYZD4PWY8VV7yhMJxrrQlYllsBQvoyd0MWRN
1pw1uoVIqhugc94+Q3JGzPcnM5Jpndhfw5t1+MgHtfDeaJmQqKsBUYnsKPisJiIP
JJWgIOT7QCZBLp4mpYH+yxv6X0V0LkPuLCT6cXXCi+yMTnv6dpqbMIXyAM2nzULB
Olaby3pok6KTKOB/a26i8HtG6Yo5wWm/JDt7sZEX4hBCFrgwq3SYYpoDBWn1RawX
jbBhjtpJyVHpbbk+2yqQKo0AORucM4G/bw16Y5ZNKVjbdxfBqym397Tt20GI3Ft1
HWsljKUGE17Txp9EzluXTokEuQ8PnUKgQmh0UDVXk18Gg2KLZWIE5GXD0P1sAjMx
9SO/r9tsCmAgas8o/pAO/ReMUMi1TeRhUG7dU6MWIwKLKH+iOM42XeFsoP1GSXcd
srP+pEUylrFWCJok3MPTyqYaEPhQMRWENL2SFIFz1XW0TVeLxq76lur/OY1fA9SR
F6s0hoaRgnPbp0T8vJLbU7tWfGeEcT5/OThqQEDd7HWchlNfW7nJQxNTWi2h/hyL
5UaUU/KXgiOurnbUBj6VMH4Kasn2Rd+wu71+6gA2qqhaSM2vQA8a85HG/nWKgxzf
Wm3ZsbBZ0kIWEI9XA9kZ8hHeaqScr9CXiV+d2DJ+2Zsu4Uugx295A8QcHnZJiK9B
9aQe0aRxO7wH27YaLzzu9ZrFo08LDs2+r46Gz2mRkn1qRxNp3j/bOJVtmSSibynS
zKlJVsAEiHDeUiqkIHn15uuBrXrtSg6jSM7k1B2wE0YvPHYia8NVvUlJOxfzGtsx
FSGlfN75KxPIzJl3o3xv413y4aNbD6x+n0WSETYng6XWNT5Efhi6qymhnIivCYCH
zETkFi3voC3YQ7NEWamrmYxS1kIg7QlqBd5fkWg+KCJ8AJUCW7iRc8GUd2bWHzdW
1lE+stA0CA7YRa/bhorP67NSxTcBnNh/pb2+Ke2HM5oHRaTnVbA2tP/lNdxglldW
xkLpyxZ0Dk38L300fwu5R0wKNGi7aULxZtkBzdtYKKj0TDf5FcylRKOZh4BdFCA/
bD9dfk0Q35jFGDhwEnDc9eATOexjlMJvyxvvXeLvxZk5HQVLkztQQn4MVZChxbmZ
t2BUxtHOZ3CszwKNlkdmnoCZW77tBLd00ZbhcHiW8XbkeCMUvjuFkAcCtQjKExok
owUpi2AYbca9Oc+mKjZToKeLh7DBv0B1zR3I7LO8Od2Ye8BR1aYjpnrVbhKyxF9w
npCjDwLq04UgjjncdM1WeyeqvavLntoQK8Slba7fzIZFmUZnuqGs4kTDjYaxxxn4
dEMCqTOS7buY5shiQvS4Di7lrBsCxnjUu4xEBsa2WCpDqUU9iYaLwz9Tv5aV2YTf
or9kb1pjFqybs/5PB1j6Qz5IFXQa/OjOdhYpZnCCKQHx8OE949eO4DDz8RR+51hy
p+bmwrDxAVRZE+EL3Pu2Wwb4o7r9wVPqoOk+TlMgbXyT/LoQGG0QVewVcQTMfJvy
UDurabgPNINdfz0JGB9cSRvRNHTFYxL4ruNs9JJD7WkuAn+7KDivDbbZJZpE3mUr
akn2lzL+Hh9gCkFEXVf/E2z/8N9k23DXohS4w8LE3130H/AYgJc8+kQKraLZelYr
LQloLofxg5+/+LTu56ageLO/5ovOEzycRapc8Yg/gTZw/aL8Z3KnAeeIqvomdM5S
nOiXld88ffx63pk+6DVi7pmBeStlwyXMdStn7Y4MCWS0LaTKeAfoBw4+BP96Z1AI
2nByhEagd+DAMc5sP2UK+P5hvfuCBo8JatOindXkTFEZWi0+7ZaBn6PfqhY7nEbw
slXTk1CPlEG0kuj+sKfpm1Ebz6edhqxF8uW9qja7CNd5waNdhyo49RbvNWjJ056x
B4z3ER2dsQJcFvwSu2B+BtJX/iSwdCKDQi68cHEqwrP4c2gwvdevE2CcXd5dBA7G
Of5SHKTidUSK6KlroBPXKFW+6RoqVYDr4h/AKoMBiERKHJs8NV5SRYCVFgCRD+Sq
+n32UxkXxsGK2WcRkgduFTE9KXGKD2wNg3swh9K3oFCUiBDvSaKKoHfUkDhlraOb
pB9sC7H7iuHyD3Ny/Ob+ScxlpQcNUgjbxkR0wSf3hHc1rZl+xquPLJCf7bloObKm
9wAnRwDsS+NAFAHDwBVJiFb6Uh/oeEBU08OexHiqKVifEm7EncYpKeaA8niysGKQ
zyWJRnagl1/sUNVt4KAp2r4/U5f6p4pXrZKPAh8XX1l3NbnVBwDqwrl/yEXhcBZW
xjWhzsZt7xJfaJ2yKdDUWC97ilkdN2vB8aHrdj5i8vkXwLisl9hXtsSVhjLyCh+S
SVvr2EdK6JP5jCZOuUMdF8WKPQezSD4Zoq0YYFHe3amH1+f3ul9Xpj0n+hf5z5p8
MTsPwHOKpEhg6K1M8L1Y9f/YA4ulV70ATkWDKZ9QGjSPAfRUqvu75JhLwxKsw/MZ
CnTTCDW2y/nJyaX4wQJrdfpqsPioSm6j5gwPKmRYn/b9nhs/U1uR0iX7ghdjHORk
g1mBHl4e6UGFgH56E4GVTuhFFv5u+8kG7YJ5eHTAYlhowuyeGyP9Q9nH8AMmUWvR
d12qSnov0Bd1xtVBB1U7pbDABasLFil3D1aT6ZYKnuj+M80haglRVzXHIvlV112L
gI0S5WLOpBN9MzF1Y40+Ar6vpcGD6oExT4Ojhlkjjzio0BX87Kzk8VDEY/F2TAbz
dQ0kXLnJIyS/3L2/jkzkYez5s9ox9yNIbfMxxDvpavPjP40X8L+/DUyXOd1PgiT5
qJ1HAEwrHcAnl0sig9RdFA9KQqkSMAS+QX8/QOFZmAATLetCzMG/Ih0GmQPWWnn7
bx/QA9KWFFNekQ+mcgyxOxUuYgSjUMfTB7f484FCJ3zdCltuiGr+Tt5aK8Z0iSCM
5RWcZWUF2yCBRNtZaPvKqE5yMOG5j8u9JDPNOVG0cteF8Y6698Th99vXKwUFiqfQ
7NKerRZJPpht7xcA1rwEzIF4S6gQc/nUUp4srWWx75lrXVF+EznR/SIb3NMy5uuW
3QJRi2h4t3dAtIxCTz5mG4izKaPY72wNvMXvrg67AnIyWKkdnGF5eWjb1gRGsMwc
j/JgosfB+kKZIaXO/qgxCkynbjut70VkrtS8Jj0n30aGsYc0454W494mN3uEhNIZ
+rnTi1OWjNizpPAJFs1N7pX7kuQtrVxVSns3uZAmVtGjxCaMfoXhu2o0oLEbYw3X
qbTnst87TQndf6648fb1uZRuNuVGMp4YBeu6VhqSZMtKtirGyNGLLQUlZHVKweKN
0J4rn7c0FMUrXvZp+vsh0+XU5RCNZj6TdQ5uCAjrmjzH1pbnZz176BsOGg+H5Jvy
er0eZSk4qXDqQMckMc1SpIy6Lkump+nMKE58Nzj2qVnw1GJlaw63Hu4SCT424+mp
VQNb/6FMr5hd2HsoaD3qHy9lWXENbzF1q9z2wX3dV85Y9YADWFju6LYf3CEQC4kg
Jc4ENWK2iQo9CDn30C1Q/LXNqHey/7b/fZIaoiawjYbwunbcybPsduw/IHghDBpf
ZHQFJe2oxDYmhgoF4y327xWBzqG74dJzi50symsrNQrsx8Kn95qWaf+bC3KNrfPd
VOQttdVIS+rn0VIVuspqOVgJB4Di7sBKr+z/7Hc4S41fj+JnWxqJZd1jE0pvcMQ5
4fxzcDL2Hy1ui2Yl2WHZ1H2YqtibCCD3N0hm6FLDYxYZhWTKZ6XpJNEcbs22wSl3
hPQGPlzpe5htDrrZpTqsKB376axk21MmyfThvR8eB1+6p9wUxe5NE+8W/n+yKJxt
WSAVYcUBkEKbL6qSWjm9MhAmNZQVY8V1wDoZK2btJXV2z7ZmXB0MAaZwuiqi38Jn
tCCRS8Ft8SqeztiTYkNKi8u9YVdLGAHO3aobDZGq9tlplMS9ZJ2QWeb5PcnnZ+VP
/8nwXQOamjiW1NGdacC+GEdxrkaB4iuGRFiqwA3UkVhMbBWLnvV3HDoowIevqLz3
Ww4V+VuiAO0Ch9tZuO/H88HDoH8DI8fsFLACEYp4q/wOvnZfjk59LMp6qXVJWrvv
ClxGX6lu8PGQ2K9f6rdBYOolmmaINYB8kULy0ecVJxkjj+fCHjBUiHn7LCsCcxmX
Sgf7lDh+IeP8weHbwvjw/0Sr2XLQGc4Nkgxt4m8gmVtkJ0irI23EhVUWiXyJlXwi
XKb3ft1klNtnOgFaFrHr9jR3cajTs2Et3O0jUhVJVd+u8Wr0kKmdrMFUwYdjP00w
PilhONDXQU8wA6h81yYHM6GPCiTXfB5gnwdt2ICnW4aOkcD006SDCUTLtMo+o7EE
8y6+jXvcwSMTbwArAp7FOapYeaBD4VqgfVEsPlOA/cVTkfEpxBLS8OzElvngwjoO
UiO7Wgac82aW51JplUc3tbcfNNKPw0NcnOVek05h4gYmYvTFAJ29L7xjDQzjnxe3
oEEaXCogLtEx+kLugG+Eusynkzy4gHNaJpcrJTQgHnkX5xrDZZp4uEkV0DfO5QMB
Q2fBNMsRLvXfNQpvhqej0TVWKHMosX8+1Y1UBOH07cp7OknP/XchO2AUPQjahop/
+gBfskmVimAc4841oV+xMgSNC/n+4LwjEOoSWIqYhL1t3jtv395IaJcj1JHm6g28
pmJSVZvON59aFYScGKXJ8AVd84G1IlMGUXaWsO5IZGFDKQFnbBjkvW7SinKBvVRv
FRmV1hHrs2bBKt9fxMo5Zhp6LQPUqDOBT8yhzy5B1rJxJD6HpyvCspzn1cRSu7Ot
KjFNIVJvxD4Rt+3LAAKN7lueTHj76qB2Jys2FzfqqDNV/b3cyCcRFlueuX8UUcUh
hbUyP6j2mnIqFtsZbNkOvQjxLKCsOX1hUiBWAC4IH37GhbRaB/y1yp1RvsoAgaCe
jbrISUp43k2fgIiN4bhJ50UKU5HqY+uzYk/IsZyFCAD1WXtQMX8fCMglt1mt53zI
DL20qYeQm+tBx+3qituwr60cjaKjFz9ORoUXvfXAOFZ5hedFot6fSqm3rLnfD7ZA
mNGKe9p0Bkj1lxuGEQWAMyzUxQBlo2XegG0tw6TkUZPFxz6QiV5Ayrp3HMqEfxpL
32tc7KuOHbqT7O4zTOaBXhrBGGQGYwx22GLBr7lT0K1EtAt79FJKLbNfeU50w6Bh
kYmCvFAutvhGfMklXxXuqV5LbmGUwUeVxiOW4EarPVq1c7MUC+2RZnh+l/GRHRK9
tV/RZFY1hMO/FpEocAm7WQyVd91+xOIZZj8t9vWP1cHSolYCGhoJftp36LQq9Zd8
zeclO69UO9QjAgw6htUJMcbuRIih1+jghvqtiJ8ct87Mil0mzbEfp5pU3mgjKGbq
8TXqsPEICxY8KmfDTw+0zSQ8hMXDnSj3M4EXgpq8X48ZnppVjn9NofMOhsxArnCT
Gg1bbFW2dWqHU7VI/diFyojHqe8ug2SdhcGW9B5C9YzV9GuDBiVTvjaLSnITBeX9
zntVh71r3raWAIimclrdGZmduiU3+1y6bw06V3bNiSZqqshKjOWhKnVI5WcwH+5r
yZE0pmU2V+czCZoMcEApl0j3rvJ6zTL2XU9CuY2/Ew/NiF6KTFnceKJiw5b+2OyZ
t/9J06/oqyGj5pjAXzP0rg30A6g3j2p1mQJMHnlTRqwEtWlw/a4OUegYz7+7exCj
dX7jRAJMehySSeDBV5nHKpq9gTtsVtQ+CqaLGWWhoONb1gqy97jq6Rr57OrgJh64
5WEYrjSO8GBWHCB6cKbgUE3uq1P6VKkLTiEd0XOcqVwHFOzY7BWT8YyW5+Xjzewq
vL4EhGxU5ACf5RE69whYB0c3ExvBSoLXkk31EI7KdIPJrAMjnymrOTTZ4zCTFy4U
HKIHwkXBUgBy8krODG7OdmMbqeQhR7ScUeomNUsjbsB3kmpfCDHPc4cmimunac2M
2RRcbvNURuuuErPVBAPoFJ9RJSKmQ1jjz4Nb2xwZjlhxGQCtlVkzVKfutzsLo9xT
17Q+OOueZjSvHrKImFN+Lt/aBNAcf6ho8KpGrK+CplxZeFnxsmwDgVsJKH0V7f9a
fqDqIa+B/OmhycvkBlEOXOCnfqxvXYwApskUh52zLHJSfnkqDqCBXcehI+UGIhXf
Tj9No9V7PqoXMWbde1f083cdLPk+5Gb3OAw2HTu+AbLjG2Q6CtP47pt3E8LGtJd9
hBxQTRCdJ7k9TL/ZfGVzIkB5oqwqXwmOCZVqjx9o018nxJ3tpAjj4b/idR3+wo1s
HQA0DJQXlogUKV7PBZ1Ofvad/eEjowi87pBQa+LR8Upz93l3Tnd9RyWksicH6Pfj
lnWjctomNEJ/TElz0JfliPTEWTxNseC7gb18xP1uOekNlxtJt4RXcqboqwL1hRcl
eTznuR1QwICRWy3oZduVFhU6ZvRodjSXNcKyg4SQPNfPnT76AAGAT1vasgAFA0ov
WQbWEIo/I39WrtSvw94s9OPL5pNS3rpbRtlCa9/vi23HmBPV56tyxRpHAKFc723q
qfJ1iJkKoOg4a1T7ZuieeT5oeAiiezsnkKnL/ek05zungN+ZAHfkblsNpqn93DK6
OOFEmgKimm+ZkqK9Tq3DWBfcZi4QtZxcGd0gBcYQgfVAxNLmnJ9gHJwJbt2j/Qy7
UnxHtLMC+C03y7Kj82xC8P+oUSF0p0J6HGHL56Cv6WQVGK4AHG8zH1eKdj5fQORV
obZGxlGbdIPhGmAQEZZBnhOl7v3LW3OzHUrUKLc5gbg46cECtTMHRT0nUGQNHaTs
ChPT7F6mKsSs+AiVd0vptVNDDUdRlrPdDU/gFBePAVI8jouS+rh6t5Qa9B5/FFS/
WmfggciCg+jeQzBZiYW0y55rS26viDLiKfHe8QRvKRDcgc1SoTFahf3IHxqzeB5h
tn5EnJYEY3GgsagsJnxxcouodcsjgBwIZpi+K18VeMn5/SRn17JVj9W3YHDqREwY
iNVEalK4SMc/eknIDbwBrmjqIhvI5bQQ9i9DIhrTUQlbAk9O1spXzxwMkdfPaPS+
bM6ZgS+0hKU+ai+4uTEbn5AaTcVpDSgeclw1MKVRN1nzngLsLtX3FqQb77QnFF4H
7CXEM+rwNpPelOWIz/GCf2tujBbSu8Ke2KhF3AyxdEChmX+KEERIU0A20tPGvF5k
pX0VfMY2kAZmca8/94nztslcj5lRmrxDfqTbcznDTGgx3wDn/E3l8q3sAwqNQz0K
K3F2gaCYFngoXMhT5VclnXzUcEuEdttVKkDHZ9RLErL+dWfTQ5XY3RxR7waxr2Qc
h2zBv4XIs8gIbbGWf1hMI+AL6dQmaXEaWqxPV/S70o4ku4JnFoYSGEwuGrStAyvF
2T2l3Ne3lZeZ1SgAL/Yn5jvpfgB/L1YYnkNaePoEyX28VJX0cG1nF2F139HvUrxo
wD9KD6nUL+jrLyqXgmvToKuV8owbqx4xDJEVU+zNWgdhPfn1VJiF6LChLU+KG8ar
3PxSP+QQHvGiF5S94rpXyeePCIMlL+U4fLEB7AEAgB6LXAgjDeOdG9BCFYx/Oxp9
BYBss7AFv/+AoO1nbJXpGhurI0a2ABB+7+zBl6Nnp5ldmCidl5uTRGckfQmLkGK7
Oh0YDrNEu+HerQrepKZJTH8/nhBnlNbWCaAVH+XkV2ly8OddUQJvz44dYh8yWcPl
IGfBkgubSPP5XsXdy5pxTEbj839i7TXRPXEKkpGTDInolGUEQxZ8EBgaGVqlEFfz
OZh1T9BbvTiU88GIy+A8XDzM7dgcEgw/uFE1XqWHU8YHGH6iZ3fozKvdfr6hoXIi
YvRme3oY6bVdjApFYNm/UROtDtkDclK+FBlWwPo6HM5hCUjXPiXTNT2R+jLOckD/
mWMnmNpa9Jsm2qMedoFtFj21DnkLH0nmkT/3Djh6OZ5Ivt6QBWy2r1yZk8FKhXlJ
qnMhjmYy2iHMXA6FpKEoNgeofcOSz1GYe3mVWqqRv4pLuO39FQgr8vn9ljUsZlCp
jUK2Ig04Rvn8+gicynduau+KcvZzseVVEMY+9o1iAawr7naZWinBWLCXBtEoP7yF
pRDZ8r0ARP3zGNWjBE942E4KS/R8Ejwyt6p7LYuHP9RiZ63XyN74MgAJZBgvdiQC
wIkmsXyZSOScKWUShZ9rPvhMQJ6qr3ANCxmvyTM8XwQ1IYFaYC4ySfdPZCvMtEEU
/8+1ZNp0ldfCweIY0B3VibvHHWzvGjpDV2HK4wsmIUlBJJFPQtmQzLI2x6WlWPeZ
0BSEhY6hK4ERsoIo8aExWLtcTH3hchCeX/YW90BhaJnFdIDffORmO/6HYgyr3eCR
KwruuNFYNuhy6JuP2vRZJihE7aVqiv7JHWSBdfBqb+PYhvQv9D2nFCJfTqdAay+f
r10Va0CBuauxML9lh0HxszprlQT56uyAeQ89oWKLeBMmz2ZBQWCTemjILGe83PIC
xAtgZ9s8x/KioEjSB9xb5cKg+Em2pPMcwnbGcEOT/yLTML5abow5Fafcz8xj6pwK
qLxQwUzhMkLe4f8G22mPX9lMBWl82iO4JNVEp+0zrFtLwPJgBIwYnRmPd5lbrkx0
zQqTVCv6BzQcTT2XM4VtTPhShdM5d8oK+gfMF/zusfcDvvt433G8McFnoSe6vVYN
AV3bQH0MJuceJ/W5Hm1IsOFzG8/bfpXq6WVBiB+jhFk4B9FDXO/CeO8W9hTtfffN
atpESbHIetlF/H1bwxBcoDMBL1R8UMManEaU1sm5IDw6DA6aTYf2ULo44hcWJ2l9
9HgPFq4/2UUY8KPmlIJxe8flZ9Zb9Lu7dSGWaizCbtZ1DPXFjAFriAzpU1XwQbZ+
Ly2BxYWBaANYR/61NT4mIQUAMJ2bLhm/EeIec++4efdZdzMYxjLoHUroG0rl3b3U
dE5k2aRt2Ej8ZfTR6U48M2gD3dM6JWC3E2LG2heg9g3ssHXAkJWiW4ul/E8Ik/Q7
l52m3BvOU/QLh3r8f9AVm+rtKuqiWALAtN7o/IRGmzSn5oolLjIfKUZlSLB0n//P
bOZ8URWsxLv4jHo1LGGiu5kbkBbZL6ZylU6h72xt1Hbw0my+blYDpaPnS5XrPKGS
MQ7BNwdoPfy6bYOiKiKifBekwu3oHK9n0Gf+6PkJkYWr0sP9GkUtPnw0HDZ65I2H
3Ot1vjVWHkMt4JXqS76WAI5ficCbpbvo8/9grBw8UDiDOshXG5n+3nhxExE+1bkR
QTUBkfn45jveHR1+9VhzCWo6/MnEpDEqVKHi3Im/lS49+hLoZ5cGTu21LKiu47dW
yY4CImFWmWzohc6hbaWMT0eC6xf9f9T+SAOoyzbtANyAQzawtHhSVYHVsrReeQNu
gG6z0zCNEVxYeDSErTtEUxmQs7xZkfjzJslclK2ooOnLly6vl1dXUP2VcySp//3F
zj04IcckwLcHzRH/ZgluJsLOQ+S/grMX11RdZcYNqQSM7oj9fPdtBytRAUPQMnj0
UpRu1Rzp2tgBh8PN++z9dXEc0lxTTKEMnkAb8eYA6rom+R7CVDdnsIgIheX6a2Ef
zhkzkf1tXyjtdFfZ7NxzlPbOPaTCoJFlKKbDBm7N8cYinvf4n/GvWN9Q/ml8S+mJ
3+MnDGkB84/b0CrEMOGQLoo0P8wJGI7K3wpSfjZKBNexQBMETnzmhFWU33AIoS/8
lNZwd4WSsLFky26zeAc8Czj1C7vaUwZkqF+ZkXE+wopxWt9NUUPAUGcrJKiiqbC4
2f23llBUObQxT8viyWzQQJftMOxb7EDY6LBXaCuvvm8ggpjXvx0Fnb9gtfroqHlB
KQzxgiCp5W6VuQQ+kpqJQk7xQfvKUQwjeWJRQBRre9GID0bfcbXWNKo6EbCL7jmm
HHrNNtYXjJxNyuWlMKTyVDEDq7fkEnMI3JUxQG+b+t1MmzaV48VkOdbg+pCLOKbv
zbOylyM/3Y0sgoyt2IU018oxOomJoQeeXJ3X8WWBTrEGDTLwCN61NcS1M3Q3dGyf
bMIiZ5kcfzCG35OCnyOYao3g2BIiwtbcQxT4a1nloO5ONnFp8qTRwyDy7bleqSrk
FTkAyUWZ8cptCD4NXRN7FIC+q+lNvWoYg+GYFgfCbjZeRJB3XPAuvNI1j0tPfODG
i0SH56H+z2a5ek1DlCx0dTqCBC++OB1yztx+MeIBYn85azWrAcJ2A+dBfZNiL4/H
xdkxGfgsckrttgI8gK4+RsjCWQf2M612C09N7JxKY3Ds47Z68kynQrtiywQHK5kt
e9Q5Cs/MKuqIQKE8U39xXdBqaR6B2Ibclr04KGKG5O3T5Ez7i26jPr+MHH1oucRq
AsV4V3h+wl8v3nOQ5RvDl50sZo6IUXtYL/RuxGHSpclWbUzIGVgPzeiQP5bBbKoy
5N82XE8SfaN7PqCAfmjjnFrMzd1gqHtB//IVXlBlqm9ruHTU0dDKQwcrH9pRi2za
6IjTEVZMemfT+c7Pv+mCSAh/9rDnWEOHoX/zqzUvvwARSs7Y5V4DzTSQYdNT1HyT
3ZX8plvUSOq/aNXKsVrxh7WqZOEYmrp2BhXDQ3qyrGqUOG5BGty6amgbxgUm6aTO
HqgoLiwUcl7eBy14UO6sVOJf0VrxQ7uo615YaXA9KkITL0SrkfWRKcSmv2cSWog0
lJ+6D85Y/5COLQ1tK4eqgANOAPmteHJoWjHHBweUUCksExQeASI35gMitnu7SecP
jiwqomS2ZsSMD9e9mvU7XUojNTkzK4MK8avuI3Z8arslYBfgXGjxl8QZM434yH74
VZ0uGRUnlS3+rKRAMPHH7DBmUDubDolexf7JsMDLH3DqQzhJzoJA3rbLl+ScH/eW
hgLW6GXOYnh8wYoGvCt9tPN6ePv7GGSi+Tf4rE2IrtT7ecUiWt3WD5hSPaoVZ+Ms
Q5svyS4eGf+5HvtOuVleVHKaAJkjBukazDy/wrbC1H5zavT8roc+Sa8n0389WqVZ
fiwy1g4nFbl1QsQoAVbSzEWJObsXJ4qRsQHaOabd6E9X0EjJn+WrZQE2UgHGhMWR
iyh1G3e9M9myCtkast/DHj30YEwNsPSnSQIQN9AJz0NO/M8ZuBRPqPPOQE3bm5u+
XCC7F6VDXXxV+65rC7XMX3rlRbg7Fr/H9MKay9zqxnFoxR9ziOYgKUE98pb8Jh+E
ORV5UhCnqSSs/7PY9AXemYREVFVvgffxZopjR4zBFyOWPclRBpsCE6wDbYp9x//s
dU0/DFhXdmEviVxQsxBYjghisBLefpKSquxRHEMUHJefsaYrsS5I8Qiu0tpF32nc
OicZy23SR4thfEuvxYtNRiWkfyCtGZRkjFyUpZ8jK3ndP5/ampyz0FpTTOyRFTYy
iDjzKBK6VahQ3w7FcXSoIEeUsAN0EzjRcAQyQUkjiLQmo8tun6LyTRAwrtspJE+P
3wdjaSk/0HEKINxeWA9xfEeoCp5kD4vjUuZB382+Nh1aO9gZ2v4s8tRBxJkdiR3t
Ykg6NZ2wOmWDVdgNX+oogLZLCmwnx8+eklkfQwVWHiazwqEO/6JRKEHgXoE4m6QZ
Js/WtNylN3SmC/dE75d/dnnZv5y5LPQVDjHdIrhdsH/B/pH1nmAYXiccvB5ibSVl
u2QiJ7QD+tAe6xiIeXs4ntV55zrN5mfOvk/p3vAPh6PjFa2mBQ02VyH8SbQBeYEy
V++sD4HmC2Zq3v1onP+3lhixq35GeD1ak+uewvh1mdqe+sPo1fwpdkfhAa0Y0rJd
Cm6y+XrAzFCS8q0vYcG3RWNuh8PiZW/uRQ8SXG/RHA409RcXQEetVh8MH0cOG9nm
NnpohGlrAuQmnNKZ+AsgsK13j+De5NsvgarXJtHbYqv7a1qpF8w1cD+kchi20Wss
ZoZj8bPbJ0NEUH7RvBnomWBEfJ+miKOwrTW7fB8cpmbEmb4B9IK5Us4T6J2A5z/j
TpvzLpwUTUYOQAt/6172fSScKYwGibjNqJMS9mCyVBxOM/DxMKPed+0C2ghyObqo
RzIu+L88ZbKYBywG9Z9gd23MT2oxTTCLJVrqoQQ+8ykjNcCvmVbF/LeHOJgdTBfe
96a7eXbvITvA7xn/DjOGfpMxWMqbSEUmdLOUo68P16Nqc7i+C+d/BsHN3ZswGdxf
AiHTpN22QKJYiL/uShYhXzVAwTSqO/VYK/QiQldTzIJXDrSXyNYUe+A4D7HwEAtu
ZqdNAWvD0zyK2sSjA6zDF1bewsODrDrPa2GpIczgnYlF43FhGsEKO1iaILDVd2Wq
0PA16Z1aI3arFfqpdx644GtzcTRjttQZnom+YXvvbSZgTHN3KXNTT0AgpO8agKwN
oexX5POAK28BzzbHLCBUesZRSew43iGaupyq4GLXirj8Y6kbMKzN0JOAfFeTtwzW
rYu3oXGdvGkSXlNmglYVM9+yAsbwmWabkaF5fftskjoDLZqaC/jFT7d+ufzh1KHV
f5EPqIB5TFx2iVesfKG78HqD3DsWXtvud2pjrsZNQHLhM7pjrPAtPy0ETqF6+ew0
c78ogTtM/Tn/zklwi2KC2YFPhwukdvO/vG0VbiuZHA8EgVjwjgJ6k6+YOurzoYcK
zwQCqdAnI0KBa1J4Xjj3tDaDS8SwbFWAaRgp/rUC533Rq/AZqM7pB/midYvrfinF
/tmcKLusgna8OKDsi5a3R94RLv5Yfqegwv/rsgCjleQUQXpgCbdWCyjwcJYUudD6
j/yxbznBRnUSY8nVI+hthw9CjSzr0LvQmSLVQTAXcpFVsQbFWi2cLD/6AYL3Pv9o
4L7CUyP3FSpVqeR+gL4cZY4t0svjzNOADrQwEw1nAOi6a/RsOYr6bCCydibjGgMI
UaNsZ3X7cf5siAEYLnX/vrwTuc6kE8Tjf+XJlNQdeAevQ7zSHbg3s9e8Q/RlpvVq
8AUy/6mqx63jSAfgSVtoDjnpfLhpAG5Uqym/FAFW52TjeWvaNYzAxI9oHO4imn/n
AdRDusqbJIHdXRQVN7dDAZqYop1NBAl31rihgGIaUuh6thjwo+nI3JK+UHSKgmQr
5/bCRn3D0G+oEBrw3qq8rYnzyuqEygYUF4y1QZUdFBZOIgfCrbNFWQpRRYw3xMY5
aY3yDxC03gNgU5ylr9cfZ8T07KGc0kXKq8RhPgpOxuS+2e/djrmSU7yoTjyHCwXv
1hNd0/S3GKNGgCFpSElnvoaM/jCE4FqvJIgpXxNq/mkLpilgCDCvXlY2+iFa3Tvr
IEw1RmBSvt7qyhZMf9DRc3yrlbk2kxQLQ4RK6vvJZ2m2EwZ1WH3KHy98c8sVgHvX
2fvFBO6R3qf5FClh1b0dZzGInKFebczpO10ePiBbmM/6BQPOLT5cXZT8rsDq7Qg+
q6VyeqSWmnr0Bc2nCWEYM5MkDMRocGml0qUfMAFYNQid49plBhsvsxOfOPHBMXnj
kshyCd495IQv+H8Taqs+txuEnFTqZ4a5Esxy99e+wqsNybxy4DdxfySUUPKrE8Vd
4OTbgOKm2Ma+PpW4CQ8NRE/Y/R1rNB9gnw70gaCbLEQxLMeL2BY2Taw2YyDCDkXz
nWrwpwVEuz+5NgXcKyJYean6Aia+6iCt0xQB7Uhz6IM87w81UFDrzuizu17p4Rrm
pmlS89Umec/ie83sQLJjwCTUAC/Ps0llrdGhoIuy7I1NkhqEiFJ7kpm3uebuffFh
UI1TNR8w3UBv1FMJ23sJ37eIdezTs3C0sYSQdofE7Nx6omkpdMBqKyoI8/885ETC
Ggw9xDewMsMfxTYNCO6tHrKCATHThBCw8gWp75Ku4S0dUJ6UtMQr+dorsmjRsah6
zILt9oEhLqWv4eziFVxbK23hmFSkG7U+LNeLMjyAzqZWnUnmQYWv4sk3n6a+KSNS
ldrTpLumsIyUfoGe5MD4Dry5IPFVXruwMckUarMCkkMm2HLlyMfwRZau2Qf/LCEe
SJJZ7KvKNPJUklXzbqclA6Q90IopiH6JjnQqms84rgR4FozIgF89enFUdt6NOaVf
TcJaUKn+EtVhS8lD+2CLqGSqQ/016cdL+NBKbb/V/E3XqfsQaX3NydsuH+jGde8M
E+pM6lD6ZEv/I65mKPZPAXFaz0o3pROuP0hT5QLRGVF7LzEgZHPQyLNTfrSMtLrn
v2e6swf+8722CRQ1q8WQ08hFfr++yHL35eSX0OLeJqhoF5CDiAG7j0Y7pr71CVOw
ZAYCG7PrKDSNsOUzxZRXVpkPA1K6vi2bfB5sML7Iy5ukiOEGpy8ACAW3AgozBfM9
Slhs+TRSkTRjLKWKLVZEPKNA9nN/y50Cix4xZDqyWBnuhTG0hR0tXRgRFtBt9OmE
FDlYL0pYtyxDASCJEkU1VzV9cTw2UhIUyp4Bz0N0IupnDfDnnxOdQsMmU+CowtTG
d4G7kMRgftsjLV2jyhWVVPGR+zUf8qMdIzBeP2BXpVqoEkNncUS1CL4XAjCUZ0Fk
1M7GJboWPpL/woMrp3uk4paVv/B20F6wxfCFFzkdfzbrzM2w4Mx7FDVNDRih0K+x
Br6gJ0KPNHxGe486TaEFONwYU6gaoKMcVt3/98E2Aex08cXK9nGdOHZ28vTVxzM7
H/8oO6nvTUmZEXwItR0cNxRqCuMkflZpdqnuFmWsk7En4Gv62k29cphWmAvHUw0K
Q+Aw0XiezVmT1ocX8Nw+f7FbfZ6C8G7yZcx+TSEMWEtptytrcr6rEJc2jnBYLBSQ
VXM3aREgYlVrDElL/lvqSLRpZzIJmFKa+HwvMzxxNBTUWRK+StMjo7HlZt7JDhNI
bHIrk1zAZvc59OZGfJB/GPAACtKIAtmghC/cHHzdtTM2EJ7Hfz2GyFvH8qWaUKS0
57Twf4hi/sLotMS1/yYB8k2sgiygOsraFx68FJM0JCkPkkQ5Y4Y2Xau1TtR0yPus
pMo+QxRH2u0EyM0RAR/W0kRzZtSmMmBG+lL3e5MkZkhJA2WY6qpD8aSa39WpjJ8R
FlLAH/bi579N+EGiRQ1eb8GB+PUHBlCdCvJUuVWmnChCptIdJxO80bvtbONHOL8b
uY+HHhmenMmlaq/Urtjq37RmhOwHa3gLqaiSQ+iR1+KFkiacPRYqYZy5s27gXVuX
vpgfrY5Dw5koZ1Mje3vgLuhQ37qUPj8ljxn6cckm+sZkSkrxitnABVj0vv8E9fcy
31jhW37FvmLPRgnavyvMAz4rB4SZo62yZerlPfXAVd2GgWUV+A8QDbESlhIxeaql
gS0Du2IzqQUinkR0xHLLHQ6ePYauUcHNUR0t+ZOt8r75imPh0doC0PrDSUhm3EsY
DuJPPPe0FIhIMUlbx+cEiLwRwEA3zpEaHfgKIMj9rW8=
//pragma protect end_data_block
//pragma protect digest_block
A6HAnt/ZtrnQnG3G0vSOyIKOZWs=
//pragma protect end_digest_block
//pragma protect end_protected
