// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vKfPHzSuPzOQYpAovW/PYnJDsrc72gf3qXJWPU9kmlNrNvqkX+SVpgQtXJtdRjtloCpmh+iTuFuH
6rSOqs6iFGjWoDY5soQ9bfyMUlJfGIk+u1LMpp1u+ZDJUJhC/uBM7qomfMiTBxA2w9GM/XbVSXVV
Nh2oZ9dPKtTzqup/QM9Oyxxxe/VWnd9xvlQs5h8UpK1AVWOomQ1jDE6/fto+lXRBJsg4O6Z7crql
07J2u0gYGwWib5aMiMVhX6sicqanADwV8XEnutaw+8fQ/RSpenxRmovxgNdv0CKWXTpjQeziD02o
XiwnIsfb54Zqo4dAMIkUqlDdyNhGM/D5kNTKdg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 37104)
FsUqGzWbIefopmjfwCjtqq6apB4ozYfIeH1OmW5QreU9M1US5tydbutztFGQ9qZgXxa7KYrZ0pS9
owxT2nt5a5gn0FHfeZgnLu1IE7Vv1c1UpfsFaqVAwa7WWxNX3fTU2DBbyA008cietLGD2MnAW57h
0YXuFsdiYqLU2uc8mLy9slRkMPi58pLsK9A4DuFs7yMB0Ix4HdV8/jPbfWxXG7+IFf2hBwg0iu8l
7TQHxliaNekpIB2WGwkyMT55E9N3QHW/RShBgCxDGHrWR+1DnEoseNizI/6gGNHTW7KGOldwklz6
DxzPFl//9m4I4OJ3/pcQh1QmvvgoGU70sus4pt10kGmHYq5vOoUplH2GBULW7rX1VSHF8ytbKxA7
NCgjV1zpMngSZli5fS3eGag7nRIPg8a/rQcXQcUi+jRQlX0OPzmiGVkCY+YrBO/wDThat9H67zcp
Ghg7PjC/qIg3KhafVD881cPnMnTRNoDkJcfJi5oOl+fB4c3CotdYBFPkpcmFyKQC4Dz5SKO62nSk
BU3ZfD0csXNCW7UPpstX2lJyL1oQFy7ZuV68pHsMOOOVkCRr/ANC+opV01hMjBDK3xisNaVyIrJV
MRWhnNszWJ5H1hOBBE+F83EEYqlyozbPpar7taZjtw2pCWa+tcxsl3DYTKBx3oH7uQo9l975DkRw
BfHwh5zNuRuYgR8UwUXKB1OiqC/UMiha7dUaxE5zkQxtW6v6S8b75QXteDnmBBBeyaNn32P+BnOf
lsavcqpBo5dRnk/NlrPQliXkMOFOgM50IT6fl5LCXrlkHAZ7zG0bzVb1ZYCJekhyLAQaLN1QopyM
KyCkGJ/4nbhLunumN63KVUOPAy/d6RKZtXFC2ByIL1uQD73HXOTXUfTi7eqN3wfWA1EkEMUFEi6u
QZ4hfjDWm98QOKTnBCFQYzwmUZdXJ/VN0D1GCi5fMkBqSg7448w+r0EGkKF2KpL7ZtwgiuL75mOa
XHPhYkGpKXXp53ylY2MihGozet9qYMaMPDk4uVPE85US4wJUUDFLS1i7HIKuYG3z28PnCjFcC7GF
vNrSL+059cvh8IGYrq7zFS4O3rH14GyMkpeJhVuFCadLiQtfJwGtl9n4qZJ1krLr1PGSk8XJG2Fs
QpN2tKIVI2LMM8kDXZq5h58rAyKj2B5spsVPEN54rp4jvXtzrJ2H3jdxdB5gvedHCebF/UYmdel3
vq24rnh++kAjQzzIT/H1R2hdanCl05iBBAzwUVLpFarww27E/N1hSUkVBp58p2UpkRRUkWyJcFGA
1AEuslesBTD43ONuqgFtRANdN6H/xaFUyGO7HTyAywv6uwF/ChKRF0FPUg+UjJEWNG4bGSFZ2hYm
HNjB1VLX6NkaS+Mp8fqL+6KyCZbWD42SWNHKDxPkwLPwZ+nsGEKKEdHPDdGHeh9EXRIDpDueXa3h
q9S6eqed2S0hC35T7pJxnJgj29j0aO9WuKlQY6UVHbYjqpwPdOLJ+KMPjZbJrE+jsGrxiQMZ1Dmc
Ajk4H/OXwbOjgQPAp4DgNpx2eIJR7TFiHZW23/1FLCAc2eSe7CnJkhgv0dvT/py6YhlIB0dD6rrE
f3E08BxikKodCJDlVaN0AKHPcM7wW/rTzYESRtNIpVIovSsdKDLdBf37eIVmcNT62/RWaZPtV94C
cJhOiFMebQvTTUklVkbDgfHEqLJ9rX1H/SSglVNSOGdjOCCKfdeyP3VjjWEHPkxdX/bRulOFMtQx
0CY3YOm29MjNl2WRd39T1b/pEA9r5RvdWuSu+NKGBsBFXwftelbOPtjOU+XVPDzeURgsiNcqDeMd
zlwWeRWxwd/9bldAL6Z/DtGxoUICFeQiTB11B0y3sXN0lOh5RV6bkjXmwy5w8plwRdWwjziqPlMI
dDizBypjbPVQFnFByzTwlWNhPgzrY3iz968PwDKxue+5btvAvZUcY/ndtOF4u7kJ9I9N3EvVFGLA
0szh1+nkwsF5/5NJANN2uCUxpT9jfIuvV6sBiE2MmGT08pW69wGU2lPK0j7IeBsNMofa95fWZJjn
mOhBqH3jPdnXgSFzEY6vwhaii9CkbGFyOQyprCQS9wlNymWtyaSndiECm7gPWUnVdkWeufsnJQOl
Vsq2AtCoPGT9ueqWDoP+pubWqnSdDZqyLaiwH4qu+FvETXakA18nf679GsY3AhhhV2FwrVn1qd65
PbUiIbrw2mbZO2MbkTWnh2a30ikwvuJErx7rAKVl+B/GS/2ILpcPGbCWnoZIN88+C2omteSjPmU6
gnRMBTNXgPNt16Cg4UOpwvrE+r9WeKXAl2e/G44VtfTvbTdN6/Kpg2F8ZK5n2ENKmLXHADof9C/c
m92FBClvujdhFc4F4OReS9sJYuq8Ib4nxcAyjCtlI+ehrBXPdMaHIQTyWKc/c4EO7KjN8Sm2RMLc
wCwBKiwpAign2iEMcX91WgDpt78yAtyL9nwm8SpIFMCm68K8/0Il09XfqSXRaVA231Mc2zSgjgG7
YBSmG3e/D8xsAj/q+c+E3c5B5gC7jUXoTQpmaLTYqbpG4UfUOwFdq0tLs87z1DC+tuWKvygbgdl9
G9iWsHtgqQvR4g50cxw89SZwCb99rSoox+68xg2eGQkml+gwOLDjr8BVsVz1xCLrpkqERpBN/kdy
ggRPEkXrzEz4osfg8MzYXh74XYRLJIPOW2orWwUOdlP3OwaeJJ04toUFOB2cvNgN7TKcGNbuFNMO
ttISrpZnUKN1OjMjgtSX8AqfqkMnnEewSoylHwB/Ykqx88p1WeS5TkbqtAIQRei4j3PFsIJMqv7z
LNBJMiIk/0mqv9YbErngbrSqsg/reX4HS28zdKSn+VhkKMNf/IDIC26G0IJO6jZMEiUcA+upxBV3
InA0Y2d6dff8r7gCZOPOmvSzOzljqZmIo0mOMk7qhH6P0gOesqE/yls9aWttnSTtVFIIRX6lcDNf
e/3uSBHfeeIn58Tcv2RABDwc1qbp+Ph7Zl1rsURUhgONz9kFUf0vFyrh+EDKTwDR2Feh43J1EeqA
rHWnmtjenTZxkKqRUYQ0ZPTgY5pmrO7ss86xYy5xLWJCq8FTQ4E8hQcSFOnWyTXJn1zpPjEOiG4K
wcgC3sMAoGxOsI+lTv3gjsVaGGIOe05qRxLoKYc4/ok51vMf/HvcZ6O8R0I+GxjVH7cqy5wPcoUE
85zKTdZGLepzNiwi7lgT3DTTyrF23X2Xkne9D0ctJbFOaX3qQ2kaUB9NYBAcDtwa5NUVWukmUxVQ
IEQL6yqFutPdyjjP/uHNLZ76VA1EVJAgW00Lam1txkbUg/1SJq+k68B/R+U6MeEqxJSyjfdTpCcT
3Bbt5RuHUDmk8Y/mPGVHoA6kF9Igi6F9DGzQAVyICp+Ulp5/bt3MSRJ+zhKQ8mY22AGRK36WkIVZ
MV8x9BrdpfFrs8tPQK9Z1E5vXmPgpjZUAmz2vNzu6AhbcdaqI4YS5pXWcv0sfLzCgvOh7J4JbPab
1KaQK1saxb49e8qe1n2dWjYkG0SHuW6NTND5MXqOHmHy8DdEVZrM1vPj7Rv/is9Mq55xP9BaONga
wSP5iCJHAChJPl2rFSjM2CkDhWk6zs6Syi9pB6JRvSxvGzCguqOQRu7qETh75kw4W6NNc06g/ufb
r4Yw9zukLGxI7QcpWxLvEIiT1Wnha6zjzMcG3QUj+T6pAKebtfsP43kLhi58FzI3lLSIzkaIqZik
IHHAv6YYVx96Il+tzKTtAimU/wIDJyi8KhAdj7LWPPBFaQ+ciGes8QB78dJxvJcYMFKv1TZ0HPsD
6yTZlv/yK8XB1gB1e/T7AGGKoBG20zLNbiz5t3th9TJC4bZ81ypdFwoKmUFFkdN2K9EE9MbXeRQ7
wGVawwbDGutHWJhMS7W1rEOfcnhFYiSQD+SLgkVR+kXjgqXDEhfqsXgjw/joViWG8LVEeP7AvFD5
csyFt/VsMgCV1tjqTa9rVP33l3GayehjkalORjqpEF9iEgjeoVwRQ5zYbUIm3vLr9IdqiFGAhqSQ
oDftb3uH5RUqdE7NeiPd48+OHc463yUdhWuHiPnHmPN5bpHMaebqxw3Vj6q78xlQY8Y5BCL4/E+n
BGQyczu1CMat9QBaFhuXYGyoD446DMPYQ/m+7bAEhzNqpctOR5ImK4tnJ3bz+ukxPQtkX3qAgTGX
TU8vxa6ut286IfCNcK8bka1aq68WbFvo3Lsb3/OMQlR77UU9Q3UWI2L1aImBuodalp+REhb5FyBg
RylQcJ0w4/mIE+bj4sVBAugO6ST+tFvHaA/d42fV5Obp0NZZ2qsUNKyBYRjjM0jf7xJSFT8KOs2C
PGrhCGkPYRbX8eT+y4e1PKyOCskbeGyugSeyjeO8bNOYsC40N33Puqne4ABiokVRQW1BUprzJRII
eC4pRu6JwIBAwwIY2EWphTgDxsIE0VpcmFBqq42ooN8wmZl8TIIVTuF8AQQXAojwKFyuFD7WXI0L
95wAYnI6OLIDN1bF6phPsmYeO+UEjENqiN7fYaCvdRN3pDh1f/LuJT3saXusG07kJO4FhJEIPAqL
qWGDB2IiRowk2NYYcFHU9EIs66aNFuuAEQhfW4gCQY6ZU13wJzd9keyNg3hFe1lGD/2CdxW0Y8Jz
VCOc98k6MzhxglTgctzYM8HzPlleEJkA9dbcB3jaAy10IKSpMKNa/QXZcxPjnoK/65kC7Em4vT9k
g+QekX6c++ui+5ohkh7+dPqJcM/eONxxyoWpcyg2ngx4btcYvYu1CG5DMGqKjuiRo+Bd+j92UL9H
sAtZVBcPgqvO7UHdg+S2qbgVc06s7XJ818L9eQiLTHid0tDePyHVzyJjrgrO9Wwn1fAtQdecV8xf
mqe6LvbI1PBuGf8+/L9TLm5yo8n2X4CAxA/leI9UGFxG+9AcirY3bC94HGNrYsX5ZBe2DRYUMri9
uEKlzApKuXEudfSw3lzCt0P1NY+9kp2ZvcGJc4QUllgo6yY62yhe5iUEWdGySVSpQRkuhnc1gVwr
2s4GSgCVh3zPF0hOG2dseD6pm4oKI1GPmlKwxNAsbBCnooJbU+3mXtMyfiF6b2jwUBlYdpbkwNjG
+r8EqGxW6NacKeR8nb8vZSqM84M/+KFXk4Av2FAFgT6lSQXE8cdH++AwrLuQAiOKYfXlWFDMEZ/A
ww9vdbRRF3r324RdN+15YveKGhCu9HKk16hAVOSXDVu8VO02RAqopfDMw4PQzZJ2s9DD8HDurahD
QBjt7yUAhSd+XFQmI6VqmlQpbjvZ6KIXNTs8y5q1L2C8x1EuU0Tg91621gnAUcki9H/nNa7Obso8
uYRQS/IsgkBhaVAsU45zvEupM9EH+TAUTpV/TndndIKUjLyCMl9bx5z7/e0kkXbZXAO47Pw8L5Q5
ZcHbrRkSAcqOwTXkrpiWFaV/16YiNZvDllJm7uMPPwc8vtJd4YFMIYWCSOpbi3EG+D284XElvxY+
AbIWo+S241qoF0xFWc34lJXMkjv/WkGpFVJBdP303DY2RmIHUg00Yyr7aDYlWMKtftWp+FWMSX1z
Jdpiyrq0/s9E6pIoK+KZEYrE1VGjIaxP9JP3s3rrde+V2J8p+Wsf0LSZmUXITyBLFyB/aCML8N06
7xuledmJVP9QlK8UyPlx8c/CkLZOlgx7hGsnnd7umPDDoVA0MnS++eoKOzZWuVa2/krUOUnMfqbG
IQDaoTHP3yG77tEn1Xzcu2eQatFSD9aDPrjh0eoTi/1a+NCFi0Nr3c8FRFeMU1wxrggxO5hjJ5gA
wPYrclWYqmfSIgYMM+pIGkNK/nB8eR27IDdSG1bAaJPxcUzBc93o3/GecFk84ZNj2dhKnB47mrQm
Xls5G63FQNi28ytjkXGtWki4YUfITxvAJG/7TeKGL+d/AXb8gkwXSPEMRmiJQZff9Zz/94N/xqoS
tMJlS1hRa1geF79hbyXMFtA9k1AYrIjQ9Mfy9Z6UNOAIsR5ArmGlEqXxUacDl3OeVLbrEJvwbVLL
dU0RiE3a+Pe2sqM2G4df0nAo3xpXxIsuT5p2hzw5FC83inWQmDpOTkaALySVyAi4KWTT4YobQhqq
ktvly2ZOAHcLIIa8K177D+OjvEuIyTJiWAvNRX/mNUkUHxboSAaXI1NxO5VhAvhYMMcj5gHdcHyN
ZIrVgKCeAc7ieUW4eC53ZZDxhExT0P+AVeQLMX0szU1su6LW1q2BEXt7Zg274ULKzhQI/mjdYVzn
ZUSPClQiubMY690QZR/EITZ9QlHhvEAPzPwcq00ipKTE/k3tYffkRWP+ECqRRYOGM9k24N2d1TBo
uTmx3JA4lYsxIXX96AJB/0NMGSTbmKsgbr29KuKFSPDErrLfyNs906UAcHssNOcPEvcksJmLVT6M
6kap6+OaLmsv9p1Rx1/tnEDJixboW5xU9es4rd5thULDInBJtRwQ7891vzn+RI/APOxjh1g+yfHn
4mAQl7SA6DhQti0+TegBpzUKzXVX6gwqBzaHOyfeLHA8NBp7LNdtNCkbZz8LGEeIWCqYDznA8ecZ
zJqiB5LamU/8ejuoGOivZretB8BFfRNTSaxaQfniKqqVs0Z1aO/UP5aNeHiy+kXEGdb68NnDE/84
Ns9Yw1X5uNbIBb8nlsOXCbSFkbtzSXwwLzQtShMRqk76v93jC/p2vJATRJv/wCiQqX93ROkpGOFf
eFwWEMHqu3E2pGxdoMMsSA0nIiVXnVW85Z9miChB0sdYKocdxpT6DTf8y5XIUQmMPvjO8fR+z/BU
wQm518dut4dwD5Ql6GSN0yjH3CoTB1XoMatOvCQNUQlshTzL6SvgC5QwEKwfxzR2yB2HMcsbU6Ew
QE07onxwCyJW+96M2kZTjwKYVSREXMDsFvNs0x5cvb3SO/ClFeCiObyv+zQNhUw64yGPUMbwZmeA
oJ7oHb7lWg6UKNlXQfaKAP6pYEMERnc5R6qagTHtGidWUS8lT3zQaffkZqeEU/j2mCHEDwzS+8+W
uuT6wHEMiw5uPDUXf06s4Nh2PmWfLeeT08QvjeqptozMnvSJToLxIG3NirpxYpaXJpCf4qSSGvcE
3M6774MOEdx4eB5a7i+AgtODvTWzq7ML5ARvdGZKj6eMw5njTA/kSJ3Hskh3IzYD8T2sciunE+BD
Tj4fWamidovg4jcAUv172GiQa3O9y1XMLgIX5CcqFqDNvjU/yoVpZou7dwYoajsjhmK6521cQDBr
Tu/JqbJq3pIbr50qRwXnkfzsg1IUPyIQOTjC7D3nKMYczGsITDadAUx5ZuBc/qzbkuTeItR9ZGko
dCbniBDOOeKCejgIFPNo9Fm8jZDlvUO5+4wboGXxXWwV68id1BL7u642cHVtKbxFRzQ/5d8kaeev
n+kGHrLazauahvadbzctvMm3KgeQ/PTXS/JEoMLZKOl5a1AORihnlDyjpdVVEE9vLXCb39nt5Q+0
UpRfVGyX8KQvik9yPDIVk+2L2N7oRW+uagc2AUI399sA0kSSJR89/rK7bnnRtBTQR/9I4V+m+FJl
OEB4hHE6/iQtfKtK+AGclVdkty1ZWZymDHREaBHDFBEIBRfnR2deMfj9QC5RU4kvy/wro9YkXDQH
sTIAYdtc1sRrLiT7Z53xRgYhqGWtUsCdC8OYUnDlB59M988x0/8fzRCdzAq/lXXCxXnpw2dUIZi6
2WpQDcmJ4RtuEGmxSaCeaE4R1fT2AsvFXcLQY1yi/AF4EcN0+5bXnUw8zGlW3Dpc/H0gbSgOs8sR
5L3RFUbzItjSyMq5AQvX/0puPuElMPet7ovqfQoHkRTiOIVx9b9Ul8MOS2HuaqAJqojp3MjZR5wS
uHG7s0/gkRIY57MZiVWRIWP8tVr4hShtePbMKklKbL4Waz4HCgvSJk5rWnk/122WZj9p5Vdjn5iW
VJbIIXta1ZgSm7r0Zl/u7PGYAEIU63K8m3YvUelPJKc2ZaRYbydU5D+V51Dm5Shd9qPMbjRR95qW
A2j10kE0Z9vwFy2BDZJSO1N87al5ifIm5J5HXTdA2ZeNOfL9i/onvGQ5PU3rbFZ/ymOS7yBVJMAb
t2UiAp1xeRY3j4X240OoCl2AiIckIdnnaxL7QQMgK6ObGP1SoPDEkn7/W0ky/AG2qawLR5Kq1T8Q
zOW1XSB32lXSyLPD4D25mFV+uiqAoL6J8X8mZMcmELF1+afJQWeEG+uaV0kjUHbBmeq1SVT9zAzW
k5lkYqhV1CTB3Hbfw7ZrcVhLNlHRbkqn+GkY4yI8ir1mGvPKKr5k9nQUa1dh7aRCtQCVFzQKrcnf
5oGhMXysosFpdnme2LeX6ddTV9v3e893XTgSmsEhKeu6Ttu913jXCFtVI8Yt1/nCZZdoKX26TJT/
O1CsY9UZJlyzuAbT7ifnktExWzHtLLCosvhspk21Av9w5ir0sfrdI6VYdwWrKoZdG0QKTzM4PnSm
6DvtEz3nckl4Uw9mtQ2cHMhJnMaNDnTIUiKdsCBqSfAdSt1s+sDBNvg1Yun/QmxBmQk5cdJX57ka
vvhF+4cT/yepFFZiLXRrFN4HxnL/MqANVZokDyfG3q+fXGcbqqrwrE8NXsOSfj8yBFfecKB8I9dy
CGhTp2V2rWeCdvA95LJ5zQ0c3H3Pc0qTZ9GZtdWWBRZeH+FCRcirnZNBGZfHCBVdALTCZboKtM8u
9L1P/iNgU0S7w3rPNfyBwRdj4dA2P8Uwl/uzrkZKd9o55CbFVNx5RN7n5gNBdVVcGZ/RKddeS+pT
ie4USj7c5UytadHkM8mVVqBKjsLnIM/4LskU7DU25BNvix0tYcfCZJSi6cNXO1MEFTKlJ28gmXo3
ukyWizClq54bNB/NfCuhw4FwDalLVP6vvHNuBvrmmNtqaoZvWE8gdMmmmRyihRyktYgCH8IvMvFy
lQcK3LTzx3klLQvhRXiV/T28vQSrTf6a9sQgsuYwOatuJ5DxF358VexnT4wPcB4w1+sxXReU9k2a
X9m5SGg0NZYVKmM+TgWmpvgKMlRLyk1kz+wfu8eBxZx+I4/xRR5YU5OLio+kC1W7/4OjulW87PVM
bVqL7yYUTVeLqr00Yk+tLOOHAkPqsZlmdtKGorAop5gts8O+HlwH+WGW5181DGf7BUG4N0RRPpWh
9oSWAaaqcambM+45YSzrnam5VPvDGV/SZ/cnvwPrwA0XxU8hAVZeWqPU1cdz79wTACU19AefuD8U
1NhbOGPdqU/s5kXkp0XVleUOy4/lR2mCl5OFhonQOiwDpX6RcHF1AGnt7faCr2qRZ+BiolXgAGgb
ECPjRwZIRSyAvQs3J9BhmJZYiZvewsbEl0eabQdNbaUHPOAxVWRf0rlVkrJUm4TkHTHxgSsSCJSN
6TA3zivYM85CgDqItgGgPzgKpu3+steHwHxu6V6ySbowjD5bAduB9x28fMpjtpaUKo9Nv7ksf0lS
mR+9/OZAKDCQ6/HvjT6ML03SzeNZ2N3y6/KkoyvCbheZ4CSIwRNzAtiqoPvmzNX5GRd7XNMe6qan
/H0AXCrudeGC2t06deVC1zrkQJ9Nc6HEqqLU9+7iajab4J4BdasBB+okfmRWp8KZB8MMRohWHB4+
EN2AOxQjb7AvMgo4DcKi2TiT6aSFtyahp9Jdl9ZBfZ1fSYIArqJN+VpiqUj8CPZ2X+3aONxcgRyP
lxd5/BGZn8V2Vj3T6632qIjFJqjuuJLa0Yszn5SzzKWAiJ5qEDPBUOGhYhrzQCPPHcsP5fYa8BUz
v7vvh5f4RsJqzA2Cb7cQ7Py4jxYtirboGc/+bDT6taN62MxFRUb4PIN4gfQFLy1YN56C1IGi8Qdd
6FzbByyPood5IcGKec/zenatm2/3qKTZaHpyFYXq2StNltMIq5koDsUFHGKSUg7kBgyfTLRKEhhs
qcfFyYrJOa1B+3lqAz0Sq+jPspJ4wTkm92GY9pjY7ZselqNuswj+9SyGvzOayV0j6Jk2fFwwdHt0
pIGY5m6WXvVbQLlDKkZF5XqU/sheaLulu0LyzmA8YlIP+cjHNSVZnzmKuAr7SfcSXv00CXru8wLU
PXwgavQbnrRwY/8t/YpYh5GSDZ8QL4i0/SIjVt0YsRR/j119PGu5VEw71wZG1jUIYObRerROWw3r
SmCRZQTcn5nHQBlz1Cb52WbkARllhh5JXyyjWsWrb/kVrbx9beFWwoXJd/kpcAK7Owd5/wxHJA8O
Qeax56XzFiYlkPqtxqxU3JCN7ZxQ+qfGMG1x5L0Hmeva1H12XCATcLXqAN8Ymy+2qK77urA8/Y7X
tNkECQmdmYMVtqP44M4g7gice78r52NL6bX2iP0Zdu6FbVfSHG/+3de1lsNHg9ME3C/wu8TMrOwy
f0NSC6nsEh6fRVnD5UG9ca8BjETVSr6xA1pvTA0CG4Hw+MOfbpwPHeP8sU/pwir4saJPAFQWKY0Q
7wpZgdedTGdL4PUfJs5fteKzxl2H/v9k5guJJUrULnZ+YjwRJADU5dqOGESJTND0ttzuxhk3qUOn
9L0qsISKvwe/uFM9IJJlXzdKeLN29eLjuFl6CYPCmV5C81ZFB+a3A6Ry0NSpBLNalEFBJgs5dGR+
o/0jnIBYPOEBqEXV1MO8sUv0kRcM+yK2R3SwaG3aOfhst0LyKO/P+xY/cWfK5lqf2goevCbBvXCN
MbETHByAORQzr+toD1wUcr9lS19GE2N6sjowhr42G8egsbNPuGfzEagcb0ekaoZZ4qzII1UpUw/8
cKb11pipjSOz4eVWl7K1BDVU0428LUiZMARuqRBBBWsBTNclWM5bbYcMQtQzMXVP4hVR68C3XnoS
uSeChazhvcDIblPDF9Fn0151rFmlpLKeujC6heKsxq3kS0eHU657VZLwkHuKHpd8cLV3M2zjxGE9
twhYPD2eiKvRsKJMcv7s8LvJpoDAScXitTbj44kGS8dCu2EU6ciNPEGFw+sBA+2XcK14ntCHzMbE
XbJ8NqkVxI7XOCP9oWuZxm0XLaanHeTHM0dGBMFX/O7JtTjGf8B60jSMutI5dw0X/9jRmay8+Bw1
4p/5HJ728s2fT49ud4vOjndyTjlNsJtgRoUKb9Q15VQqn8RlP77JmiSwDOLBceAWLkp5PWJxM3tl
dojYzB98Zpq+cByc6JXmXN4EKnb4yoKqshn0jhDGtaWPjtdxxkBiMPEEqDJPVhBTwcLppvMsy6TH
5lXrChijk7cLAozImPMRo7wyqYP9Jlg/gElHLh2S67bnvFZKOakPPWeMnh/QTSCJUps3oWUy3oAp
mrPzFXUFAIhdd53p0OcwouF6mvZ1wy4j5p2RXM9JN/hlo51oL3wUsGPcS6SCAPtWVlHORxnqndWg
RMB3sqi73t7sRBUES89Gyf8b9+HLTbxme7X9yrsnJN5HrWJJyNFo2nTrnwzqApWOuwnEesftgsKv
LWvD8+znp1Iys+HAuarSvD1IXwzERmd+jobH/pAwb0iOp6iI9MCX7rmg6S6261Ecu+nyzsl6dwjg
E2tXqVIDb6HJ2ey5QCfgDY8/UVJoYAbp8TdhYgMUgYef6+4SIG1im4WixBtbkaiCAUNBD3PDSndr
VZSvPht7YYYML37zlKrOKLWESY3AgmS/XIEFAj8Le4pCUIoh5VKHscndrg0Bj336SqNTRxFAYLKv
q2VPu1jvjTvJU/FU+K8lKk4ooBi3HHMm79tEozxxY3QcxjAT87lqOxyyUOHS3rkzN8kIIkNdfUXU
xzcQIcJ99+oeuO5CX86PXa+mvHK2w0T0ycQPZxdA2dpE4G/UCjuXUFCFQyaYhPQubx+TFLUffYqF
yrWfHbX2mMABrWv9xOQ2Fp/OhRvNRag2jOGEIaBw42uZU7sM8C0e2M9GbRVC7TPlJ/mP6Jrb2hvm
lEirW9mbZyaavgwtl18tKjxeQKdN5CA+x2K7YX4uUfdt8z6+EgiWSRJ+SDAswUrTaBMlHN1de5Gw
ydMYimPgUqI0lWUeHXqKpxnfhw3yyxm1iEo9M5jJswcEMjTzlv9idjuR9/qt8dgucc7sDIzE826y
SL492UJSw4+XnubS6+RsS30ySTJ7gCLm0dXUZhKv/MQDsfZBmYUlKnZGV9O0QGRKt1y/8iXGC/Rw
4m4bgGCpPig98dZAUr5h7ikYZiIXY595h+HG+Au7CiGF8NhtYfkesmsGyUg1w/JKE6r7zBiUaaKe
6EXRlam1KR/+27lhsW21d2jtcpJM+fu2gdkuJO33I0VOLA8kWPjHWVcbAy24waQWjeWKNzPaqsZp
esuVsXSyTw9KRoqa7IevmHWx/M1+Jd8Ob9+XbLKfQGfH/DJRfC4LLwwHB4UqkmCIefcocihqHiih
o7UG91s2qILIAYqLpN+kmHJ2ASOH4B1FDWwabMk5xiVjqJNqEJ4XcWWhCo5LpS36vOVNMd57Bc+R
MaC2dRdnG3Zr3Nsckf5vsK8L11cWvSTOw4zf9a8LVPjyGM+P6scPhFxeAeE1J+MaRWXxS21qLz9M
+eRgQPyF0yuHMRT7Qp0YIzkr2i9UMLUzmflPTBFCxCKvOKw/VFvlp3nCbiVsb7YWnyMYERk4WR04
qDXhcEEro7iSwz8olktmOi5gzonDzGQ3u7KLuAqJ821L2qYL/XEHtmFeKzdfTdnd0Kby3HT4trnl
Boicubawo3aZSIPCNw/7PEjdNC2jSTacmEh76vS26Ae4T071WsaWMqWERTRUhfM7oY6YLy6N3dj6
LvwWYZ/wpz5jfDiDVGSBuWZwbr+BnZwFj9GT2uVj1dzJfZHZmAG5fVKVphV7fquRSsr6w7xq+B14
SxPjEOllVn8ddsFtLxcHDNlVbPC+/2o+yXMl0PLL4V72OpAZ/VXEo9XqSm6C5PTxKpEz2SzGXPlr
fM1qmXoClNOFlwF8Q3oZFvc34LtP/tULrfyg+C7sUFI3/g94GiXZVM228G6fWoaMkWiUa93y2AJ5
rETHvsHuhUJu10dOqk1P1LR0Upqkb/YEhEQc3jv7S4vlznNk1FKA473un7HASH/GAe21puTWI5nr
/BvPGhR6qDDnCSlC+szRxChGIy2OfloQ9FlIWMoOVRuMGfj6tvD1trj4R0D2yeaFq4TtcF7oQNjO
ooETtUrwJGcXuxBIu9YFkXUYFS5l81gs+hvKKYbAjEFel8esZXo/gBgJwjMc4+71pbuufdSJFVsT
qh/tHFNksUxLwyDterDL5V82j7yt4bvA5CvGifw1cSAUxJlrkjSw4IHk9cF/mzLJq134fQi1I6FQ
5aFD4fMXkvVrbnZK0gMOTqLKfsOy+/o+pZAw23BNJfQOkBGGLFQhy+XfscQLyqDYRmT6wZT+5u71
SbYJgfkLN/DuOLbQO4NGbP8AEmZd4D+mCppljjzfJhqiX4XFuQCTeeZR3I4v1TjxZxZ+HE6BC2/k
vbddRb1OsSDlmGK5WOq9yYUfGAsell9FGS8Mp3MnhctCD6yPtqej2wYZ41UNvGkNV4l7i+75GCaG
rtvlnBaUp+uHO92FzZqzoMsSclaCq3R7n82/yMsZ4V/IsehYRHFYPww6qbxQ7fI9gdgwezIVpxcv
n358Kwh0yuh2MlFAYUO/+q9pkHwe25kdQAuoFDqPhoKbATPaA32fW2BWPHT1518crlYtMV7C1YQa
xUE6/ZbtYfAP3+T5APLQGgffDAOdGxj+LMN30iQdX6bs8e37OBg6jb4dpK/ETIqKBRsqIhntiWIh
rCKaDHRjTABfc+DqJL7WKswuxGk9V3GylI6oqeWrYZQUfw/Wm/AIn5ZCbKsPPTrSWvtT2HhqPKYh
i3daE56fjX/BxFWT308AmXPdqlVuRDIIOFqtKw9olcT0CSquYJseRPuBaevYg83SYFiK1YGzve6K
DLQoUVHf0taRTS5XAuInMWel5zaVWCO+dHi/4i9lbedabwzzdbMFdYtho3N3s+jSyak3qCV/tQ8q
EnXGraxMZhKSgTthaveBGbegPTNPDb2ewRINPWg3DymQaJ37XM1Rlv2Rw4MBp+5eCVlYwi2EnldU
AsFlVCttsLh3aLcGWey5Wd1wolH931pDnfkajfJewNPuzmQeT0lYKBPGfwkIFNLJR35SWrMR0I1M
T4nzoXaKpmREfSuzN9gW6nfF9314IoBtLtPhr6kyeiiEkrYkwCMAa01U10YHyI29E0aOSJUzh36w
PLpU+FzOmUUvkrHqxmx03vbA0yDZxGxAwMGMls2RGAA2gCOJ1X687DlfDF2v1/QI8AxDwamZ22ok
VN0hdvRNAGeLYscu10S/Npp5D45I2/xfdy4B7qq8p4GVbYp7HeXsY/ZQ2IctMVFCbJkQRJDlFig2
F1oPBazwbw4RNVxlmjlJ0AxPdw81GJr3rhVNKp6YRaSvqHYK5qBiuV7f0G9anGSdcc8J7wk1HAy3
LnZGdiqEnUqJW0XdYe9zlM1B7waR7P94jFaf4WbQQ1Pdh+NtKlLRGEx97cVvcdTAA0DVFT8kJUK+
LfQe00l/AzFtRwZu+j9toH+aTxpoCaqMKU/qfc7BUadZkuPzBvv06tXSCdEuUV8FXab5x8FXzQJd
nTfA6MApJCXnqCZPoaQAI0nwtITOcjO44v5zvRyQ95HY9kvzaxZ+4pC4D6i5NVwpLU12hXlahONT
jYN8qhPE+1hl3sFGLnJqZBmBWHLcs92dhoGXqfOQCA4u7LIJp+VGzNp8Ztg9qVsEoCZYgXRsFHIA
wjsIAk0nYyXvPWZl0CfMvqnGWNyRyU9KRT15691RH3YnndROtVpdZovtJxMkyP9g9E3V25Bpotm5
e2jnOEMHUAbL5k8uyeTOh7XbDcVwlde81mJvuho/jFhlR0NgFHnR9RJ5jQlNFu64gB4R60nuzi/w
SDuZj2tNqNwnE9awRkdoK5amscG0voBsHiRLKPO9ssc1gqeKfRvZ2mLv15Z+7ECbo4uPL8z0P8Mm
hD8foKqVB51o2Epq8s0lqQstTbpf3C3y2FjqAsHDtmuHfmFngVEv2Gzm5wwhvbqS1AZRDZtP0Xy5
vB93q+CCUrU4yJ0pP6hu3tPljFKBINE/bZoWGezLVeQQd/GARwM+x3JTsGDWBr6wkmmXhcuFA/Ll
tRmw+17aZTrPPwKQ63G/H6PQqplITEUhbfirCnk1A0ymZX4ZQwJLhRo8SGdX0vBog4ZSPIA76aWB
qERlxKX6Yudy3GjbtaHhJn4TPFD4N0mFHTqjmleLy0AnhPM6lIi5MaDiT7FGrhHTyxHwj/uIX6hG
yrqLG1eER1k9kuV3sVwQUZERhzwMZ7hAqTyednJCWeisrIG6vr572oWxfbHrgJG7kavz9dwn7bVc
ZW3LuxINPh0KzdikAKb6F4aW0NxyqcchdxwJBtrgLyK4WAMZf3zQaoLSzBwponnpzLmm4fwL/I6N
S+F4vLm3jW4XiyV9+DbjUibd6ffF1a0HJP0nvPcMZK1KU8OhaoN8lD9MpvIO6z0d4EYtDyat4K7Q
Bc65b277cVyZDvOhX2iATMlFt0WE2mmrYx7kfFvSpFWHlq9ka1jlddBoSAzjfeMHMd+MkpwGE69R
0PvOUtPja1SMrOTD9Nbx6p3wblcm0wPwzjStXrZEPVIoz7IYwDmudp5dF1T/l7pgQPQJAyWAYfjK
rCDn5BODpeAwPdOyQpHwnvjMJnsMmD60zI8/VsvyN/ZpHvsXNWy5kJUBonEmJz6/xVfxiPIuqWxI
2fju+1EVGnBx10vMdiVxKsoWOpqZWEeZkBAa/GZOfix40GjRSJao7aMSKftdk1mqKGvb+fRpZwmD
Q4MUMxWJZ24pz4jiEaDkU6Qov01ACt9pVCyg5pQou7bmxdzj9nOUk1JXlUkbZJIp13tf5DeekTKw
nJ915buDMPw1U9YIeSIZJYU8mwNpTJzAJ+3HBwUi+CpQzp3DkeJpRkZY7dvSMNScJRmUwegZyDs/
d+0WcLKp6soSKaK6j+rNxdhDLOYfwONHZ/ZUbN4Vi9cubufZPeqei3DqlGqDtPtDuS+PCpbfoG+k
k3TJuzcMZkqQa6X3rxW6/GYEStj7glr8F5DSDJmTaHG6Df2FxD1QDrXAPGM5Po7ThqrYNhbOUec3
8jFagOJPi/ddxv/DbShvO6eLKK7Gi6vg6fTP8xyDwuSPCcKRpdaoNnLKTgG/0LX2b+q7TdoGKKE3
GwtYkdvKdqy+6sF8ZUEu6ovEFN7clT4GcSVQyIXca7IOLujTQm98lEGQsPSribF6V4Q43v1j3tFZ
+w1jG9IN+Y3Q1nVdJj8MA/7fQ+6k7Om+ZnlCyAUDGYAY9wNAQ0BG5AYIsUVzNjkESfByS+/ZcOHt
77o3Oiol0AlW7M6pCJFys+SgkwuQ2aIiuHH3Teej9UnHFkBE1dQGzZyZmq02cd46p/YGtiZ7Dw2t
JpB9b1mXiBfOj6jhsHXFyXfYtL8geU6H+sqtyDKbPb3fgPDC1FSro6c6JaMq+6xWequZialTN8Pl
HU/1kcYST6XlEeRJXnOLegwoimoKSXUvR8V7zVu3pHEYeFB6OWwrU/ZkuZkfA2H0R3jFBSKHuK6c
fw5v1g3vg6EtBnxJJtZFdsQX7Ykg9MCNAUP5VCGRpbDQDMg3RNaYOh0/ciAWI78PTfRiATuW4K4c
kifEVfbCQ83Vx+DADC6jiORsS5IpuhAUAgTXaj4dHApmv8HRfkbt0ZaKkguvtAngL/H9bowyX0M9
QTp8LUW3vVInS2IhrJN+GUSj3FecxcfZiXoxQQ6mveSDKtgY5f3qWXbsUbDqypmlH3iZuH5GaZs9
L1cbh4lPd+OpYNnOY7LBCj1pDnjqlV+MdQfY810ti/TIcdyj9E7grir4iRjyKk+Bq81Um9gkFv2+
RlXuWnpkMdNiyGVl8entppAhW6idIcZfAAToalw05nP0l0eIicbB2JJgR4um/NwGuV5bZPiFgpBK
nMIB+FJhudhfr5VGMMqoayI4G4upXvjfN/9nK+Enr2waDRJgNicvGsyj8EbOLM1ZQmOkaKDlK+kU
nEb4IlzqbU4tdXb4PWzJIxHs0C4hfmG1UnGMTQLuZbySLiE5h3fo2ud3/DyEw0vXUaVISDM43WsH
BwEYMQ/i5i8hfWudhrald6D4H7nAtVrH+G6l7pjFega6OvqnJcrsMpGtIXcZl4kkzwlylICLDB5D
Dy0Jme5uAjBmnHoe71x7+Mjk+YWFitCb0scSuNr7J0YdVufmw5gpzFMCB61nuCoegCopQlRAFXpo
2EaY1wywZQ8n8k/7vl6XxpfhkeQRirxCqaATOThnOmGszEUwZgCdfWdCCi2UVoLIpnX42sQxlSr7
Rz1cwHQIVKKHfPcTR0yyFZ5CX+j4aMuhPH3SWb3/7vONho+dQ0p65GHtnrpZum4LhT8nVbYQ/rCy
O/M/cAaOx53pGTFSRugdrAIv4wQSmxjg5oQhqlLClWFVSLWXrrKzpqVI9YmjgIX4VH5e1yjpgv7Z
qVzgQSpkmpGvExk2ll+m9V8Yh4LkOAsi9pcq4ROajvzFytcZtxW95fIMEO9NrW5+Mt5pWnQur0dl
2rkk9pKMFdQxN6vLxqccoe1luAhO5xZO3xslsQfgnY0LCkjIzafeO+d4V8aRYND5Ez53EeCprTBQ
72Iq6w2RJlQDd517qADUSqWjSyta/tEn/8Qv7eHzwfdUZE4SFfSL2OEAzFpnWlLmwiIC2CDGFHSZ
fcqvgioadSSiUtvOenJ5AvqPn861oF6GEayiY8TlE2djx3u1yccdiQk97ZVIpXubcHjxy/V92dnc
ceqgq+ov/7tMX6ABYtZXVtvPgMrIjwsnTEO6op8+tDDkFY+BcF07FTm4dd55A64/e5/j2xiZP8lj
SjUludKuLPC6zIXYXReAPXZRf+OMXK2iKsjMJS7hHJ4u+B9bXYwGmVveA1su+/JqRrZ6N7If3ye2
iIbj2e68A9tMfRSvWPnSHGObddXTMBOX1/bPKW4srfcEbNMlZj78DSWg1mO6RDnPqmQaD+DeK70p
AQFsKZxY+qj/zeC9UXjc/akE2QTmnsbhHpPiDely7BXBUjW1IFn6QCvkgmD7CZZzkf+ISCCN84Wj
Bc8AR/dyzPbpcNem70M98wVrOSIcG9/jNubcFertNXys+D645jIy3kw6WKGyUwvsXg32/pATwxIC
nv6ylj1GhIdzSMMtvNPvxjCXEKGbXkm40bcnpJwXUnimL0l4jwQEkUPe0ovmwQaen0NFvV0MuYpq
orTlX597C/GNiAa9L8kvTds+91PjWGK3fcL12wZCvtdlVgynEzzXHHKrH9mRKvtva2m0/qHbACdP
+lVUiiS7TaxP/Dlx4wbX0u2LzNXzcZVAyeAHuMmxLMJNJ8UIQP/26DHY80tJbMRm5d3fukImr7J7
cWbrETUnzR/rzvtZa41GF3gUEWZ5T6OSSZyY6aYU7lQGq+rsfrxvbQngjHcf3xeH9R/xdTmjQQD6
HRUvr+R0dHQ+v1JudJJaIcekAErSNXlWhYTfC1V0/aQC10c+YQX0q+v8LjFcUNhYIWut4NDiw1YJ
4f4yFzIfMcFrBcuLdnLJc6C5Sei+zx2IiIhJkAblMHcqwNWW86tM9oFI/YqkpvTYmSXXYyilz29l
37ZGZV8lErsEzmeGcytnILEnRMt7u/0ihSzFbS5CUpYPKo8jgrHR+wrwbVD9ObwSvldi4HRTH94z
dZBduwwHiYcVpKAEmA0O+Pagke5jA2qP6RKZgAw65cvx28/mgkc+ifloE64J8bihSKpn1s7yZfQa
bm62/74oHlxRaNCF0qdNm3UPWx5DrjSEpg7diMiKOLKgPXdI7FceREr5fZ4GSIlxKFmyDKOrGRg2
v8ydHc4qGL6+3Imil1oQSRBNZgTTZmNj7XyytXHo1UYChhwwjJfjCL81qGzKSPBIvC+J4sHO11FK
p+eckuOx1RgIEWQ8Sd8+dCj4j98DY/NK/qZCrUGo5iyP/WxxyWNGEYGlAVLUjCS01PnHw8UU9joZ
m9W1UeKBuQCzFYVJ6Jpgkq0fmlu9ITGImJE6O0bV39wCL4bzj2SUfcabuW8HGKextkFBRXrghWnw
lyp/tu75sn6VxaHnMHFLqLe0QR+F1ZEJLzraFGgw62pndyLExtenqYwf8G0g5e09jC2yqetbWEov
FzI2nstrYuWEWGnmGpLQOnPWIRj1PUAXbsopJLuOMs52lmwKvPi/2FES44Rwqob2KrOts8QPv4o3
2FZdfC/e80IaL0pbSvtvV2oEX/tSWQhG+4yexPZ5jhrESUNAxluNc6/8XCOPbGuIRp/NynEq/aOW
2bcNVpHHz4vUbCqLydK00MsLRzIps8A4juJXcsadcqxqdrUp+n+8rRrNdKYcq/QiZSCggPWFusVp
n5+he7iNcRs8kiWjdFxXfVhBaoqXV69gpINThwCUel0nKzm5A9QE6rRsO3yZu3ko8rpIwQP8kioU
jHed9jl8EsegIRnLodexxdM6HEEDpubCkJ7EM3rzthv+iOd3KNTag9vy4bY4Ua2qUwv/bkjiXDFU
swrfdS/5zvs+XYFB12SBK319nAQ1GbuNjWqw6NQ8kYyN0B6dwsXR+L+wFtUr2kZHrvFhKkbnf6fE
qmKxCknEiJWOBfpSUhyWzah34zFfwmbf/2pRTxEkh5SazctnAx12miYpiEOkmzn9WRL3UcLdK23t
LLvGiHyzS/zgDf/l+S4UC0+TUddwDqqMK1NsSDKrPm6vmbb4We7M4Dmrdgd3+0gw+XWIHbargm2d
KS3UFRH/oYoi0DCg1/QA6VKmXvyOhkJCDhz2O64TXT9++nTREsmzP+sjQMQ7wff21Q5ByWJNBW9d
BfG0mn+e0WNjU1sK9Y05Hc66l3+A9U6VGXAmYFn5DS9GtMsPzAKYfPr+Zzl261ExvDU1k+GPBMD7
JaE/36OIQZl2dSKxwzPtH7tSR8TjGIa6SHc4timasoH1QbOKHlfmaJa2hIdTR++si9eXw5t3MCMO
nhAm0SUQSEKkNkNsO7yFZaM/GnjrRlBBT1X2KYI0ug/KzWLRvLIzJij1qIidwEMlwqtRwOppPEpC
QQUaoVQ8CNfWeiHf14D3+L6O2LP/eg7PL8yV4u1CIwg2iX4VzpYb4j/03rXsw5FVbsVbLh6Ke5k4
2WKWzkBuPE+22w5RU0L293cnMKMeZ4Re0LEhlTxqJ/IUO8nx1FaorFCEdo1v9VO9OI/TUbhSKk9p
X35+cpnaF3jYOHjr1ZiSqUvGwgk8k/1dlTAdgL7UwKnknh9dVDhbgXCAeVXjjoFVpgqQgS92D35o
Ym4bzxum2nxAY9CRK63agP03g3ot6Zk/2MfWNuAQMKQ0VPXOXW7UUoCRbcK59q9mPl0Be2IKbk0+
ZoSfHxc5VlaqsKvB3FX6MckX/lNUd+Z+nxlKFcdgb43/O4atTl2qfwLVlFHuSvmgBxD9mXdg8g1p
p67Ir8OESVGQ4L8nwrWb5kalooMNhBUllJHn8ssA4/Yoa4Zer0U8ukvuFphEUn975U9zl8OJuTLO
bLjO14jYgdeWxvFnYhiq61yksPTAB3Gg96AF0MikMAL82JLIVmwy65OK7bPuRBLeJZMkZdc8NO78
mnIZ632QjKtIBbv9PqC3QOJGsYXpNhnP+OcFoQ7lTy2uUEUBYn+DrET3+C0Kzt4CmH4FF9WtkaMC
2gv5c9biCaSPdykg0ffsECx6ocBEL37JqIosJDC8F/4ukaIvvFeVlycokduaX/sGr+zQbgDCZORH
2W/A0d1okLtnjAETl8J2tbketcWrvflwTQzFE7V1jz19yglIak6VvHqvS1I3o/AvwXhbKVgBX99U
26V+An4HfvD0pVnL1cCJuWU0bc/yNOEsjUWfMQOKgUsAzBZPQaDyfXiznsaKx/T9/Mhb+Ux6VdzH
dtSZ4LbDGOoK+OJPz/syRzgY/j4aEo6VO8DSSUFz4p5HWvMcZKG3ewLwZpEjBxg/7Kdmq2Xp55CN
iHpMcgznidYGKCWo/7d87Xfa0OWrQ8jfJeacbZDIP4btJ5PSwFXA9b/4DY15BotPBRQB6bogN/bD
11lGz7AhGqKoa6mNQnA4PqSrumz8iRWG7nDrIBDPyKmaAp955KHblafzGgMtu0vEbbMgyTJG8Bcj
BwBsizLUKh/R79GCbv826d8T54g3VNy2IhgJ8mwBCKW/9diaCpK13IiJ6ijLN7BawIl03bYwdOzx
Gx/Ft/5htXKosYLZFmrVit8Id36c6+HWHq8Ddd17yTpZzPzU+lLuC7Gb6uWq/5dK00GSHMbJKPta
reZ16k6HDq+6iBmrHQws3h3wDmcgmOiS1ot8sn62QqCGOTgba4/+BevIOCg1iyIFfe9CAiM31qSv
B8oj6B6BYKDN1pXYIWFmofw68fb2K3uRypSjS+tSTU6rtwUhp37gvCuxebBzHsWjA2RWVYnQDLk7
DkAs2UOFdvQMo6NbFQ+YWTiCwhj90u798mWwdPmxmrWUeZSWFU/2GjtXWfzTuntPKOok2R9Vdsgr
QMGItFx3ollbYD1u3EDXge0+ZyzjsNQrT8/yd7lfB0/JxgpHUKFRZVRWR2SCZerBJLckSVYR8NFi
ke/zTIeGEnO/7nzCPy9u0RThiVjRiDSBbQd/wDa2oUznbI/cuVJ6E4Kuck5gYiZUlGmhEB/BV+IY
fpjff2wuuXIViuIA0US5szNnW379JtZD7Dm7F0eLGsBy1NaOyfQtbwhuETBHkZBt6CN0yRnsA5iY
05cUGIz46XrnSb2OVbRo19gRKPtm1+ZuWDiOpezjr4zDoVEGX967+ztToS0vcxZsq00/nNl+pOQ0
ivAHZCHHa+L+S3Gnd8hjVezvHRd/kDEhHQALLcpWQ6fl2VTAufHyt5CPMQXXpD76mZ2UEpDrKyQ9
ktr1g93n1glLOKNl8ddnfIs6rNUF0CbYhG/ShxYXh/iDJmLmfEYpjQeMx8DaSl0V6sUeNjKXJdYi
vrIqqw7jfAgP0rhFlxDbKslMJ7nlxQ50tCqg2cZBqTkAaipFzFIh5+BkvEW7wJL+Dt4G85jVkaqu
9ClhCEnMsVRS5K6YD+JLMWKQPl+F2AmA3hxUunZiVtmt8uje2wfQddgIEY5KUXD4krctqW5uUBne
kV/zhXc9+zbuK0bCD8Q5dBFYcTzwH1fPVKBef4Kc/W/sQL190WPUZ9YoUDl79eM0Ip8Ggs9E2gon
hTuZAMak1nZA/MjJ5A6BYpmLRNk8g1Nf/PfeQ33HdhyCu/NMnSVVcmu/KvpPEQPt8MiMh2KlmgJN
S3W891cLUDA6ggRTRUqp29UJGxZWSDGNEPX0UPS/MEBvjEcXSdNUzIFOXFTkQnyt1YbLFbg2OVvT
MouR5cQdz9AuCSkh7Hj/ysDV7SXj6mnmM76tHlhwJbq2nPwlEPcLa2FNQV6wSQKKluiGWI/UtpPf
dgwpKySZ70NqWJrtNNOFtRyNXHy1YtbvSLcW1G97KpuKLM4CjuljqKCeBvXeiuW2HeW5yADDLaWY
z0JmO27dNNtShrSJMpordotnvVZdLUddEX0BvsSIqDD42ePnneOasZQq60ta43/XbjRy5B/zoYFf
FHut4q2HLx28/7kuMM7R4JxaaqoO6x8IChCmBSaGYUqC3KvXcufroyW9x4STma2JH2kMoAQthmQt
OaR+yXpQl3NSu0B62591lf0Gqcf+OZd6MxytquSK7KZM185vvRg2uG9jTLo/utXBaePg2+YH9ns+
lFVVhbRAdJtevZVzNUFeh74KrE0i/5fHgX+JJWAMEHDpR3X+GoJ7sZiyAsbYfzYrUONhh2tUou4t
J9jdF0oJegt+YpZ46XrsTwa/3O5fNYj50W+ycuZ3/BfbZd+Syj0pJQbecgE328v/Oe2qKeJBS0oF
30iu+V2eUpwpnPEwUZSgQsgU8fJU+G4uDqD5CycfyMmgRvoq6MjwbCM9BP6vFwzGU8kjxrrYnpvM
GlV/VXJ0yHQImfLE56iJdqhgbcprWZImugwQZGT7Vau8j3PQpF8hArkuewqGb4gPBEMUlp33tfal
dvsIpAz3eB33pViKX2oTCAcbiKnO2T+fu3v1kv1755iYKLD178JzkuCkykEA0UHOUGrg/rwZk1+T
Y3OIoG7h/i3xGx7qFXytlZjIuY7AsU1aaKJgofZw8twrH2jhgtvtP2NlmmSFPaXQ+6HcQb5dpB4S
/Yf0jeyebJwdp2qy8c4yKL4nefLw/acE/nsIPgEOD3QaWzMIuof5o0eOcWBD2PFpQRDc1WNCq/K6
doOBALGAdjdiEp7pkVlmGxG4YZFtwQPqwO8kLHOPMZgRS4cB+bBpD+Pb51JcHnsUmkLGQOYO25pP
GlU/3zXGvG6oAop2nHtjVsTrx68vNlARlSc1OGiKkSSFg5HnnKkoc1P0v7zB5RbZ6WnfDtNhQ6Kc
JeSeYbHpnFHatYhQJbkEWq8ZQ95wxbgYPk4CVu6XwOkLd7JzpXxw+H2Zh/Udf0NYXsGZCKvtwUfw
3wDRwoEsQWX+MnYeKRfbMzMekaTTbdOemi8pDTW9b1FeLXk6BR2LQmNyfivzQYQ6OsnPlwpaAEGm
XCiEguFFBlWDcCb6n/6f2Kx+EMYW1LRbvfJayZWQEAe2Gdy5FS3ISpla69HDQJH529ApLSqgFRPi
7/3hx/lj9oF77oOD4GoKs4ePTcKF7N9B+ONQay9wTkfcFoZMGpBy5P5LuyDsu9SNP7n2YvOuIV14
qJmhZHVXktGWSXp2paL1yilMoAY1HaLfu8pkB1+U6FgWTa4otDDQk5JiF3zn4VsBGDC68Py6HSUU
jU6m6T544lmZ3iRfzhKLhs16nB7RRMD20N1DaotHLdlSsrbPf5V3uwhWBycpj4oAyuyNlzfPNkm1
fE0smJl/QLGjCboUfMzY/zTVlpBg+D3Q0WtiBFRIi6c9Wtk1jhmwvozwPe8y7juFDJ7us/U+wGwR
gJe9AWkzWBGUTCscRghush0qgyy48dGNXGL+LJAZF7C2T9qROZU3+bwYdxQRSk/wwn2OxCMYH2lw
3vYq33pwuyx4VWfg7odmZQJNeQZT/YAN8jqncj/vt/nanzb/IO6lRAaklUWfI/Das2mywx1xvpbP
qYgy1j2mzWEak+IJ31KCBjFzzYGCM879194ylA69S+qH42VW0CYPkYbQ+WvTecK772S6bF72roaG
qbg9k91ekaFfibm+ItK7PW1NjXNZ+RPZwc21QkYQVepw/fZCFd0Ai6wVfnDnDVPAyA48II3//lQu
9oIr/hM5xV3oIRZHxbc7IR6GHYpW+qsaMWDWbwHHyQsr2KNjM0CkGNyGWcaNdLKgy0/uYkF+tF1T
tuHE3Id7O6dt/l9WOVWWOAZ5u2cGDjircOjyv9FJWFGIUkf04n0icFeLkwhZFR9NoNXC5g+VvrBN
95iQ7IskNdEQL5HwZkp8haj6h8J7n8mVQgZRWJb2g7UN8HVV4+wWSPoTO0DJXLFeYxohTexfwyof
SGDpGJXI3qaR1oDk5AJNWGzJFfYNzQ48M8l52DblM/QLLYdtmZAIm4qEh9bB9ZidEn1hAl06EE/l
MfWpiTq8itDrHP7sCkP79Jd6Rgo/VwOSsLdk++Vnle7DnEiojvNE2i9s9ae/fmw77KYjgJxX+RXR
DtptQkEcCOhsDW3+AYTuc8c/02hhcll0cO36A1hFp9ofBcSHAfT+pQbLFiKTbW1w1QDeEkIPiVhR
uN/vATeoK+gVB+RHsCQp+j/56K+8Yypk3PxZBYPT51UDfCz5FXOovKj4HY93t5KIYfIn3zEgBAdv
HXJL6IcdfBrxKF8n+htt/l+ePhBJKf2S4cG+jmtA2odWRkgGtjNYLQp39ZMYBgDRE/nH8gL4XtZj
pX/ALyINlYjweyFJWr2gKO4pPVsTyFCvq3BtEjAZ6H8MzHXyPvoTxAvwrsAeyjnCZTTNBKXvMvZU
ghZqeFCKN8oqi2qQK9+f92Vmray1dgBUqaP3H1bXc8Fydlp9RK4kGfY+Te1BON7gmkcItr1uI2/Z
emmS5BsbtlI68F47EkhOVFYxoxhFdAy0Je/4a5RfXUfp7Qw/onT2yJW9Fz5O2/3kYgtpc89kFbfj
68GolMpXhhzqwAOqkU76GbnzMjarOksV43ygG2n6ayqcOY5h1LwOr/KCBxEb3iWhqrx+eMm1AwAV
icDSd1gEXQpR2mSQDFgaJGRS4ckKuOjrEoeu0ai85vh7M9Zsxkn+otpTqHVP1Ni7YmjZlIct9y3r
AIjdirRDoVDJktewTYUL4+CfuJ8dKXAl2xdLqw42nTohUSvwTpL+P0JeXyvDA5KVE7EVSlpx5EDX
OSX8fELnDkIUlaxiCo94O4pRtnq+/RPKl17o9Eevc+22lQXmmYoTIW3P7qzuxywy7wpSqRW2OrWU
G6YX/amvC/Ny59yClM48lyu9JvC2+9Cnk1+q64f2W2lYPSnmafIAlpci2ddsdDK4eUxVftbkH0f+
QdpvUoK2lxuKKfiK77oCIU8aIie45qHKRj0G2EG/k+ToFjA1JakIcp7zBzoE0Y23r2LFcQUqSxLk
urGYPLcTFVhg5CKnQy8zLZrbVKVXBr2CvGdZzPHnxph+NgCBj0xqgK89eMFkQmu44VjsMcRu9UlF
dkAJXYTWDo2Yp+6UUovsrt2/BN+Cdk1xGGcVKq2nTSJYNgJ+rtnwPqMP6Nfwn+qQfna97lM+Um83
3AihQofP4wkxc+VUvaI2BHif0iD6E6kxg43pkUAve6wX6/53zntk436cY4RHNLv8w2554gJHAhMy
nRrzlUFKJ7GztVCMtUS8C1RwT6NmANXeOEVBMB8PeY0bTuvWwBDa1ZmAfCxJm/8kvAwlIPd10Pep
cxhSm2+Nx05/VUsyqsUsQLTQlYTt+Irf5FP3KZOMXYelKlqDrqJXvcJKFT7eWx7tiHhv5IriueT9
zj39CwdR2fdmf/BqK/DAMyynahvvvHcHPMVv7lkwbgwq/rDpc+oPAQJRwwuEQM456aNQyRgXJMYE
UzDPGkWvYdTFU/SLDzIMfptfx4HnwSj7gcaC7S3F7jr/fPH0EMDE4ebJ8Zv0CJHiHyxTDyplKlpW
zTgjYuLOdw9ac0ftNawzM88W+rIkYNAF3mluM6twGOy73PAB1L13pcUVfQpfePG5/BxfKWOwonM8
slz2yHb1y/PwS8679qUZg7HDUscXZPIWVmp/Q+IdxsddYGiF2FTfksYZbXble5EOJNSUgHI99b5i
V1ZuOpBVN5q2gxR2nhJE4hp8TLHtprwYTkffYCPfLaW+i4wQsAk0XONsqPQj2p+EhiPztWQNzavC
wru+/72mWjfzNTIkrR+sTJApEa+riSoekjKWnqugd6dQRyRoJ6DtUBjta9qHo7Mt4YfDKuBqz79y
0g/XDgNhYFjMjwYZX0Caz/xIz+IMG8eustL3dWeHHTEef4+SJ/zxtRzHmsvGXvOWnyPuae4XHKus
G+xNC8ExfCCeeNNJ96msaNjvHkR1fzmSVafw1EPylSBcFihdVtbylEU0BY6tHAX9SlPYPTd/Rzpl
+4p4XujE7OtTdpuz9oG0AVE5672skz0Om8zsFYpdunwQd5Jf4HjQ+ABcg3G76Ft+wHu4PTRyGlxB
j7ruTUiNv5e70tZX9Xv4pZhkw9QOUK1HkjubAFlK/ajAan1gXmABibmeExyJaE+uuZ2pjEfc2Wvs
TY9pLNd9JemhlwZImlAo4YCfAFVBFJys9RKptNZGyg9ByM7EsCxn7Hq0vOBghQQJcdGNOGiPVOWQ
/tvPnHSSB0of3LYWBzACgJTCAoppRDz/RG8pX3I4nUxPwWxhAHdRtSxTKQYcVJhMedPsiqzIxTjQ
GkOrM/1OAyGXWoLQnZuTqJoYRSEr73FC88xzyx+A5ALv5u++gaqdtI+HQ2goyf7Bg4V2obeLACNS
IfQUxbJnUhPLSH1oHN9cbwK8eBFwYKWSPNrTYCh4x8FFhqPhn8jXoSg4JvHY9wzEvOZRUx9MInNk
CmoUG2gV2JAD/TtfAm2/Ro7jJn3L+Zk2U8HIB+OxwPw1XXBked0uj4BRzpRV04DYIxBq30yGSNAx
KxLcr/K3LJtkgf2HiiYLHjJkKxeYyqnoBFJ1AOvzswq1Xg8DnsufvFCXMgWhwtzqbMysrvWb4Kz8
C+eHt4PKuXL3LMUcPr+sIP7i5UL8IEU0ZBAf04ruoIIT2kZuq01BTVSKYgx4Sy9Wg2nsu5meNtsQ
nDz1UjjYlOGTpd/H3BGFnP+lGf+sr0G921giM8T2Oj4x2H5YOM46r48IyseqRN2DlkpDNZvfIdGu
jo8NhVzs+qyyGjvQ+xMkMRio3W6CfzyY5Otit7Go/S0vvM2WcYCm3wAN4jA8jlW4uWR/A/uyG65H
5AkB8n8ShCFD4xWlszlgZV8G+y1LH4OchyQmFFz5GP9SixLuMB/1dCk4uxQMKZKmqNKHNum7rLIE
e+TSA75BmpR3lJUAsVmSTH39tzYNnhlQU1/+0K7nIID6BHJazJUzfrdlRvjJp5Pym05q1MlgP9GG
KHJorL7mf/4rwobTEMq5T2qoMoxvmRu28QE0XWSacrdQqVAL1/sF9eYQgEkia9pqNY/lJTp4WZ6a
gqG1ki49R25XxvPOPiizJeYykO3f8jJJavMkCZXxYHL5S3TB7AYZw7k2CpYP8jCe9MKzFhclBxha
jOdjzVAC499zVQlyTpBbkJafi9gYsaDmmZSf760IeAsjsvmb5Cz+y0YkOSfJ45EBk5FuJdEWADEV
5ZhKAk3Ivz1fgxbMzGwci4uRzFiBPss5Bp50ZlykIyhPigMptYPZ767JFJymnZYPJycUO6wPwn/w
tv/OTaoe4E4saty8bQ+XJVh6Y+TTdaOakL9x/Infh+EzEONP2sox9bTFetcPXPX2N3n1hzCSh1+R
TgzZvnipvZ1FQ+o5R59aUJ1J6l6q3NAxZCKgqrnpZYyalqakkxKv8JAiKtjGyxFeZXiuiwlCXLfM
9/DzsskdbYhQGmvL/2G3g43GjSOJy0SaxFYJeHglgTeuGNJTp4OD84OiYtKQcKSIURY3mkxwdOv+
yPigTTIkQXj8iztP5pQbl9Ei15DwfBSHtzZBx/HLGSBr0nHWV6gq9TGkWiCD7Fe15djs3gE+RtIo
w422qeiHqjM2MuvnwRacLynXs6jQfh9xIiUS85D3+mC5MDA2l0C+mfgFh37+CynNt17mMg4eE59R
LtUH1IATTP0ArRLLvgIVRXWNALQaS+nPHh335K10YnJOtFqChDeAhFP7E7+c+RA+t3JnPaMoGH9x
hRYpTVUYgeYNcnKXbAkXrSU3U5t64lhBqZgmogy5M3+QgUlljUfOOju/WPRcrR0DLmIs4IWhB+Wi
9cnzbUfqE3GHRH4S0gmLC2MrsCAKJ2XDIYqGjxHfLQd+UnlzyPdSCpi5WyKO813vmZ7sHAEVkbz6
LkyTLaebS5BTVDv64O4o55AYUJxSrwMq3axPHUNZM42Ql7nr08obweMzFHrrZYQxhDMCahYQk3gj
koEeb4e1mgFVgMjFNAT/Mc1nkfabRsATyPDgZz/Ml0VVY2FGFvhW8Y08MlgcJbwlV3T7yRAAIaf8
DpTwazZrnV+aM4XxFLnP4+R+H89SFtug/XnZvaMv/t6aXQHMNoh1hoQzs8f3/lPNITCvCQuAfDWC
XVCOT80O3MZzdGAiEBSF1dfKpqclsNGQi4Xc6iEnzBbQaXW7ztc2cTItsDH6coP2hp/01TXI4+5c
P4ocuBEyfBje9ygH/oZwhbCL8ZbqTh++T4BaM140BLaRdaCaNJJka1qfsLAe06kE1+1JFty3NWBp
Tv2VHaoAWyFJ/1g8ATJgX0GccIdmJhOKHDEjKCLEveugRC35hlHE0Un7UYLVRCmMcgAuUwmXiac9
tyB8d5Y6zQGQRO0Uhri9KdU1SvDhAECtL/MYsd6p44LiMitp0xoG7YJvSd3i9ppowGBGT7oryLSY
kcokT2AU9W4KcAtL6Z2Hblw4nSQmfY8c8kLyUCvfwk2/9qFwrRZiUyO4lSIb7hWk4qb26Bx+mauL
S4k0CnQ02fqeXIaxOZ0eFRtX9eYzso8YHyjlY9FuEIUJvMPeojwp1/Myz2CAAZcDh4rYFfReHRFx
B704iTPykq4n7ccHHVUAIR69VjrWa/U21cWG90ZlUmRbvzVFJdSom/FdajfWs5jKAKQpzSg3c+BI
WSdAzSsUTiK+7N1FNqrMAlJzgYi6KkjyMRatDxdSdFEB5dQ3wQVk2UYBAcjOTyBkU9hb/D7ejyhl
okXtM1DUQW8YKY2LOS4rdGAxe+0cLxY6xI7BvLaypk7imqCZv97pNsbAV6LIcGiviLz/mKJdbMrI
Cb/z1WIUoE0vc6MPtaDrMH+YdS/S3bMB7yU7ZUjgwDDuln00iK7F+RQD5wXj6thLRuy7LeJjjTk0
3PQOET17rKRSSwFrd3vAX1FYCVUJF/XMbpb3/Em+5vJ7ta0of3eFZbslbzNp8dnXU4Taf015IcGh
mGmMQAOlhyQVo7YGoSbAsnb3lUeyGlHsleQ3k/UdX+lhCJi6n/YBRTzqNeydm15hflqoByJJhYbw
Gg0fdrla6EyKSrv/snoHB2tFcOlwSi1mgiV3T3vlcu4CbftE/0eaZVbxY6tUZQtH+xme+cE55rqP
4O8rocXw+iKZhwkTuZBm2NmADp1LZK6Pwmeq8xb685210M7iAACeacfhM/jMjYllW9CCGqfcScBr
Ps0UTzp9vEUU51KMLNSju/seKnCqEuwlP80yE6/MzO8dV3eyiyLwpU5oAkjbanf+msJY+m1i/bpN
Q4LZ1UijkTVxPQwfqHF6DM6XG+sSkSm4kBnZw5ZsCd/36pzWdJHieAv9Pg8xBcZYNe73IW0WvdzX
2q9jWR/vRsBkUgvctICd8mKWi3OdHsEc9BBJdgx4b5yRaAjBDjwmXEruWbyHKr2VKg64cMzZRqp7
skH3EnuA71WNiq+BfqtoCkovYDXycMO0/x7QT9UwxLEeDsY8f6G851Ubb83a5Vqll9rT3uOBGnaS
7eFiecQTRudev2MK2gD0WbB/kAQr7H+4dwj5SGiYUs92wBPI7EfY0hsU64y9f7BxZnKBJMcgL462
CQQJMchHzVhGh7E61FLnPKy4nmY3iuxcL3OQ1zLVGSNqRCv1UugD1+QXhBueD2AwgmHNK7R4WrBQ
W1I/lJ7fj2cGtYqjt5jQAyjSRNLipWaPJJrK00o7gWmyDNVKrydyADQ+E45+TvFm4h5W1ztmLURd
/eT3O1gyeFwyjzVljHbJDmbYBvRdOUfc2WlSz/2ltuBTnqhDROQYJLHd7mJDgPmfQdy9iRjx874o
ELttw2UK/iGNf4ec8+esLUoLU9fKpE1VBJfJO9NpJTsf30pybKxgisxITp/v/ew/F4CPt7Oyp0AA
Y4yVERwP2XWyX7J/LuG1dwk+HuDEFBBJmMgsCUCHp02NY3z7lWK61bN12MKA8pbGw/rDzPHLMM0E
VAFqtZe+qFmNyjP4lp87xaE4U4PtrVOo98kNKFUVj+06Fy3O7bj7u0mz6TaKygzYbFp6AnVrL6WP
z3Gm7ndQX5ZMOed6GYZWX2ABMlCw8mklswx8DUKgaZEIw4KHlQAH3kc2CLLawtABFg+YxD7NOVK9
vBYbTTRgOdh7E/+SThujaA4MxdsyOdT4QDKj628KLRUUMqz15EmYjj2prZr9H6b8bBZSrmbvhJSp
W0vSyHtQwZakko9NRegNgqvtKCzHGzdqdNHSP/xf3g/GtUksKscHvo7Cby0F0rB56oHo/F8EWDon
P1M7WPRAQzve9bKyOPKA8aG+KE8dFOtg3XEBrucVkbKzftS8WWqmdMWVCgj+K7WJGXiujGIbX6fP
ij9XM9h3ml9M7UnBbuifoX8kvh1zsQh19n8HXPguAkQBS2oKc9nDcIUmWFEVAjSTEvvUxipjvQFW
zRSI0yF+q2VLnVbCNCdssU4ZPse1/c4ir9VknU4wtR60aZnFIcb9JvX7PzYCoV3VcKLYlArDcPoA
KT6xf5UxO2CGyj+ej1a4/+6AU1EMn3LHIdMYIIZTGuxlSgcSW/lcdH0+DEuz0ZR/6CXubksce0x8
tvJuHkBviA5dTl+m6Ak6V1euQFT4chyVenfm5nOfF8xFYolGsmGI9hBIS4JJg5NKDr30SHEAOWIu
kY/BkthD3LSLpJfq7Ca0Wy9TIhM9fMjYCDfDn9q0ZL6XlonKZy+5+gxr65PWe43quEf3go1Jou0Y
5UFnATSBjJdJc1gcT6rXMu4ISgntW2QlxdT0bG1gYLiITlT9nVijsj6f1cxnDlHX6v1gpPImI9BN
JGZGHycGcHdnoOv/HvAoPLHLCZNHTDpkBhF/Z4FB66Z156/DNIXCt80QZG2LacfyjsMEul0Qf5U1
ZaHX26gciPea976pZI/i9XklSOj/QO2GkHT3ca9zxmWW/TpbPzSIbC7taOtgrrQm89AIxS+5bINy
OOt384zEJ6xtd3FBhibB+uEplzoAe4XSlHBlrJkJRtqL925GRsm/1ELgdBLGXLf89+xbXhEucjjD
poWhIbqOnOqXNRW0M4lEl5wQWfb5CkNRBmGlCSqA5YC0wZ0rIXlGnk1O8DnuRHxacrdvfLNqt5hI
7JeICqZifhHyL6KTOKjSpdmTIBf19v/vAE9uVu3u2wpvhXAbFrsovl4dTQJIdG4bseY6jLsBnMuw
9Wez4Q6fKAdbMPpbHpzh3H6qmI0MQE4qbwaF/TMXSNboGJ+hxj2LjKS5fxYvLBasg3I8Czw7g3JZ
5/qqBWXHrbzp65RDN95NW4IltOK6jENiOr3qFuSQqO4iUUHaaETgHwegJdJx0WAo4itewohFrKib
WfRbS+WZf/8e5S08TycP/aJRmSu8Bd5HrR9wYlofS6rBQIquYsjsnGXH2iF0bsGhtFpiwj+YgxYs
nr7sxt4QognkJ6r+ddTCus8aI3GPLk6afY0YLRwyd/g9ZlcgcQLRzaNs8YqtZqePaqMWhBKBOpmu
mUYgziYbIwwQJTABtlgo3HrJ6kxngSz8LLkfPAtlYD6ErhxXyjTHHztLCmrJ2cd4QL2Z7Z4lhdGv
mTEVilEvd0Q8bdb4+bpOpxXBU5oLOiU/tK+Hz6kVc/fHFUm0huHm52rJ+c4cE4szT2IWz/WemErk
f/Ho/mI8ErgZ2vfDJwxJ94lw8dTd1STF+Up34U/VKXh6Op+DJypJXVFMDwgxfGlZZfY6CPrnjZIw
6n8ngiQyEz7H9reuWQVfyIsKE/CVIeXuxYNhhMYVezNE7N3d8uVx/uWUg7G0JTDRc83Rp6Egs8PE
wNOKuH2k5a4jC7Wb5j3hOpB3YUSo1KBFy4oSt2uF7OXQN0jpu9VRQSJKRkJw7vSP/vXhs8yrxld6
SHMo2A0U/VSyCPHhTNBKSuUnkWh6mN2NlUgouuQUrVuOPpDFMXBAJlgfBiXHb//mB/3hIGvdqHlw
4ALdKVBTty/JXeZ4/xZZ8RPhP1zNCxV8vagC6sAmt7wV8FSkRsNWEk330usmQtG9v76zIOsKISjC
BmJydhAMqilUFUqOo3094oKyxR/A883LF8WH0Chwu5vXSSRrVCa4CCkth9b3mYS0AK9hwJNGmY49
/1djmoQqcIMYgUJ91u7NzGt92feQtw+XR2WpKFId0Ng3/CpKuWHDOeTuhuoOC/FC9kQI7liq5pSw
nt6JyH5Gur++6v0kFNrP5X+NxQNW4jrzuJUDwSRGMEYK/l+dp5vjKqkhtze+xg6yas/1RwpDXbqt
im8TBIit4U/WQCxHottlTJw16HlUwhqxz2kuc/v3dEzlfOkN5VcTVGoVdLNUv4Rft+uyXvOgLf9G
AH7eUz+ZoA6p4KyREmI97ADtI/oDTj55OXJuQ2hnzqEW5Ik6oKsmfi/H4Ke+Zs+JNhiRBLXoXSr9
jZrF9+m4+B0U/D37jW20CDzlx0O24/DwIqbYRUR/Ugnb1O18Ht/ahv3dbeXjJu3rRKhq1WNzap+F
IypleH5gdfx3sgPXlCK9FIG6C6lYQb6z++NlMVwpsPZM+4Aj4g9mnFn+KP2kEoe49+7qz1kH9FI9
oLjqDS2b3jI6ckye5rZTcPkaYtunMV+rmQAfGzpG+bAxdWUxQ27iy3KJxFbktVfEEjQi+ucUEcbi
tT1Em2iTK5fIRSHRghP9uxM7GtrN701pFEM6GoT7d6GL+MeGliYBQpGnTen1kka9y7B3pKTuIona
mpRpmFp1JkT9tbSoNwo55ETJrBuYc+PUxTmJ2OEGDXwcKpLyHlgEPNcFvtRs0bWlYNroxWOQph+z
6HKZAEYBIRt/XfsOviriXrWWBUlIYQPIb6KrFS3ph78CX2K8CQiFPILqwvYdDaiXywsUYBYZ42kY
Ahlyg88a8/xsB9KIXxKGlER2AXdqWusSlssmXmZRYHzuVIjJiXGVId1c58pebxYaDL5dpLaY4TiQ
uRf9o7VMFlU7Ny74CrxWt63z82/FL22HEI0SRugM451Zg2kOLfc7n+wway+OShEvgDU29M0PxkKu
K0WC1Ufjk/9BVsyyaqPuwGPQs3bM2o8w9isxNhk5jYq8mLeK38+BD36HDyR3S0PsrJXaXq3EuFo1
gTY1m/rSuXfpQA6CvwbVhkAszpdSR7SDtwykIb2s/EpEXNWOIsh8OnZlgpayO+9FWxIQk4EsOpOm
cogv3Sxe1WJ/yk2uSx49pSl5J8VsBp7C7ocWZCCqYXRfDFSJUm4qktESocIiCVtYU9qVAj8kcAyQ
FYbwrow70BUECAqZN3wnqShiNOAASTouujf6JWOHRRDKOV65MbejoXqNwKldxc8IDYnoA/7iBP4Q
KG7W5Lk8A3Aw58guFQE/NdniSts9Yc0rocHsfm+DKXfDXiXSlnGGpNhbuH6cin8AH4wP1HGbswdF
jnG2a8gVE672TZOYpPs5TRmzSJODRT7G6Kw/rNiA3pgC5RKbUbWOG9XWKp/IORmrCAHV309JLyih
sSM1Q0DDsutM2nO2BRNtaUrmx6LnE6ORas6W4MKJl+LRC5QYMXtNWz8YVPyaPVuSs9f95uY2Cfai
XuFLb9VUs7CsbO4r9aY37NG7za2uN2xjTPq7sY1NKgyD0pNHPTYWYAbDRklgGZEApgc3RQKy5ZD5
+XmabNJyb1t/OBaRizQ14x+xilHITFfrJ0IAFjuvOIgUsu8AkPE0csl16yZe4QehfmEh8oYGyLt8
69czDUSI6GoGH+kBRA4en4Vt2UZqH0Kc9K6V0/CUNw1wxEUiuy43ueEmSOUxvSD6wK9Vw57fMCgV
tFy9YEeMHeaqruGwOxs718QZEDS/x4Du4Wf0a8s8PljGTi0bCWkZOwnfI8n7wExlhARyQXWRQvJj
yDESkInXCB8t0ykXa9p5whcHUk5GuYOBkw40SG7+u3YE1a6MjQ+JHVOPDN8VEJXaR0GrK6wqVJFq
o9LenFsMuLKVpCh57XKpnS/EeaQgFFiOC8DDcNUhFLkRTf/Z4mWqiivp0lhvSbf80odNlWnM7BQj
rEtHbd15ea8IaZ9DvSpfqiB5auzyMsRYUlcBz2njuUlU8pgKtJcLTi8I1G/HKmotDjMABFVTHzVg
yuWqM6kaZDZ3sSWygRvO8APtPwKk6hAOsGm2CJWee9BUPNN6Slsd9bZU/H/WRhkNzAn38YFfKPjq
U/oA2Rl1F6hdb3dqmQt+jGTEu0qJTENHbCbDOER4HhGDpwTylUu/RhEgUWoTWShJB+4Jj4yl6dR1
Tn8KO2meMYogsVtSbsEOYojGJ2y3T8WHrMriqK7POG3rpM+l/FYym41ODFu/PARyJQAR70edKN/W
DL5o8tFGIm6iPzKJC02SYy7VgE+noKB9rrTwUx4WUjl2fIw3tVb5hyFqVtTuBmxpYipyNw6H2HWa
i3uALuG4VTTYXf6jxzcMfkUsW43EVlKPiKHdkangw/1TGIcVWfbAN2vHyne1jsTI+bP/+JGg1w1Y
ezLYYKyCzRMvw1buhVpK8pDjXFw3zfjDOFm45Hwn8zZUGGs7JOnbQYYQj0T7sn7EuqmMdVoEufZ0
HU7d4ZY7Dm6uQWnfWGPA2Ll89UuM4PeVr56ARVbdYcBhXzs9azJ9BxzOoGYtKjlO7p6fJ7Uu4IiK
3KdrGfqX3qcUfX3v5RI3wSi9WHJABe6byY2IKONZTW/OeTd2gd6D4jAZi2LyTtgvHRCcditvQCze
fB4cMDSX8ig6svtyjr6V8Zr57utuFFzUd2JRLeoqMXD2FBUuDSb11BZFhLumHRhJPmqWeosEYpWb
baoOAzCI8nFSXuRNdgEVmo+AoY7c9F1nyDztfAEAIn7SJOI0T61wJp+pKu5QYhOve6GRLeVqDDaz
kvpaKSwltZPjpUU403NKZjTclfiSf54erz1vFfe7hrAhE5LqdPOG8rhak6EXefWUWqfIhv5HZbHB
PSFMo85tk8Kx45Io2rsTF26aVQVBB9OuFg55LQ7DOLja8QBmGOWGz9OhqqARx/+VcQdjbmLpwkUF
gjbkFVUR3MKo3cTpgXOOsUiYsr7fTf4heR80/M7DE2fS+1ACnlpY2a98s0pRiVjv6Qv4Eh/m5J2Q
7mc8A3lB2V2ojEgIkaObJF+R/0EI7vWkdsnlt6DlZ1/n7PG442H972lC97unmXdZSOHIEgj1Yxkw
b7J2l8WqmL0HlbmaBleiE225FbZvDHytD5ja3F/jvi6gr72ij5JNPaxb9oUOHsEXUwzt/0dvG6tN
cPZTJuqtTFig2xLsp/BpjN3Kmd+CRSjOAvPmYgbqkS16fnJ2dZUHYRbg6Z0uwfUdJCT0BJKoeqp7
242PozwxvrjImeqIxyE0+jDnNeWDTVydvsbJrDWQqxR0relL3jRrdHUETKfLqS34EHOm8zZUGX8o
0vAbYTsV+iXj+4IOcBe+XCMfdiWy5H/wbhFjymmhE4LVrU5zjduipVCqnDFo7AYGQuB74cJ6sUHt
DX1caRnMBwrfBgDJlDu3FinksXCqWOZjr5KLxzszVHPRiNMAWVSu40sbNxvq03kN6knV3JV5hkL0
UXt1FcTLQfCF9OPX1ZWAGC53LoKFn9fJ9MSU2c7y7UelZvX1aye7AWJWb1uqt1F/1KgfMQy2NcJP
jcEgnEPQgKWC30ap/HCBUAQk0sUK+/VWnEKsokNXBMxI8LcUv4XT++bh/m8wYcx9AfQhOVj2vTOM
Z7cMu4mrRb5YiAx2F+Ii50seSt4SNDlq+oyAYriN0oIeRyVRANgfcnQEyvSrfepo/tPSmdHoFCXN
RDVGIvVqgmrjkZP7wRyuEGtn5RW2acK3/lgImn2bygbyD3v/GOqvvD4vM0dVr9D1NBfc2SJcEeBV
iimMsKYWMZ11oZjOxp2uRY3bEgcDc6L3yU5hnE4vkfDzWaBG1WOZAVJFJ+eTGFbDhCyLFtCmfmgA
AnYpR6eXb20fFZ2Au+WQGizrQNUVngj7a1VUtfK6isQi/vW78OJgEpoo13v6yHFcvJibm26s6woW
PsTFYNuT0wKBLq39wwF0cIatyWaSlai+DI/Ul+pad02ZxEQHYBSdjpaNDIinIPE45h1TdEr+24I6
DFjw18Pq02ErpJn8a5z1QdpqFjVTwDCfVyENpbqhyo3ZLAiLn5zmKJWQDZwoBUZJwsFx9cWYE0+z
qrfcqNUjI2RvP5UuZTJLBRRcm1rvuQHWqz4SbSBgvqDPlWzY7YKDfaBiK15VCAtjDo11VCQh4LjS
ZkY9rBd33ckmhHhhkii9gSLDNQrtP6ZS9lUUfOtI7ZXKs0xvycoa8lgJYs1xMQ0BYFKIxhmls8wY
qAMfHLBHMOBeiwg5Riv0QobgpdwSfXcO5s+NLQcRv17fb4L6btUrkVC9ptheEa0bHod2vfIUBrKs
R/89BFUCSkQx1ZfJGKwPsC+IYbGgkZjey/yKL3z9HRjfLNE0F8hNMcfkF2aoEWYkfd2vxJ8AWvAs
8z2gdvGZdvmclPA0U1VkqidsrvcHyT3NPekZZ9U6XXsaOTpjBEa6HsUAxC1hr8g7hyvzSXsmDLR6
ZfVtkSYtQKozgmcowXF+MRR70nC7E6eEooKAm6gvLeOe0vfptHTffOmv45EspHBWboUMtSQyiNnj
p1ya19Kd7f2nJA/VvONYnYUME1hJCeJUfO14SMMLgKtWiqw3VPk64OSsO4oGMPQ2xxdvzmwGECPw
cZqZuA0FFFroK8kqmt/nGggyFdjwTJJiT8YZ/camLRiGzF8PniXeKiqjuuldYMBWOhiwNMF5G98f
4eocJyJSIuQUsFvXGhiVwGmm5Fwp9FIgfonEnnNxdhDBN4aAu8w3askcnYdhYbUyBaSFVnv1a0Q8
HughEYoLvmt9xbTTB0GVWRnkBIDprzxfB3LgA3LnxAmosq4amfZTz4OC4qNdbCxtPxzLdu00BPEZ
wrNC5XaVAzpnEAbV/nloo2rinWR8gnLaflfpu64FKua1nBb03RPAL8FhSU9x6yPxKkvzX5V77eFN
BQhi3myrQ7zfgoXSsNfViDyukre+CAx60p/JaTI730XjbxsJebbqvrA3ozq1bnGU+ODwXWKGwX7W
QpbA3rR4LGpXxOT2jeCx8pPUbxWT0bskkZimydSteUzg2ZUBSqOjGusVH/9ayzNCWSMtcxUGZEvj
JbDGjY5HpDGTUfOXhvAXIFlcbpfYNS/YsyDBntf8VFCkE9wMmdAlvjHjEL+i4N11uXliqIh9G8p2
ZI4IFxyD5KLZSrCvSp6bYpDsAUY8Jvd2tB3DW4B0pfH25cmGcfHo0/7RlcbVNi+yrW10oNCxNhtp
qYsGXJDIxCjqROnTSKpLuhX0kyJPlQMmsnv9IK2w+1KqdCGEGUtn13Yd1VlN8Qg3SifzHrFrAQSW
z8Lci5OJwUo+pLZypw2du+EppH8RKeV2JFGYtVOS3yXnBe9delD3GLGc18SniRIyA5QGvDeUcOZ4
a1qWvGjIiUrlrV675nFweAdmj5nu0YbVtpoxI7C9EaVHRyUaMJ809owZZ38arSsDWxau2ZYqrhQS
ISBRIljSHbcI2AT/CLIvNPV9cphunkGv9D9H1N4HgOn1X9JGhFum2niFpo9owoQeB8FuvJA5UZl1
fs2RbqegoBCyRpk8kceC5aXaIH7/1XgRRbWlLhxhw5nMebOYSixRgFJ6XHDhDxjyr7WPAe0jvyLY
cZKqT5mYigDZ+eyoAhjqPwtBGKqGNtcPZJiGM+69K6h4UOh0jp8KSBIaivpd6cVrjTowjPErl9M8
5MkxWBPH3zckyBX8B+qUunCMdEHlUMg4YHDMs5bglbpW5CRrma/BxJaFiJe6hi52l7yTAHs9KCiI
awhB8daGGWwULrqpr5pH2LKtJoTUqzjtAlpwDn1cVdRq9SKKnzc6SN9uKo62pNkue56eCA2m7tid
oNo21/I6DRvohl+ybGZNZN1urk29wzGBDnrgMaDaMseLXy3rPH4XKQkLzlC4Ua6iX6YAVq33+ZTW
rY3FBq+xrBmhNcUlqlwrRg5i226DwDuKVBEdqc6mQ7w6sM3L36aJ01joQM1TOUiilgqus6GAZImo
LpPH2fOrCA67yo9BUrAXcIgCYB9OtKdgoSTS+Ut6hHJQ+6sKP9oP3paaPgdXNQdmnBIwH6Fstd/s
WXv80azUsHJw4ZRsDBCn6dB+qB3LgJQt/9Yt9+94LDULaDTe3/fuNUtmkT8VKrUKHL9NqVrGX4aT
CP+EcQGI5z0nKoTWRSWcF9aBKS7IRJoD0AR+snmK2GYHs2im5XZLB5LS59qu8pzJWO8FHoZf+cVu
SXHHWNm+1pxrJOd1gB5D+8OoTQ8ug7f0P+8uITnLmkTFdKkfgWrQ33hd+KJkh+YX2du1MyOhXlGw
5FfsM4TdhCsBALDZ/NROYe0FTp8HSxKNIbOszUaE7UrebrgXeWXRcPTa3GP93anm7VQiKsS8xEhj
gTGTNvcizE9jONRGYD6+h1H6edi+s4ani+fOID7UkEvaBOG1Q7I56v5vK9nfiG7Iefx2hJ6oaxGC
0iXKgH8AF5+mUh6vUPEnp2jUwCExXtqtGfmFo8FFK2YnZa8Vi7ek+8kg0W3Cj0QGfOKblzPaPens
U0xmtCJhimjXu4K7aMNxh0PBAPTRRoPRMSfCWUNUyYKKhq0nDJnSmHR2aYVYtRvPa9tpFFeTca81
EWZ9KZ7YD86+WX7vMQV1ntcxUNxejlReVhZmV8HPj7t32+7f3YjFLZshrgQHLdko7/u6A7C9WBda
XQg2FkdAHbBa4ndoAQURIIRLBdp4b/ulDlAJHJIMfWKCXZM5DWq8B9HuYH+jrFviU9w8S3ZczYjl
eCT7AVx37E/uCTSQ6iC4cYavdk19W9NVsYlVqPA5FPvJFzGC/t/OWbvXik9tFm1/Vq+ZkR9ehVv7
QuDmDQcVwLv6hrQ4Zn02gLuR+3T3gR3pMxUf72SrAIcwjaBY/1VnAJLD6sA6/XOMGNVYyGDtjEb1
rApePoxKvlsFVIrEOFpGtD+wLZJjsvncucc/qO9FvDpDcf4tq2jj184qflRJdzpWH2bCXsJlxVix
et46K7U5tht/wVEpAtsl2BGLDjyCQkvBigr7epAa1+FVQT24q5slEk0mc7/GCTTFMy74X5mtkRQx
T9/SijMDxdK9r/DmpjSnYw1m13rlO2TSKmrtp//LPz+TfKDmd0JMgD5W8MMyyCmiMtL8GcXWYS1d
zQQpqVknkIvY60ZWoQm7zKt5VnaYWgmLi+nltEP1B9zyRugd3TnJlm7ZjYBALZM52fVtvnRwNT/T
MGMDGJTtYtLGYA45pe/9F4tXFZcQVxwTne7T1JbQYZFtmYWwsOuVK/YpgiDWBGn8IiDEDTN2nG+F
BxB4hZBskICPlcJmRj27vK+6M16T+SLviJkxJtz52uPshsMLn3UIRRsyhbNfsf88Bef4PBr8cXuv
6K6/0/EIpVcnenlVdfWtEUajclIj6BhR86ly3fpck8n6eLDElcqm8QGf2SiepPqeZqzyWejLUfGC
8lRZLlHHZpJQAFz83xh3qOHRrPDSkSc6gD+fPxmSvZvMJmPOl1RXxkbT/JkPVuWvCekXMq2/bEo6
HkdAcgzudF/+zthSjNtZlujo90+yoQ1svRHYuHF8tqPRBfAb4aEqMOe5qeitjCPbsH9Of5vNJGUz
NXMWuuILiZzBndQ6NWyAh60dNd84wO5lCESO7M/Hsn7niSGTks+X58SRtu2SVgmMuQ80KImScFuJ
B4ql81T0jb0+5BzxHmd+nhLL/Dz+/6Mn9/LIDV5cjaVqpXIp/qrnDCyI/ZZqtYzHoTXjU41X0uAt
DWSc0ZIHOeSEui3mNfQO6kLCm1wYnAklwc2xZWE6nT73+qmZGtDlQXWGoqFRi7xiw135TbCzK7Iu
F4+5jSYoG0v5mFpm8hK82ij5zFQ/mCm5XeDyPpTqez0gtOlEvSkkfsKQf3qQwRJcfGo7sUAU97So
Ps0Ad0NgSZ6wcs2esJUN4ZyQHuTVfg21LlXoo7bZ+dRfKGY1fO2AComorcED3cDrKFiu1vteG7pn
9aghGTW8NCvpkjhCdTEbaZsoKgM8Spr9QF/TmEf/yoYNn7hX9uxYdoFj5gDuMC0stWYMkAqnx9sU
ebGQNsoH6SwqCLwcZUW/g8y6mgq5hO8VjHhUm1YBiXlr5BAfPfX1Aqz2wpSB1Zh4YaOyhokAOnJm
4UiXlvUHHo9r+pAKnbyu5sVGnlvTyWzkOyFOYi19qg0wKtAxKqvXnNEsfqXUUNkbDTdZQPEB2G0E
iKrgFRdRRcxcebb4a6368PkxdpJm3+trL5tzYFlQv8huqaibeRMALuRv7V7Z3sEIn1zvZ4vii+WM
J+feqv5Jc0WNE3MxsYc18T7Kq2M1Zq07CZ27XLvJMIoXOlsVdfWnFW7pR3CfgUdKUkgWxTcVsG4R
klND7n+8PbuyeUsnQJTDDvhjjjsCKq3nt0odoZm8eq1jvhXfz+nMKUznoY/VDBvRjNFXap8Zybr3
lc0ZdD7cWkm/rbbD6F8rqyZZUHMOLI48xS6PgRkue/OOAQEQEsfcx2Twpk/FvTnh5hKZgtD3w6ah
g9i07T3JD39uBlCp3sFgc/65SDeEUeigsGXFrbdVaZ+rJSs1uz3gy7bN7SXa+0jRJx4pHFrVfLcK
SFot2//1xtC/4gPM+Nu+AW2prYtArqNb50cnzXvteQ1lcncfao5t9Jtdej3g/sxm834xqZdNNPcN
L2dBzReCcBRRsNG3OiJnhIsDsTPiO0bALZBt883/MXr5W3TWdP2Ngjx+DqcpBMPBSnAQGGFPguIc
qoYosVJwL6uZz3tRYy8QZXvk7sFfxNyfaOlz0x5jFzAGUfjjRwzY/LDn1oNQlgy2lCInb0y9nXtB
omzZASjKK2mdbfqXYFKbLlG1Yk79SDWQd+eHaBO2ygDxJtx6y8FaeXWRX4Qk2EL3VxwtpEKQ/Jo1
h4ca0IrAMXtozO/xmdI3M6GU8R0Z1VtaNFQ8Mh10Z1OFXW55mtB7WPyCPWtrKh9H06zlMlo9VVg+
NGpSEq1fuzEdciFbqz5ArOGIBDBoCCkC0LTx6A/nNVVjGCDk4NijaVFFn4qcZoa1vRgqodFnuF5q
apPpUJrSVUIaIkLeYD09Yp14ldmRnV6GPWr9czhy/ziyoweUpY3uAZuQfR5QgWgEQ5A3qDXl25k/
km40rDdIytf20zqoujKUw/2vc/kKlPciu+JFZNx++6Bm1ai35rDEGyqSXq0PRx1fMt+cyB6zgVDx
tF54ypOtwqMZ+9dtKGvxXKmFShGWAsNBjWfEtqmlfvms2QnOv01YsIWihwVqNmOqfb8aKL+VUI4p
QlQTmz6okpYD4mV2ZY4HgeSFZUu7syAyl5o6nbVTs1DEvxfu+CqY3/cFKFp2ZE5yQ2jGvpfAB+gp
2GIZMjNSTDAX/+up9UiSFP09goRfQL29ziDvWoPeWn8JuU0X9rmHcWPyD6/rNhA6hIJhER6jspk/
evEfFI/k3aOTTWg4h1F5uWjkLSErRREpqNm1imatXUF0Rph8sqZp2UFVIwZXk3KL1Mw3MXdLxJpE
NxIx6wglxgEi2Scdtt8AgIdq8urfBXV1/MF2DIosjdUfeMlxekFk5xnyRmwxl1yg/HYpTWgburjz
EIOu69CA1DNsf8n2fxYD4+yn+FobLNbj5ExzvYpKo0uG9xEcGI/aiuexbDzY9A1o82pXTUUbOZen
8cbNT94m4uy0aO3vWr+TEyZYDV7Kk+d0CWJHIJPP1zNsoR3GEfHG6K7MVL/a3xba9WThLTsg0QMR
uc3SIKWPwKLdLd49Uvc9isEmTKNTbve+ABPZNvgAgg9hAImvKSR29wt1sGCU3/cigXU8hb16hMdK
yASCC2caAixTl0ZMjl1lXVHzuJA6TaLgSvvai8Z7s9wwA9/F7hcYsMtim8fPWII9J1djQsA/uQJS
/yk6KyifNYN4WHPbi5Yf34CWW4GWLIyVJdZT5NZ8r8JatHo3APj9hTI2QTkmpXu0ercxOaUxxmKg
C7FHL5aWsFg4AvA2EfpjELckg8topY5hQUKQJlLw0SqjjnXr+YI/Qe7ZwWRLVUN9jMWmk4jJjAPv
DUGL0eyz8D4Qs0Zi4pbdPJZWtzTrG+50oVFGI5biVfRqeiPoOByPy9G+1JubQmuwmAWh/fgWZhw6
XpQf6Y6lkmZDj30xzhK0V8hj5Q1vtyIXiD0XG6fHdCFxzzyUI/a70W6Q7TnQeAvLtvndJTcrauOK
ZUvMMPP5xlAiNC81DbxxUgO+DKmF+UO6R3MMBJuNEVaf6CwUWA2IVSYgssgTsOplZ3+mzI8Dux7D
yp4HKlIgY1xW3wUiAO67Ae5t5khgWcwSLVpu/zf6TSnpH2rpXrfOJNc6e16Ho3+4ZDwzfSrPcgbp
+qWJwfLHo8uHdDP2ioPoPFBXq2KqbCQxQw5DlQlW5bqLwiiTPSzpHsEhjMU6XiKuZEJz6UERJlNR
lczSggeBcQlJcL50qfe5ahi/y2YB914nA4Gu9KkiRhwkoSIAkp4AvlzosnQCipHDQcqn5fe/vrhs
0c81m0Ks2TN7Il92yD58uSEWMwmM7wK55qzi3vcwOlNgEWy3ggQoehMNPCrt9Rd7dpIRsDMIZqt0
+Q7P46yH+5rpTjqgzAKAt2Hrq2mzDACDVnuL32bKntF5j0kLQ+0wpDJnuvJCip8d9AoZCyj5DAYb
u9mdkZs1kAFUEUSEVWv1tnOX6vjwCSB+87soLNB+ugLZpInimnZHbkrhKmAz8uJI+2BNRteEulyZ
DN9YaurbIOE+kWVqAnk+fihOvBwYgGcpaHolXqvsgW9xYk0vJJjnge+hF1ZBRwNa9XcfR5YVZUYh
VIB5TFqlsJnqGt1gyp6C5IJL5B8rp8vwxmFFGQBn1Nq2/01MHD6nXzqQLO20EfLuySd33DUbG/y/
AqSvGbAkfwrgXndHgcFGvgkBViH+lcp/vZn+/pYB4IWYEMRFKqfojcS0uoZhOpCLzfAjKjcPd7ia
gy8mClgOjx7pdP43QIJ29MNabIJGj+J9IdBc9SPujRpdX4qb71nCTEaWcitl6zW2NmKWlN6o818i
MEnItNteUhscIuUhXXc84ka8BFEKa/7nZ33uv88tnTh78Pm5n8lXeVlGwKmIHVevWcvKoPkWkPdc
UBqN8Su/xcyMszdNnBZWPU2qIrFpBb/bEgP7WgB7Ek4wN+/PbR7Thynor3IGe59j5BxFew71pzKj
7Ostwac4zNoD13vrLESdcWCHv2eSgQoElUMwP9/8Vi3F4W8rlyI7NF6N6PLZm6uzGjrQMZFKLSz7
fw9KTP8DyBvAfepR1tbwfzSGitna3EDI8ur0MxIzPU9ey52zUElAVzhNXPkHxVtEErtWjySKKyFO
eCdCn4eYC54KYMd63TV51e1N4R7U3VkvhL3jWgqRcRQ3+EMLLX9lAdqWnPY4DrAiAS3l2fUahvOT
L2hGvox1wMwpwo4lr+cQXSDsdTPQ4gJl4vDtzvwxo9NCjKprdw/IrOoiVfgkp8zCFJtYC1gbuLL3
44hvZe4x5daMo3WC2hnr3X0zzk9cOZNbBuWxVqBWW9xYX6HvFtlF7En2/Xpk+mz2fLAQiJ/QEj/P
oQ2n+e4f1pnGCMeO2NI2jvGyPKWcKgkATirl3IOlAOZkaBNt0XhSzhlw1mmtoqP1zW9JICn7z/jb
MQOdEEij2TB9kCruIQhC4iZkzpOshVhWEIymxHRuKyDcti4vmHrDTvDsbuNwNPDmesq/EEaR3d2I
0T2DvxvhO2twGUkoERQmVA57ocPCauEZYABzf3JDWlSkh5cM+7zXHjpFhvMxieEezR3rLDyxZtmw
Nd0hpwAOZ+uWClg87NSE14cnxVUeDGtNjSwNjTSvJuCMMwpCj0xPNPlCzzuArOyBalUJKZrZCksg
idXazA/7CLMH9sAfTOExcz0RHecNHSeCsJ5bGxxmg3jnAgLNIVZkDAB/oiyk41mm+NYOQsK+D4mn
yvxLheIEngRIRKVaRChWk36yMujGQj/wqyvZOIC2hlFBFFiiHkeAyTuYztkIABLRSpDJghCNWkzz
fKH8sPZfV+kvMEf5caf78gu+6HTNWCXQpr1F07Geiamx0YNwgW+6eZ7KnrMpU15QHH4ML2a8YMAL
oz2Kh4m317l9oKPVN0vJJtgE7h0WzGvKhU++NGKaRiV50K8Ew3Fj8HzRZxwYc/azTjeNIlXAaHWm
cKbzjUdvc8DRSCpOukfp9RYZWdgVkZr3Cz7FCHVdnAieUPMFE5poIWGBLpGAgQa7j7XIkC/cb12g
8qjH0RZNI2VbSPCz0ls8LaHAloq2OvQyU+oV2HaZtBUTJ3JAY9+WnWNrK1SmE0zrssWYGqSSPE3v
mVa3ER01j0BLnyTEaVzv+XG/Dj+c2CMrVrLIgUtjtUMWtFY4jCxlTCZFLIPFdCGzj+aCmu57Pn4S
LyDH97G32IX7ccMebf1UP4uO4xtgkoaHqJRUX17mDYqH2EQQ7yqTPuuVU/Peu+EKYTuFEqBnZmnh
8+o8Tg8IvmLOxCUmYL7SjvtuWA2Mo2/zUx1uPcYto9NYhhs6HSQWrYZ8Vt9bTExe+6SFqC8nvBON
pLDObtiErT+6sKFwFDKOnpcumBuvMDWzaHcDWuAD/nYb6Tzdz/0++d7QjmQHdY9kVSEDS9RztlsK
Yf1tJFY10Wi74dU1e9iyb2c5M4BRZc83Q2U9stPq72kE9Dr9PGs4Lo3EHcRnJG9sgf/ACfIu2wfn
p2q83RkmH0YloTyxcJD1lR7t2ySUe8InoWZva1VgQt6FZ5Yi8BwAfTBJ1ssoeAD6n2ojx6+Fxzou
iV0aeT2hMiCqcH/2gGz9jYjoLeFx5kdru18BEOfY2FB7YMce4YYYsUfEDANSKu8mvo9g3kkSvV2P
2UndqqNphHvLE4TsG9vZeCVdiJo3oIeu3gMqbqLytPjmyqTziw+eVL1lI6PEOXpn17Gzqy4rZa1/
xG3GZ52gpjAUX/zcxx8AbQyQliUE+J+Th05gS5GWLUba2bmZJaBLEkMHSJvlokktyazbMcC4TTpb
KX8lRDycFk39JxloEX4udwNTQm3JRVayG5e9EzJ3N7AXIX/gHVRqwKvdNYrTMpt/vokGXLN+tcoy
L5QrQsB9VLWlM4id9IbXOwyR8L4tZFFXLAGhIX0teDnTpB4AblY5F2zKA4gohEyHSy+1y1PLFerM
SVcGU9lRiJBUdsIpUeEX2JS7VFaCui9hzrIOhffLdDNS8gY/zu6ko2ggHIleZFSbHdMW9/NG229d
e0vxIBkMBjaxhQ3B/OwMinbHPOeu0GLI7GxGuhVqBI0lVCf4cpbeVGfGyXeB6O4pCZlbe5QVG4g1
0BLFrg0kBZJgX7spqVzKKHipCFbb55pQO/JjKaLBNEBswphPC2wLxryAto66JpuAmHTn2X+Xnkz8
1wDC30uDbEkbCKSojCfAwihNgQHlTuW1eNhmjK9LS3Fs3DrSodYogESgKkIDNewHs5yAkfyzODy3
UxtgQkWiWdK7yG6rV3S1fV9Ft8u6JFwqP8S8Mm1RkCKKoyeyFKb4y3NQutlHXQ5uaVTOTN7qCuTK
6jxuaqsIwei9cpXwRiHOp8xVJuGUVLPyWDFDjhh/y7lkoymB7SuDu8UzHZt56p4Q9Mu18w1oaptF
v6pZVBceKJqxXQBBtjRX5F2GMdXerrFq4hAksHnnH8Azg3lgxv7MsCbCWXvtmq7lteWVciJ9fPMv
5j8VcJ6PcDu/VAhmY6Jrm7nnrgrBysrWeudCOrp83qIJmKAWfK2Bl6RhLyw1E2PCAZnETcV9bNkh
q8y5WFvhjUYDfRXowYMmq7agp1phHLMH4YnvTWlIkxjBmevu3AfEiSeV1urR9RJIJAY5dgHxllvF
v7r+aMcawka2Bnq6ghNI3vVxyHSShS8RoXVQ9pW4vt+rLC6muZFnIG+fh6+IEPW/25aOMkYh+aCw
jvq+p1a6L1j4H13ow/98wqW3P9pWlmFd+jX91sUKsrQW7a9vZMKz7UsuwCeagglfmUj2CC7HklpR
06J3i7JTZG/iQnXOZMT7zYqZIoRcC41+NfR0kwhdg7R7RxaWdJ0xw39G0YJs050Fcmle8eI4vrNc
DRFaURpSJDUEe1rqfZ4tPYHzH7I/+YT/sI5ThZqyQDGF+yZowE0tvp43cXBEYlv7+h6CvM1acvXX
Xz/qsdhAhU3GCBtNjlsTyt41gwed+13HhC75ORNBBkcRLO2u4kmLyGv4VCXFOwHEHSddkwibMIy+
+bMkJePelIpTLU4hqIF66iT0Z5HTfSpqLvlHDBgo4fWNJTqttOTEZxUv5bm8ixPV06gzo3dOIF1g
l9mR8d+IU4LCuqbm155pW5KBpiPXxNXL0mik+a2Zm7e3ZJ/DpQx5BCLrNYTSHIWvSqNtj78SknbM
fJuNaV4jwKM39GvBmTqbZAEQWY+hOTqmjxx8rEWDlgBSa33wKqTFAeGbm1eqKk9oN91tLCJ0yjRB
vrgIBmDcQGUnIwrnDZQ34SF5qkwPhavCwrZsVZkOMa0VtqxaLIfpJCOK/KAK+Kx452A4ZsZwKCcs
mhRATcj0BKYsBIDssW2c9pHUertgUTyp+ttlSLemNrl6MZpuDIT08xSnZ6qIGgEo5zWwWd2BCzjV
6jLwHQ8XKTzPiTij4cq1FTS+RWvaW5kDHzBopr+NTD44t504QBZZc2Xsit2Kw6CY4D7q/E7kW4tG
ieQOmt7qtJvVo2cc4yI0JqRcJWzoTahvfauTGUSo1f5Uozu/t9P0oIbdEV2MoZLiZkvQA1XaQ6zw
iPmbNT+ieZI+xO0TqeMdDLJ52srt/p6uL9ug3m9+DPYocTdTu3KWNuqo3nXranNfuDSLGzAvjY/4
JD1uXZCilVXJ4mN5tLbo+C56IaF4RXPaMiBP+U8WWb7mw8YXc+OEolygRa2ICvpWwGyof6SD5Vdm
mvCD1WbUL9n9DF9z2yMfwGaYYiMgxnXB6jfqUvRebRGAezO+E6W/BdkhaQKEmokFs6aAP0g1TO+s
8BNWmo6Phlfjhpw0+CN0UoiKUphQTUHU8TRyIxj8djutxMitLNmUBElGgGpCiROrJj4Jt+jZL9bz
+tDeROtjnIc57qXvcNRoI3c8LKxKcLDcTN7FRZhWYJW28kGCYZ5J34EsptFkbcR4bDOaIoipZrWt
1Bb/hhgdsEaBcURE81/bpjFwpxu/0lEbBfeEeHkwK+63Cj6W1JwIDPjsdjJF44bud4SqdZuk1e1i
zSWwiJ5b2HRhorLoKkVUNonh6/bWlnZro6zchVNd98lhjJ5uGKrAy/eEoDLGc69F4YHXv4X/vCp3
6OM+Nd3xDLPgi+g684GEdGkfwE+Zx1buUwAB4WikqCvUZKPootrm7Q4apjvvnTphQ3ZAenNcc6Gk
pNMFWpvQ25OG+/Wui5QNn3QhVRvcFahFecveCIK/IjvKfzVONHSWxWD8tHaLPrbwj67QGve6zf+d
VxdOgD0L3yzVznccRlOo7lMEn3J3q0w0SlpQi1zSZkZkJkJ7fAuqpOC5s7fKdU0qmMoME86n+gfY
pSepTVuXwMZCQy4PmV4D54J0xgCi8wSadq2Iy84RY5l1IFfwZPxOj4nZy/DhTqG0McDZUZjWREJ0
vtClTVw5XbHlDRfgoe3pPhl6vFvGLwOuPQJz6VME6ZhE1rR271UJqzqhHmxT48N/k+poS0Cpb5JG
YndDh3SVLu8A9gceMoiT7TQhzTzST6UfrLWYQBxJUghAD/VLADN4Ns+bz93nME3VkElvIaz2/QNU
cpFalQwiTe6oqzeGKzB41oSa2iu5Or16dcw+04oW4IAl0pK4vKLsW7F6m7RBQwUi3Gx7LkU6QMKk
o14yTmSgV8ujPUNu5uYTJtYK63EzvLQdlBUbwtEX1Wz+W6CgeJ7S3chiz0pR+ZkCGHSdNo6ECZ3W
Xsd+f7z5ae0N/5IcUYbI75Dj9cSS314xddJBcbBlwdK58jVfdA5Oa3TcqQUUWvRv2gthbedz/ZP8
4PPxeZ/yNXWTj8PWEqecTi+kbGEYZaHjT80CfHVNkM4tLG8qH6pFmvE2zL2iVzZHFWEWEhjfss4E
GA7i8fbrvCLunyMFewzOXIMdCWNoG8S/VQK3WoEGdvCUeAqERd/CHtTXd2HcQkjEWL+3c2f3bI2k
iob5PGYKR4yt4ksYiGnyMKeGdGHqJV3dopdPHbqeq+pvoyDA91z5YxfmhO4ZWZs2buAFMaDgkH4d
S+xETjlmVrcw2ZFLn8YPtbXAz5oBv1SpQzeWgHaJNfVpWSeyOa9z/8LBio2OPQxoI/KiU4kvV0Sn
VU8kA1qgoxVpv0M/fIHUDPi+QG9m4KXm0xjL0hSvmo3imL2pFa6yAXnFG0yN6JD28K/POrl2PI9p
+mHtiSidAx6l9CdAn9gdDcvLr1oi+1Imo8WE0WXoQv6gmE4uxmZS3l6XUEepjqDPqPSwi+NbizaY
pejzTXFrPJ2JVc7qFFTSQlG5s40Uvbu+8K+XvZ5ajHhFIWSH+3IE/tigZne4OgdIu2tQ7LbB7pAr
Hvv88fPKOkBbRSiJ9hC8EFgvSipESWsQPgvMuBjjtf/kxqldk4fbaoLqLbKN8dTK4NW3rAwisEdr
ZSI5vJsEkB5JbzMTFtod11UnR2PWDXZpUoMLUB4iNjoC0RrY854G3RNWeEaFP6MwYl6H2n5rYM1w
Ag59mVwII2IABqVY6Y1LJaochuo2RIXO5Kq5J70rcAMuWGMz3gWYY4N6tgb6MrUF+pfiK1g71btK
KKadU1z/FXQJN07gdRzXPjAo4WlWaobAwexjZxmqrWF4r/8rJ6eWs5nC37+GoQvA/VbZejn3s3qL
xW10EX1xMGIvz6r8jAmtzigL/1ZnJ+XwyqmmcwHUMeDNE786PC2UrC5yLD2YJ0fzBO9pwZtRGy0g
CYQM2BoITh6d09i2fsT9+UhZ/tJIytFXgoBI1Q8YVJKJxZ47GI2YE2i7EqMiFa5g1O0LSMN1D5qM
Ytlc8c6Uzs7MN/VWNWAIpVt4HEOvu61ibBsCdS8aKG++PU3NWieCeedyQPcq1heMcD0ljrJj
`pragma protect end_protected
