// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
bTRtnpWmav1lsfUX/zT958O+RUOlqG5eViX9NI6rrH1beyl45pL8JHyGSW33JyuE
m4DGb9ZCeYHt3Xs26jALWkxGh4poOpRgDq1+CegZrfYdrKl3Mt1AJ5x3fektRFaK
XmubezWReqMzuaNz101bAHwpuVG5sxSlYZEabUUgRU8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5920 )
`pragma protect data_block
ztjZBTP+40t15XtWD0EIFPVKwwwPqoGuAF21LLwe7RWGLd5gSLRejgk+n/BfMJPS
4yw93EyuyPpJ6hBc0z2aKUhovNYO+PENyEdlwbggcGZmuEBhZzgrwxvJW1eqOceF
EuUTJvvWh8LZCzK0lpCp90rGBVwcIN+nxSDv72EP/DeW+DBg6SgLu7t1VYeAldBU
AH1ATMgDBzORcqY/72EzyNnBEmaWWZqlorci22VTZemL9eB7G3WxA1S8q5NLpLS/
SDcyjSl7clWs/rb24QZdjokCVBSQZ/kiBhHEZqAP1bRkBrYsMldtzCCHrBKvkPfw
B9o/x4lBH/4JclzyLLRM2z/RVUJ8fCpAaZekfGo82ZhcGevGz5AfVnQq+99ZTtrn
lJqXr/HZ3TuOrenECy3Yp5mxwJ4MWEmvYQ2uZTGDK0q03lN47axE+45JhF+fMgfM
1NBNpkENolEqluj+eHxGCM1keljyQtHuPWjObDJIJu7wuJ7mXC+04aFg6GwpD+mL
u51ifVmth6pJj/b6UVgpA+mljCTqXL9Ri9t3ekKA/62XZCpXGDkGwR/3X0F26Cl0
d0DerkzRdo+bGGHRSL42/gRHCC4i+kCF41Y6PwaGKU3MoeiBYNXmhrzum88LLloM
cz6/ymheMgx27w8rNf8dQsJCWfXYqYdCi1NrDxEJZH/KrbGmlV+csNHz427qdcyQ
8Cf2TnVm/3E9DcDhomMqeBbVfXGaHzxmqrO/5PY8NtuFqCala/UVaiXQY3Vzd87r
7ru9MoFX7smgZb9ouA9SqARxcfYChLWyo9CcRVuc2qOxsjINZpLf2LzlpMhHZrsQ
N0rPf1lb99p+A17J8vYMK5uFXJLobu2bZikJUpJV2C3VYks/sPYwRNZH5pdw1sVc
2WfbnmIOnxcpP5AGXEb34Cx5gGUS4vB9rHqr0PM3MQ605is8JNHGjtPe/YYXrXIy
tsSKj7ctZUUaVvVm21ql0GAppppWt79BU8AZUy+Ltun9vdILPOWhXzBIBVuA/uQ0
8901Fl1YxEyHdQPI3NY54GiJGeNi1CCJOu/eRH5Ai7CeMozV7EUzTA9X+A15hT6+
wRVmlX/BJ9q8WxPTVyIubShZH6Aiey+uloxp80t7oEnjGGSMTKwUZ5W62RUZuc2o
/BjWOhNao+sgD13zOqitz/dsTNucW6+eILP9wKOeQ8oIsxXtzBBypImKq6/BxRhu
8pHg1ZB46Uy3qvE9gXyC2t1cuBDke4Zm69GEQ5yOlcWJqB7RiLI3d8EwdmySL3oe
mmYoPhbKpWlEdBwYtJ8pkYVQ7he6Yz6PojmBjxP8uxBq3HvoWF6nMkZxHIc3fuIc
15jp2knqfwjVQ6BWKeMUa8fCEzT9k4i/VsU9Or0Xd3CgOJufKeIrw5e9EKK805hW
hvojanhMCzQE+24Me+G0X79eGDL6gAl2FWFZrarhHnuGYZOTWnx3R+6H4iXZocK+
Qq6RYuPZGVCJNdR8Se+5YaB4yVfREgA4atEP+V8Xl5Ojh4VqgP3sXG9GJ3azSQ8M
VlE7hXsOFkAGd/dBzP4MmGzUMV8tUh8dLTIcJv4euZp5luNLGTx1jkXEJxdINgo4
8rRp0jDr5N/d8V5WvclJpxlUfEjT/rCAglJL374HaMYSoemNK1r0qfKBW4GapG6/
D3nbsGI9BnnLK6j8PONrJp+kWPbkUJR9ZOA5x+CBgU7GgGxk0QFnwCeLc7oJRLqs
s9hf/0RkXdvSCK7VpR+SOqrVY88lWaYfCsVfrpLuKpNxHO6UbIW0pTeHX/g6Ap06
WOy60g9wdjvEWRUDgQY1OkwQZMoS+4M+bnu2HiYpoQRLAM8uiF7mfYonXPXF6J7A
n1MuDGYynuQoPfeybt2fseUYVioUvHkLrwM/XWZz7cyKRyUWxU+7I0zUA0vEQKj2
4KLY9+vwZcQNt8j3yNJiB7ij82bUuUl7K9vkFaLs7aMvhgD4eW0OL3CgVThyETPh
MnChwoxJOK60SQm4bViOxUzs7iHavTRTc4hi9tu40w+/pX3jdY9Dj8AYWbIUOu5V
STj7DHmTqvRpw5z7M+ezer0c2mLh0lqQa/IYqVWWgb2Ud/Szooj9L5/SLi92mBAq
lOmk1AT4iW7f02X3UfQA40n0XVpdEe24RFI/bt+/aa+O5f9Ur3KeP+OZ0ZWt2c90
jVdr3ZZuS0txGKJn6djKzXgJsuB7ZgNXHinPNvIut3dxidiyz4J4AKuBI8Zvyo/7
PneGgKdxw6xosYnhWrTEZDVQ7l20UzZ1UgXZptevAxFw1YMNhppPJwD4AlrEtoDw
0x+zot/6CszcZbpQwMFq9sm7O2DzdA7NgviQqpz+rVF5RDWVmB1Wde5C52t9BbvQ
Nbc49CTJISPpKwcz8wOWg1Kr3hP7HvVmBI/x51QscEt4Tg1PUvTwInHYmsS9Qmib
jLsLtQeX8VOM7GdYcNdsIGYjUUPtiFrD1c+cLIBdcW0qqTcS9qDYJifs0gkJsAPs
3/32QUYfzu7X17odei5oIhZbD5RiP3zwCRYD8uT8aSDMw8HaULSCTLQbmdGWO9es
9Bu4tU8P8H/J+ntVOsKUwzU+QYp1pzFc94h8XFjTCdd4+r7aliRykurpvuV9LJMK
cEKCRLmz0T/l30T0p4TimF2rf/UhFijyFbTLYvYhoBkgvW+JHIFDldBLu+6izd6m
8Q0kj/c0YkQci/6lGmJ+gegXo+mS+fPxNi+uSgOaHu1UnGXH3ryiDXOMZ5FLfBUE
zBNH6v3i76qQbXakf5Z96K1aRYm4JnmbSUwg1h8gVtUZu2hdqYiiEGw4BMmc/aYo
aLoghdFMfmuDnBwZShSoOySwAogDfIwypJw0MZKOuJcTdFMBid3GUlJw10zBKJTP
EUpbOpaWCE4KV8wE27daYZMs/r6kNSsLLbvypiXZ5SCi3grthamVn0nvgH+3l1QQ
U7tm5dmhydWOLBiKo7ffBvIgDW9JbOBSSXwSiN/uN1jO8rMWL6+v3nj7oypFyf2f
oBvP8Rma0SDWENNFXGnoIknHNcv8nQvOBASMGClfJffz9ZCNfp2r6xZ55mPoVXps
JjSb0l/hyvCgKsyYrvj5AgpH8nOk9qhcMtCTTrflV/RPAArzEemX/JI5VQQV0zRJ
csY8BzT7q74cyhgnGOF+0psjSzdxcaaUjI8KVyV2N2kkj/TyeF4poqFyDzvf6jFL
OFcM5yHW69Qjcac4N5W0uskvC+nAwELWTg6S0eous1uBNZ+wcI+S04klDlXKwiZc
rfuaF5im3ECnP0fCRwRJbXGMTgWtiOwb5JnUFkn9ZXq0o01vIoQ80QptWFtj4Gvy
mP2ACGHOZLecVXWtQbd1Mb2l94NSn2o/LL/2ihf3sGRkBK/xQ730MJUMQGvrW+Ry
kPsPrLhwpRdWna1GKIeUvGkek5rOWZpFoynUuXv1dVZDmbQh9bzD+cJKKiNOPgLD
zAusYXtbjyU9N8oJOr1+dQiCjp1EXK+twlwadVhG2Ou0BpHo63ttXaLO9Wbb0y2X
w7+FMd931O193cRdNUEl85Dw3RbjoUNpy1Jc3FV99tfgk/XLuW+PvkqxYPIMR8lL
WsMF8J3FxV+f1S2RI6BFdedxXVC705NRLX/TRwl3tYiXmf7ArdPt2zqlUDsnKgI7
ej7zxadCHzJAvEhisbdvm+rh8EB/1N5/iBfLYRXHiFLxKl8JBc0rruYdiS+8OYet
hDZiYJrD1OXJNF8XQq9GpKM2T4KGEKWp/jIIrGG9Wy7yrF4NTDXDtfDfl1H1bkJS
NgS7Gyrg6QJSZBczpyBakJbQtzSkj9Jd3z5aN8RhRrdrPIL/PEnAVuG7VNiPSO1g
dskFEVHqdw2od81Xg/KWBOSApHRwigtto+efu8S908x3rNNZrvSNMUy0FZ9z9FPx
L7EmwMiy73PyP7mz6v2rKvKvp+/AtSZCOtGMtFb5FLp8QQp8eUkftlBW4D4yI5/K
N/ol593T96T8aNRNwkRMcGiv9ZPum2J3z7C1cJJ4pvYbD2qu5dVPokIj/8iQQsTL
df7NneQBQKi6rjOtVGaIhcSp9aAhGkS6BlLCXZrHUhK2lAT+3Ogc462E2FyJu5Mi
e5yiJL+M1hTDXffy214JHlKoBYKM8HuB8vXfgt2BHXZAHUF9tAoyeMn/8ESEEiLN
wULBLMdfFThaJmXjdihJDm8ZkXPrSEJRXu1gZtZ0eP5K8Apvle4FiB3T1Xu+Lceg
sGxMNhJWssWkc4WcZXpRWNBkP9OdSDXU8NRbJ88SRSue0fi3Vuz6UhhXmsvHP0i6
nppwJoupUzuxC5FbIu/VKMtBhjUANBZXDbzEAioxGl7/VakIPDqJjOXoeO8wcTV/
KzFbfIHummJ+jXSEYmYBoT8wDZXrvTOg7WxQUP+1j2cWP+27X3Ccn88KH+dP59SZ
yKMZkyyvcj0R0sj/I2Dy9TrZ5ZBlC+ld0gwoV3vTqg7V8BKq+KeVsd/8+E2FcsJ0
mfy0QtbvxA2ZWxbepKn+b5B21NTOOg3r+jvdarWgaNQeakIx3Kd+DGlDBFUU+1PP
U/EsM2ZDjdj4KoEtOHgPO6o8aQaCJnL66AC3BqbkZxTcwmKB7mv7avPw4hrQj32k
QkFquLCAQL1B2IeLxv/pcl6ntaIOLGD7XxdW6xOfWQjfZ3hae2cv/VQXGxGakYou
3Ou5v1xgCJhEhN6j9SAYAZfABDMp5KSSbZLZBJ+Ej0XRZCTRnfyR8kWDAstKLLph
okAi6dDVEnQA5jqffeylMldbpRE3bnV/9q8ekOS00E3HxtcrNfpuhWyJeqjPIuZm
FlIGzjsY4ZWKvnzp/2D2XWttW6N3XiXYhk4MIGAzw3m3aKUwgxWPqgPs4wgQcjyy
x80GMaYzvD5cafSnbk+kGTm9oWV7z+W5fEQkERS1lCChBnrPeJvUW15hIUcKRI13
RDi3u+JyDi6OsQ9Du0aLvV8j6xchWxsqkCXjFW1sQhg5RqUFY7UT/xYFquRLM5sC
/0JhrzVZM7MOU1n3SeSolIafAfukMpIFffz6phBnJrAoOS46kPY4Nsp6jwN9qkr0
0tQ3Uy97nxkj9Yfomzn/YdL5ZI7c8erk3tbkllRrN5BqmMq4tj2aYSp4hP/1m8Wl
Mq/E4RZjnzDEb/IejkiUWA05YNdGjWliNTpgaoDb6hOJYvZ9Yub69naJ5XFNqS0i
v4ZvwoWSotKrkXzothN3BiNlDTlOeGuuXZKXdbBrhWiOmcfd8bvFeiJHcoIgsz7B
Vbe0NC+VTnqb3BgwydiNlhAdKIIsLxVB+WHz5b0A3Qww1d7jK8lYESqr+fSJ9gKV
/Ls9Sa71G7J64kXge8PNU8es4qt+Y11kJ2Kv7yKQ7aeiWTmEqpEs5tEaTvb3Wx+d
o9Mnc8ce3zk79SXuqsdhABhrHy+oleAr1b6azU2Y4iKaKYjTccI7O11TG35hmX5D
+BfpP/ac/0Qpe5UKhcJxEQo60U9FQWZAEtxJoGJEoc4+KtjnI563WYpCcc21f+Rt
7V7z3V7I+CpXoYjtomE0m0N5qF9N3z1/kZ7xxG8AUDIsfHLQafeCnLazYQzUhnl2
18Cg4qjNM7dNTHfb7D5HFPPrlA7UUU4DE65nrQejxRRUFES6Y7etqcJAoxFmApnH
WUew+BiCV7W/noQ1zRGpynf43tDj3GFgOztcpk9Yw7Nt0GVvDgssg38WfVzWOlkg
6IY1vDEd2xzoV6EjX1dF8xkyQkJ4RkOeKfWDOi0EDihu08skI1s2LQiMwkoPFhZY
eP7na1HnynalYW0GBjTfh0USyMjYOtdjgGAhdkxkQO+p/1BkjS0tWWNtci8pOsiD
vAl4ECAiwSVNHsqwvLIIZ7eXDKXb5KluGEYCGn1E8oumj71eyw5qauBfZUKCXgGU
nnQdclJAwnGnesbRvLYD6rlbOtkCB35rh7eEAhIYiaJ37tSCbFCVusw1xAYEVpwX
Bmw3wsMs5DEsS6esy5NRjSdqO0LJCwPEI49Dx3NQYAyJCyj8djwEa/Z2AGJHVcWU
4mCnLfylg0xQwjj30WTlpF4qi7tDg7rwcla1T2ziGxllqu5xXo0iqwSJjK4RYNCC
3uoCTDunfuI3neQap6GaOg34ENaWO3Lv0s5HQvJ/1miMitGnUYvcPvmctnrCylCa
7pw0JHsPwURPx3gvaJZei76rv8ods+zoXGKAHJzPl00lgmPdMJiS00xbAXieET8O
hjkgWuq06QUd3B7NMq3Eatz3AYH74slRFDGDiFJdx5BWKCNgIdjfbnfUiC9s4YvT
pdSyXgyxPNiVa8H0dLGGwf18pNWUHEX6AHFoj8uMjKLDrr0sNsSMMzz15AipubSk
PazT1ZHgxfZrNoRUhOFtZyV16cyFYGFyj7SwkjJRwYYgrZlc8cU9aZWCRC5W1EC8
ItDAZYEvwhcluYE+ZH0Ko6wqebMxVti6f8SIg4/+TxdU2JgR8ViiuDtZKScx1p9O
UJY24IEvkbI3dnuaX+ilGP9eSilwR/ujvqeEU1Okl0ea9kb6o56YBYqySw91zlwN
4RTWesuQghSXYNiDDvtlugXMBtTLy2GriKqHEQvp0Y5kk8OO2VBvIVR265/DkPaZ
rIgUTU72lEbR/8Um+CIirOmQJhMafz6nl4AP00+iVFGtZPnqVGRgRpFlipd6kFZO
wvpCbSXRwG5JhWPSxLeQOkNXw2DiBDdl+7UvIlTCwoNxl/nGoLmDEu96ubVXP6g/
y+fuy+J/AEldBwipF/2BvBDu+CyQqTKGLzyiGAeShmohq9vi3s9WruphBGhq7O6M
FOZyFVj4xFQjgVpy/R8A7J6V4bKk9EZ3aI1e8Q/kjfp5VaZAJqYInH/KXmPtTrwT
r/6xkQTF42Pp+XPLuXAX5DyYma7oEEbf5RTL43n6mqNpHQ9agVxoAuM2sAYGLgQf
sAzU7OSHujd3VyoNUTVfkOy7U+RDLGu9Qsc89bjTeNANIGtWMW3Le5BkYnuBgA6a
3pHk9Ai/VGBLZDNXcnTzWs3f0IaH74oAqeDFO+kTKl7GhMU2LyBOqXNB4iYe28rL
SULpufWGyj15OZWuv/wo8NbRXAuGq8mH+5BlkNDohVpqWybdeJpxorLrug6V/AMF
+B+cr5n9MBIplUgMMqwl5xA+sbfjT80tAkBvy90WJkW2pMPHSy77hgnP5Q6fSHQi
JsxA/dmczOLd89W+sqAJttdy3PZ7JuHeqptKtyNK3kNihgfPgMCkxYozBKxf6ymW
S+DYcFylAlZXXudC6YnNJGrH3FgyGpmbTfLYyCynKz7DDWAyxrYOnek6tdF6ucvk
LETICpjbESyXdtMh8/1gp1Vhfe02s2+KoMF7VXAIObVZlbbgSO1Kjd9gErrS+JUS
6i5MQ1Z/Hbk46hWrKFMS7hS34/GoouCBPxKjcf4eNvoZndkRAdUfsjZoogbfk/pN
khYSWX6gFWF2sERPjWXrffX9iDSreW3Q1Gnsb3ES5V2Do+zOTur/RphmywvN69f8
HlyAiRbVowsKoePIx9VY6VzExdpGoJjsANEvGW6Lrzj2UYUlFqnMZwe2NVkumZR+
dnF/p4wZHlopfIBJ7IwCKCRmnclHPBkzzXkqjQG7wSZ3o8jKQNYHZI4RaP0tYlbW
844YCXf9KDMRNlIx9fZs6tOes/EaCIk9iFY11FUoyL+kDlpQ+8qalee6brnLpvnr
7+tCpSJaLTufAYlAbR784qI8q+T0XONBpZXQ1+/Wci0g0IIEMhXs+KJrPANRy/n8
J5CTpPdyJBQzG91mx8I1YqOFGcRncmZ+g5CJmZiciu2vvdFrBJ7xLEfi9FMNkWpH
ckRq1HSXDZjKGATTJxgA51IxvGomYceNMI/VPo8F6sicjIFBpKyJyRJvyXtX63fD
mymiqxSXxhOPu837miwQhg==

`pragma protect end_protected
