// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
cO9NOrJjl0VJ3C5iz5w8PL3F3bKtgXVMbzj0Nx3rmT+NJL3cdRXdsM3kOnwz9nPm
RhwsZql8dF+UKhkFSz3A5kLJ4JBJ3LNMqmjA+xedX/C5B/v99c5RUNFsFFsg8gEW
fDvxcKGcmbhdORdJBeobfBrtK6I5xVZiKcoBh/kv0djsTCxHkxKS0A==
//pragma protect end_key_block
//pragma protect digest_block
a5uIYTsZWzAG56JpDnl/SHeVJLk=
//pragma protect end_digest_block
//pragma protect data_block
vuJjJdzMIZ7aP00mfkoQX7327jp5e2UL3NVQneYKWDWy8q4+XplPKZ+5b4w50tSg
Y2rlB8EIVZrK9Is5Dh5lTBbwNbaLXV4g6BoiSryVxltJ9iPOZP3ZqRCqFK3ni4zd
j2rR0pfIR+tBqYC/0Yo7tVmF1pPJnitz4NhXTFmfRVk1t2tQXuFjmJACDyqMVttY
haLhP+8yaU8mbBkdB+gvRR2cI7z+OAddFSW3KB6Udolr7NQAQmfTwMLo9U9ACx4R
yqrty1qiyfuKn6dvu67QxfLJuOjmDCwiR8NEDn8WtGzQBwEh4N/PKDwKxv3i3x9e
gj2RMwDoXkyNC6urkDhD+rH0Fmr+86isEZeqq4mPRvAINc2wjm4ZMQzPj/Z/PPcf
zHM9RXzUlsMD1k+iBjJEUav0zWt6vRwl2UGuXhzgGL1KAeI5dzT7mOp50qmY7zoi
inmoW8nwJTBe+90Idz5L2sz7qZejUt2WEtabM7quDenqfkqkzdgzVGnecD26gui9
gtkIibg2zVffLJJLnGsneM143w87FTE/4n1fQ3WHJKi1klW+p5k6Caljs06S6bjL
7SIlxA/CMGCV92U43tnzYVypSAdj1ehFwLYXf7a5ovcLrDUrEgKJfr7Fd1mUdylC
YhoD4gXuFGKa8DYdt6xyOKD6UiOyu/3hX8K+lpL0N4/DYbY8PrV4dXHF1FwY9IVO
8VySVTm0Gq0o/EX+ZGyxfoeljZI0aoAT2PLCAXtaPwPGBtUZXNvHH/Xa7kkZq93P
WP1Er8bBNOd2RySLzUHjGQRsTlRGNv9aNeLNrTSIQujgPDN7NcnMadEzcmIye0Sl
1TGbzkJIQuuY5wPMK4lqNV2B0BLdswA2x5Nr4eChn3zEvEO4RDsuAzmEwbQAwYdH
KGMBxgl5C/+q9NWaWObvVbwx3JBQet2QxeEWVprDfoIc3gEGTvQ12dDZHvdni5cM
5E5OSbIXBkMC41uLs4ag5wrH2m8/HIgVTc3f5NNjUi8g8FnrgbVABuUk3kw4KR/k
SqJ/QSNDttlac74tNDxtWahyRYAZ0kNt2YYVliY+LEhmSMDs2Xl0iyzBhqDL3cul
OMZsEZ1TmM7yeOmUMiEGO1awYgut/DUfXTdgA3jBPatOte+Rt32bTl7jIuSRByDX
G1LpUv2hhX2C5TcUyd8V0vx77LapYr/g8qvztLxBLN1nT+hz5sag/wt2oKnglhMv
lV59HEDYnjpnLKBpmaOPB+hwowZImF3cen3qEZlMy50cWz02yjaJguOcmKXZWkMS
E8/70mhQOEBEha3RYgzi1R7FYQsNrw85Xo6iHSjmFUyGSD/klJ5Xh8Pj54Y7nTf0
ig4/M8lil4Z5gVTH9mLpH1gXYkfskE6RoZbGLKbpczq/u0Bzjj31jn1cqeqSgewY
utJrToLKZPP4qdgRe0B+9INT4+rg+qldyjsGyTwZ7WGectH8CyVzdEvyax8olIuE
1BMcyj5pxZsI1hNPUTu7eiih8hpnD6j07Z45kPRtmWMTirFKh+iHyLBwviNRwV0V
x7C6MkAvBrR4Rm/Z9Zp0phUhWzSqmQ5Q55gM3xJytr+Uqv7B2sxi/M2epHFLDfu7
RwPPAFPbVs8EUGQBarQ8e7MneD+PnkFdtQtYhDNbC5tUjIYMqEt3Am2m//JeEMyn
46dve0yodLMsJP9EEloWhkaox+SLNQ04FJ2fKBotXZRd5W9FEIK23ApVFzJsOUPw
siPsR2ltvRa+35/hjFvAsgU+omjh9BEuB4SQhOLYoXm1zkngH4QJNAqpHDS0hbxi
w54UAkn/wQNaaUe2H4e4P6a9gDh0RaVjqQtpGpKYYxSyn8qF04BCx7q3/7j771oz
+1Y6y6gVmmzTZDLCnBbSlTjfyssTdjiz9DSNWUXI7h7Ysj+v7zktpIyuxjxtkbQy
hnL+WJGzaNz+I6TFJHS4f4pYr7lVAk3WR1rTn1eDZTCMccwJi8piw5dYE4FLI5Jj
DDj6kMlqOLbGORUPYoOWTJcItZnJbyTrFonOfWyzuBkOmEzKSqWLxly+Agd8kAL1
ACFnqDCGzf+bxxQ0MZkF1yU2Dzfx+9mypF0AQi3vQztZ4mXmXdIeZG/yar4MzpKl
NKZKUBFZK6n8enwZxxU9GS3NzA2bxPHBKrcKQDrE0GvyY4wGt6Tk1eyTPWvDAkcR
qOjegiuLKPWgl29LGRmx9Qfd4KnuWs8Y0C39NTvwoQYKdjsJ5vEOeqUfrqumrIjL
LnMwdy2SjVDLLUn22jKE+LIRX6cj7SeN5MiCF06v8X8RTgm8A0e93dFwpfFBGQov
QZiIa4ubnnldsO5pKTcmDqhVEC0t70J8LBUEs3v36eenue+MdFkpuhndnl9onsjo
hw3Q3aa+K+Ikp0FEgcnpbbCA57wCMhOjpiirJOSAZiLc5MPK53bLjznCZBNhbL2I
qbeniRI5inO08XbpeVUVOkTM16yiRKobBHB2I5xmJBz/dt5tYkuXoQbZCR+7aNlV
R8cAsnDpTP36eslSlKH84F16kQhgUAHFlsP6EZ70FNsQfhCDJDcmI4HSQpkCeVvQ
Dip6wsScIgtaUiV2ktDN4U962K8t/B8UmFjUHCByVWmMWnjRU2heWdXa/oGzcmWy
wKrSMkGiLQa41qkNcmY/DCQ3/m+P++2wm5GvdOsEMwzdQT4UnfGpKz9+xnpaU7rA
ZE27wciSY/+lupu5K5npOONrQhvZ2pZsjfAs4IqUlWS+zDDTzhxnvISUs0Ebs0W3
SQaVLhXDOLROEQKEfrSrBIxl33CFw9SrQFFD8tRo/E0+Toy8S4preR+3/kzGboHa
Ta3FmyGwKH4XkEFenNqpkXzlXs3dVrK2oytlhgQYuXb5ksR/Hu23RtkdfITKevND
PLK9OCI1O/73T87R2nRpFx7a8BuAD74nG7Mq+e4zIYS91EnmjJSB3CzHzGnQbveN
cufU3U2wPy19pufR5Pu94s6Tjm10wg1+UcKqasCXev5LKuK8/DOtx3YX4cDqEAWf
6YBbDJADAp8+H4YdOI6bHAp8eY224o+bJYLilaHeZZkSWOUias2cZzFXdUPidmhP
bN1/3Q0qD/YVkcSrA1Q74CbWtObh1H/dB3BriHvtFTuH0oG/TKoScjj2Vc0Q0Q2W
eJB5zQU66RM8681bUf1Cu38HE4DMngd1owUz5JJmkiq9tsExRPs5WPbnygMdfKgQ
7rqNxCJbVOFiEXFVCkKd+p7GRWM7bL6TiZvHI+vf/KEk8kWfHS555gr7bz8xbmSW
54o8rBLXvsrWQxzzKdd48d0LprtcHNxzwW6I0wwANHb4pVU21wi/krNYCBIVyN3c
9cfSEQVL+1psT07uxRrOLB+3VN1XLNcYLj5nqDGWQ/s8hO4g20jUIYISTOWb9r6n
oh4D4jqHms2lDpLX37bWrqfxgY+Ok2zw6S2mMmWJRQMEoHe1UJim4bkn1pxU88zB
PQ9rG1vNOXIedfPrmGZjcmgI6DgoVEhxYhhGDEHpI5vf8VRMPavt1TqMmcwMlhP1
3H2AeLSvRUhpS4imzOiXZzcIvqRJyyJT6pK5f2kPwVpOcDISTUUtjxccQAQWIhTc
4eq5/4hdiZm+mKuD0kzpl/+yG35JljdRAoPN12REHoy4itZH1QeClgJmmv7qWKW2
a5UQVLN7YrCQwD9bd1jp0qf6Cj/Dp9DjrXYjP+re+SqdRt8PF7WSzWvCO1LJz2+W
8zCf5AVwk7fcucuH2M3XNMJhxqGG0ohfAsIezLzncWua7N2Xt305LZpAodg/NhgS
ahYh4lBnN1q1da5GWGe/z3XSUcosMQCs+VZpcZNTST5hnG+q7lmzptqlk9KgCsCc
BK5sNjb82nOhpvKvU/Mz2vT5XTcMu46CsC0kLY2GYhLLeAC85azmJbNUdiY481Gb
He1vo76xF8/gK0nlsEOef1KSnDC5PpJDkpgusZAwLtBcPvhCZ4t1dkgxmXw7ZczR
h2JiM7XLm2Zxru7c75QnbWrStooF/4F80BcQQ0WwaNSzIMl+R7+Y/wMtkiiuYBNi
tGIC5L6QZphSgxNHPg/OMdWBwVXVjxoaFGVkZuzrxF9GBKYGCbDrueqwdr9KV/pC
+UBkl3LVn6CaHYQiDmXN/x1xM/nhn8cQoKoqY29Yqa/7CzRY3uuW9R3X/ErTGMjD
2mJ2+YxU6wKJc0lTadZlo28AbzQAbNpKJaJpLweLcpHKc30h0LxAm6R7FgRY+q/b
W/pwhrJcXTZ88Ou4LAZdxW0+BeqAqB5+TkFYjJnPdOnRLQOhkEQaBDyYnrIBm0Cw
AJvUwzC9DbUbBafZzws2XDuLKQKi6lQ4VpY3h1rg84aZ8y53sTuhEAXkRZG8cWgG
tdYGyE2V7I/1cJis7rdKIwRWY38cuBGSwqYAMwELOykrrRjbqLubMMuALxnQaGUk
DATC0ibXnUOdspRzBXUmyPrZ23+0qHqbLEiETwr+q0fuLKMob6fh1D9o6HyCrK53
okhtS2eXdQPXyT8OydiXXqcTlvQJmBaAcgF6N9/NNmk9LF968IZs0xfEOPmgwsxx
xHou18O0VxrrXigQSRbLwZm/hF5JpLlrWRrQ2tZMRXbg+hIZOpKqGmZydhW9LASQ
wJsimyVcq8JQUsC1Mk7MFbVSMnRGKjGK13CkkUMnyqu6KWdw5o1tZRx0XZ5BPwzA
etYGleLkqOGpf7WD5RPQYF7KyiJhfVVzbyy5skRCB5Zvf6hxkkFXGOJDVQ5RHGmF
wVjuQNfPHqNmdLp1Sp7W4fEkPrfnJHbewMvvyPTwNvUhxLYN5eqRUQJGluGcAbyg
GcCh3l+FdG4OYcXpODO8X6SCgez9r+CMJ9XZXIi0xTt73snX0fYxXvObyM4ouh25
niEYmDQh3407jknAslRhZ0LmMWdChXdKCpalxwxNwwvfqgvShFeQ2X3E8EDW1cAI
Z+bb4ClFJCrDZ+8sHl1Wqwf/aTIPxmjTTT823wMoAxNFXNAgmsZXY+g5r6pBmLeO
5OS3J196FxdoNBLCbwan3YCnt+YxKfSEwQb4AIGITgyFT6yi85cC8EHYVNt9Vxpc
gmSzRJgJ2kwhP6VNK1uo4ngsrfdfied89epLshybLtpstLYklYbIlZvC3mJN5o1v
v0A7yztLObzMkniwOlCJ/XY+EF2dMf+/uO6AWhXMM+OwLBTOsltlQ6A9jbs81fmf
5fSbzF9cdWBNTIbUX5VdYdrvc9BkGZ55D1uptY10NXXkIyuHm5C4ilZ+59Ah6dQ+
oD0YZEn4nAGhuCXk2vlaprPK4s4WdC9Qpwu9hBn8IZyTuox8KLO6Jw437Gnp2g5z
6CtlD26/fNpO14PlC8nQil/7e8VFESn1xhDy6OqIKJpaGt7R6LY+vxGN2W62lxF8
I110PhT+2GvMQXF6R+7wND4iTzZnNWpr1Bvh+SvVmDAqU4uVAhJoYPFA3OllnwCn
lrnOCyun/9LtVdCUWCBKFtQo6/H0gsC75S3ibfJHcCNdjX9r++PUybXjPsfYDoV3
WvlrenmnBLcD9eefx1z8EovgC9ikRkZV87ujB6u/eqHjRE6JsP0OfphbUrLczLCk
WVJOieeQNWad7f1xYKCs+JqFi54fLkprWiTw2JRc/Um43JGZteFVsPzgJEfJftBE
VlGD1kJOdZb6Ja/Qf0vs/7SM07MRNkfhVvBIOxUs4TlG2jMTTEmQjiyru2PnYu8e
8aN3Vt3wzs7Yb+NizYEkH0EE1IzvP/YurP3b5bGPaJpyFll9sKFYtreq5ZyCEs07
dxxlENA1O9rXNmgsRWbIMAZCXfaXgTnA4VXCfM7p0AiNaPAVVAdWj16yQvGBZ39T
LWsyMvWA56QbvEI7vjdxPyT9rN2qs5wI5BBXmFmLXXQ7PRc31JrFkmREfJgdCnzg
CiWjZ+KoDpqYBmTW929mwpJ8+A97GBdNLUFiiW4WhrtJnkzjwFJf1MsjrOvr87rL
/W896KvPkCkr91YH132lVzVxLNCpaqaQTRKsDGUts2fJNbiMRV7wiBpErakwQCtj
fxuyqvyDUJAfA4Qb2QlyB8EkJpPz2jFevTNlp/NFLZFWRCHVcNXFGxSYaGf1x9C6
gDHtTo0mFtqX51mlASZCyWfitIQkV7gNtMdssxj0z0i4eAEGgcgGrsd6kqxfk2lb
Y+/g6YGxuC2E8u272hC116+g0LuLAXTmiXFaowrEDnhjtGsnrCFo+RnxR9k3FSpD
Z+uldOzpI6UCe+zXiJmJHC4UgOi5psG8YaymxvwDpWmvKqOIZQW74aGt0RnjmYEM
j8en4+MUh4Zqi9UTB9U3gQrpZA+2mwTthv69PONq3VJA6aoKnUiApMEAA///GZdV
kxjRAH53GtemXYXJJDPMxEgdGoBbtXHvvRqh9q8ORzP2qzXY9BKE84yjmJekeH7V
0Wd3qF85vXcTMfa06p1WAMKARNBiH5QmEK3768A3f8fTQp+klRWb3B5huH+ur+xR
aOqykdes4wplyVjMoedCR216Df5B3ofRn1GzxTrY2LOip6ZI0yOjRTEPdg5SpiBv
EEthFOoxnLsYY7RTsBi0k8FneaKg6w9UzQtxPDDwaiU1ZZsxHsyH0Cg4oM87ScL9
R4I/kYjfJEADcD5Iq9W06DG69pCU0bZIpR+AjWnH7dKn+8FyPyEkrDCQCFLUHmYY
h/gVe6Lmw5Ans9MloeAQclx/TYifr4DAMrBr8z2WQxTh5kl17Vyh1vw42LjCo5Lz
9wiY93ceLg/C5oBi3CF2k39N02iPYSMTlHZBULzf4tBq+oxAVwAKc4orTidKWOTh
QY2/y2/OvIsbahIL2y2OEVAivL254WhOEeoZRdqGeQjKspFyT0nGcavAluP7wOV2
SSPe0EEpKuRnuaemWKaiAokRwaJlRFQBrhit48aVqQmJNcK4hyePGxdjH3nLqaZC
GLC60JWY6LFLL3a4yM2KQL+CtZSW15Iv2btW80Srcw6zCP2Z6e1F6Y5zrYC6Y3O8
Kmsnpvycb6YBbff9Nrtc70XT3yDwDZALM/IF4T+MiGBk5m92S5TLiA2iX+10jYab
57dplGcE9COuy53EDfOy3eiGoetnKm4WePq05ruatO5hcmdbt7X0iELU4MzFaola
3gYC9it087szg4gk994Sodhy8NCdnc80xZHxsor8uKSOo6UuZh53FRwBBJb9aktb
c8TlnvIvg9XP18alpFPz4fa/I4nXSGWftBV6O80bzd/yiOnzKP4KdQqE5oNHBYN6
YfTu1V7EljF9hl9lnc1kH4sp4GAtz8qKNPuKrd1YuKfl2uMlek9rhdnt/HJwFn26
mzpwDGB3aDyZ2yn22lH4GMwSSurWuDh36h8zhg/21zOEeFYjUSv176XPikOCMAJC
lzsBGNWZVs0+278uxIw859ToX8xoPrzlZx8c+5MGH+ASUB6urchfqivAOB5J5we8
DSIEdLVAe+v4/+aZlBkPB/vIPlGXNgUL8kjh/lpRdgRx7zFqSijydGrfsDlu9fVb
rYcDFSzZlg9PQi23hH/AwLiTa0dW6qUB3tGR9dDmNye1tftRpHeGMX8Ndubp2EVP
v1UEfAyyJRC1Wix/yqbnUiRxTfYKheoGdVU//vtDqM8X8ytoyVKEXQF6yoMVKiEu
rqy033NLJfboHhxqHwMDWTzXlQGT7YwAfY3kjtO6U53+E3odIYKuxUE27Ais0YKp
YgIslKAHlb7eFopfAQjzHAxQ+vqJZhAul2+fzaoTt6HpR0HO7iMUgE5u/aGATYI9
H+LAFrpD06Gjf8Y5+ALRVUK0RWr98rMgOHPfrpLQVayOXioYN1X3XscYBIMYLRF2
R5wn5lFGAtzl28HNhQy/TS0ndO+S0xe7UiKJK+GK3gx/r1s8x42hhCn4VZuqYUAT
Qp6AM2YRejdeSjDasf0uXliPxI43IiWpdYL3jHREAz3+d38sSG+YY4lYgS5o6Xsv
bNjpGtFOyC29umSslhFftnULa0/EpJZ0pH6XYQKIOoS5QvQpXgr03Ha02rEp38OX
WfLOJJkP6lji/CPEaJwDWcwfAq1RveXM4Dj1J68uWX/8vbIUycLpPDJjdvTwU8S8
mKvewDoBDEf8qcj7F8CyLrFsXI9dbkWLhErufzpFBqjiZerCHrSp9hzlLOLICF+8
ZtG/AK3fxzoaW70XCYUTEo2RjjZ7Zncg45J1gLEZFpEqyk7OWtkVM2Lmqc9wuEti
zEABS5YtUmkwS3rZKoy14dpWSExm+/Abp5EheTEyWfvjrqleAnFHLVVGYMdFJCse
RJVD6X13K+qfH3nOtNTHageT7zLBXVTvdcqt1yXsSDtQgZG7rTVmxU0YCrwRERa3
nHsLc00xIIKgNgdNADhI84ryR4x3WFVBN5pmyMf/zFbI6PZS7r5LTXUgHCA6BZT0
srDV9MIsoJYP+1OJbuRTOanaO0wnnbR7s2PhQV/OgM9Z+83ji2cL8ZAjANaoChhp
9TNElHSoe4HSPx4z2cGNipArHP+f8EzafbEAq/nytUplzfBTl2A0C5GN0snrVKdi
7svyY6Bg0WpPHAQmEGpPjYQJhLoR+8yGIykmtWIVmzoG91FdiI4Bi4Gedri7Tt02
RyL3sOa/v0wABDohPblMKUvfZ5t8KBYkcxUnZ+rjjcfbtRALvbDdrZmVkYXqMvzq
8PWxpsXgM5434Z0998OZ9R5MBmwi3spo/J8xSnQaf+buRyKRwDtpWo6eFd3ZT0fK
SYNcBACkbZKZKLB6WQRuciuiKgsgTSUsCCMkXEAT614l4ASbfP7eh2NJcEp/11P+
gWJ5SzrgNwoziXtX9dt250wyPtPVhguQORvhdLNkJurkrUgXmgojNjojVhVMXhQh
7hToCQjxNx7WYHH49CskHXPIaO/HfNE/Fc8fXtzsDSWFB+QuUfEIxPSUICjaeoOG
3b7PQ9aAHHkY5XT7gJQPEzyJ/CgSV0PfF+RVAjaTtGw8or1uBusFNphiKMFBEqso
9JcCqI4/rP0K7IyfsjPA3QJZ4iFzGkH7Zx5EAtUFLjdi1XJ1q+7xUEsvZc82Od6i
Y35r6ZS5WlG0GajMghNhak2Y/O0lgHJOk4q2+wI23+bsb8C7VIc2JqD5bZUKcxvb
VRZA+rAeptSULzClBO9nAV8NkimBeoiJpMidRdXAfP2QqTlhWItM3tDmELt9KB0h
Ln7Q9+WKZ4dsmL5LhXm3KNZMd6lDVm6Pi3/78xgaGBbRObz7X3NvrXgW/9DzpyfO
ZkZ0GhbuywJ6iFiYATdr0aFulv3ua1zkUeEy/6gX4tNWIP8kUTc5G6K3TBQuubtw
g7u52bJmae9k3+3/6FZEOpYyx7tA9sh22gzmbg/7PsVCY9pWlniH6MnF8VUosXe4
4mayfsf3qEQZ49i9yMTiD/Xfnht31dfuzZ3s1o7+FlafY0L+Mbk7QLi90ff4imYa
QVtD57jw2JjBC194In5NUUZKx1um64FZFe4/if0BVbz8PQaFwUi/xBpHoqYNcYM5
cKGXmG+tVyNmo3GKR2/0Iz8Io1IK7f8VfwSFx8CztlqmR8wFvpNQVjJIWNIlmNTg
MXxHvwnWTeWyF7ifPu+ejhhFGzMOgYnS6Qo91fQn8W8fSysrEC25yRg63MxSMDjD
Zga/pgGCdkwG2TLDZxgRc5dq2BBs7sQ628zy8iCfUiQ/ia+yT8UcLsx8s1gGWs8Q
3bcNM6pRSpzdYkb42wjsgO6+5xipJ/tvapo1qdGLuq7xI3ztZBQDhWep1ZVC0cEw
y1uz5ojzBgVpUd96e+gYpYpU3z9CMtiFBBCzWWL/Xj7HzEWmNMYTiZxjrfodrUbz
kZ9wqoXOfaRz4Az+nkkj4ovSkKyXRKobn5RBWt0bzq+tegwIxCTsVZBB8z3h2TuN
DzpxDvyJCRpY6/DjdTjeihO18sSgTqZoO1kfu4thbra0tr2KwagPwH4kz7QLTYnC
y6lh1WUG71lih3l2GTpyMQGNNFDGEfjhjDq3Ehz9H6C9NWW/GCWUs7Mb5roUQuEi
w45IWQyHU9iNrJbTHYl5fL8suj/+OPSF7OT2wAQzp/Zs7/PaXTberrFb65KGCUUy
gMjLJf3Mi5BPgrHulANBnUxBVYjLJmTrGUEKggK4bHREzs5IMH/IX9KTR6JfzAb4
P0+bl0oQ6jWRTBjNmAC7/EqyoHFxjheRen836MqpPrk/zVoYCQdOT0mVS3/rw1pX
eJyYgg8uH5nd47eCowCKb5mHKX0MEPOr5BquJbuI9q/VKSFy7YAkJl6wuUEGEy+h
TpTooCaXvqSzPT7Sl3NFwRee6vO4JrADnn1OE3nVbv3iHy/tQiYR6uiqqiytNV8z
LWO/PIfK5ww1xE1vWA5ZQleQyxoDdkOpXk6jGmA/g8U1hsv9ElJnb4Gqs5+41kGc
zEDPHSn5cKkUU5WX2z4LIfT67IvyIGEHKFcQUMyNXGhcwyZG2mDLdpP9CkIODUPN
6IqSWTUJCItc6fMpwMaeFgvbuPjghlSEan3dKWo93xT56HZpQqygmXxC3S7Jj5qr
uWVVEkBX9D0m0ffDvI2hP1ROSbFBeF2MlB8GGE0Zh/Zq1yyTbEBAI+pp4WftB2GQ
kwG6w+8AoCgeL1ikps6Jg/zcwLqkrOE/LcTow5rYpLxkDfNoJW7e0ROTIE4GGhIr
Ph7+Dx5xUj8M/hhJhCJ19fejIYtQTE9+G+YBtwQV/JfOo1/i6IK0CQHDVUMJk6Fv
f4kS/BffKc3wIMWH+3O33oOMXofTXjPndD/I+CgAvgvgC2EZQ3DokTMg+hn0NvaZ
UgCO89h8yNbVfK8IpPWZQBsA/zWegqdEfo+T1PuNelrP/o5JyPqOfSHTBy44mFvd
1eeos8BJ9hMYSk8/PFnfoRD/wnzCB7irkv0NLVzNL0jIBEZlpDdYIILEYEYLVmlx
miRpshYDoEfOSr+7RDtiE0TfFK97AOhFELumAlcMFsiYBkiSLfgFBQOgoZIiqNNd
y2xstC4lIq7epy/FRxZqfwww2E6BZB08MTx91cb2imue13m1X9bSdeDHKiBpo3Qb
wzRwLKYfZ8igE+0ev5mWSOavNZKyat+vkiETRFJ29yeVzqhfb3jDlo+TVnP/Pmrf
z5mD0kn47jkmYtW6EQnj+LZQJH6E6MpBz6Z6d1dWuyGxw4UVQ/22zXe97KdBSOuL
zTDR5CaLcMGJeXXR0Ti5oECLSy6NcljDtdyyPn6CScdWpFdgbxBzJs3RRz5UtOeV
TwY//ltUhCS/bdUZRCpJjTGxthYix1JByYFsYUwsqxGAE7eh31XKHnYjGabGLFoU
YJbguNU32ncZlM+XLnwIOkQ+qiGsHqTKbKxbSRZSdThoQ06wQ3iXW+pOMeJyfp62
WImkbr2nrOVhh2lLuJnGImKhNC1oIbC4mI2ecJz36rgcGg/ezrYWe8ZUsKPrSnQy
L+W2YU1Efsc7oXSzQ1WiGXDBgjdZPv5kirrTS7kSCCvEVKqQCAu5vdPyAvY85M7S
3mZyWqJm5IaG4Htr25ob3XOKOslx36C9Idth59ZXLR3v5bryEH2cBH/B8r/wfsTj
xKlThbx8MpoQwKqDbxbeuK0KC3k1wRYr0MfvqxB5N/6R4gVlFNTqzaSkc+KhuYGw
K2P893ggFzNb9ya7XkZr5TRXUZMhLPUNrEn5iXOrqIKU/wcQLYfqpTCqp/6Ej4Mx
oIpYESayNalLsJeIyuLSSetdc0zVUR8IwiNOJwQS4ACddOAx9bLv9VG9tz3DaUIe
omw/ZJ0PdmtWdOAH9FD/O/Ue2PLopBg+kuLiF74fkLfk5sDX/QN3tSTq5yOaTs4D
gIwEPCkh5wPC+EcebIG9ygdb44HmLNH319Ea8G6fR3vLKeb2Bgil/NSTQVghVWqa
cDeUJ8WMfn/R6ZuNj2P8Hgs8wCjah1E+X47536SvzqZ0pzeJHz0I7piTqY44EJi/
nyUrm6iRyfkszXO4B8dAtJaBP9wGQqDwUDx36+ISd85gF0h5YxYBQ9zB16Irk7Vg
jAfhsi4OTWW/eDAA2n1BhAtEROh8L2GMQaiEQ7oxsaSTCIxA1h4SujVusMZIhaLq
QM1S90TzFKAubb+/tXBp/IG+MdAOOoWrD/papZZzKkp0175aDCbWzcxt6PN2sfb9
Cw35cjJKbpa9FuqP4ahWBATsU8hBgP0Kms1wgOLFyYD8eqX7XTdi8Q2EYwx0rH6q
USTzGqTCz+3TjX5kzyclJs+6sLf87Mruc3oFPPMOYtzbT9BFwp85JLZ67YhfofXn
IIvCV5FhB2Zm6bkhgVgRKeR26berzwjbfVGAtflTEKmGoB3wYnn4x4uRAOUmYX4Y
sV4HZUCvrgTVLxhp2/pyZ8hNuJ196WZ2N/vVAwVSMqypWFcp2Ytl0GT+IEHfvheS
c+77iQM2ydpVTcRPt+WwkfpwWP1ZKN7HdKJoLXzSApKBLhjjGbBlqCvNOG7yI3C3
hh4QYNJFnjFtBu+8xGstNJ8N9SNQPkzbTAnCmX0s9L2IUPhNrb8j4uhM9Nf84uVC
JKJI2qCEiU7ZAdUsIThqMLh1/4U1OI9ggmUZObGPXmZ6zlMmcF/832//LQityipk
cuPmdrUkU15TtGozRTNk4Mz6SsAirU7a9vmG3UvcCvz6obNgUs2qAKR6dig5HWiI
+rEv5pdZAr3auQ2m6AVeVB60r5U0hbDKqMvXHSqO5BS37LdcMitosqBcPyxfhdN5
QamhYkylR1D6crzbXQgSsXCd2shZzo57hWrmswNy42XcabSNWG+18AKLGMJusLMu
VVpMWxwn7G+0eBwaCuqbAok3QtMXgSFPpOqTxcGpPBIJCe43CxugR3uyRAP752S1
9Lmqp6L980EP19dDIy5N2iNp+D2CnjuAhNKrvU8mwFs8EqGB4NEE1rYS/v3K3CCm
Mk/EFxGF0m4Tz92n/RcrWErgoy++vomj7uGftJpUKNLRP8VH2qK9KxGgJZ0KvMCI
ZsNzDet18uiLUZRbNHbs7ADXESQYj8ylPhg+GKv2MwZ9+Jmtj+TlHmMnoRiKK/2A
g/qtZRwIi2jRIy2chYXxEL2yybAUHrUZraAoOYxta6bugApDbV62mFVlNWhInNQW
peNNefSK3Uegiz40rN4TrCec/xpZuyfDo0m5oEeDkMyiWJP+Z9lLRNcg/jM+RsUf
7EMjTZV3a1f5LKAx8GRUQ5tVofr54wfFNqim+W9iYS7wOYW+gzfj3Y9VSv1tVV6h
4qPIB6X721GM2t/0FnmvryJIG2euiQ56pMqBmyFALBc79psCq3QwEJKEpaPNN3c4
90jRMfRsAgFTD8O/GzipXIWn45rI+tWe6Mb5XkVZo9wuHFh7gu1tSAhm95a/7R1u
dMHrmr5RlMX4vzCHEGKfHB1maRuD/v4fiAWwlve6Xjgzfq1Qz//Knb+emQFUZ9GA
y8p4ijdxQLR5Cbc0yj+DWpzy9grWB7P1DEaqBZJ9x7uZNfPbfuPQ3gtcp/0QzYlO
kqlferzrNz7IM+PVljE7n5+C61r8HU7/9gyh1gL8txXANH5DuLYtS6g3zQ7QEX1g
L3ftZF4hcgL56qi7oFt7COzogV7lJbkkrxqC6kcCgkSQ0jUoZzTgf1q1T+KclU2v
03j9kQqyTtOvAROem/d0Q+Ulg6wrWb+C9Albt6bgHY5r3DJ7WyvMGhzuRhLMCeuw
5j/BteWqew4eTwTBGkWbB76iDDSUu6yKXO9RNVTgOr6CR9eVup4ErlrYbXEcBZti
WJvZ9naCvTDSFjwBokjj+r2wcjwqtuuIjC1B70mCQg8RVd0ESKiau+HHcWuKFiQm
xe36APTbWbAbUl0ajLQnApADJsk9Ku8OH3Y0CwyZ/09ci8jKpE4GLZgtKsfv6v/u
5iHGbz2SRWEZWQip6cnBJPqWW/s4hleyMQxIKUDd1Bsi/nWgft/NQbvQTqkiBM8X
q12wV/yxtPAoYoWMUDU0ZzPcChIrH9XcSOWNPwCqbwuuqzrsjuEabOKuAKDk6yGl
h89RIV8MPW1IS6ONDPegaSxF8y3C9tFOibG/Q06Yki3ZQ1nAMulYjhW3fBZCpXHh
cTF0CNh9Gwl/U9Wu4/JbCpvPGpR+RxFQGyabHGPfRylpZZmxPdcOfD1Hw8gs66AG
3bkmlyeKFyw4OV4DfvEYyyrjfsHzEdQHOfLDlUX4mWXt/rd6vPkbeOqFCjgKebRB
z2w2fwaRHRDABrd6mSGowdbcnoTWPr8a+Gk8PU0iLwSFuRvibtKTtmwOmHahQRRy
UsW8PY7HCdc7tdUjLzOQZgYdW9q7fpZkfJUtpMin6Ol8PPk2J1LywQW5t09MmtDW
J8u22i+NQBgVAlhYdCjCMXRaJVIcit/icEakrlPUMqu55Lo0EOx8mZKuDnv+PFcv
xzfkrG8zzGT4lowmYH81EDBkGdl8hhYlLYIEu6VZTGR9Yfgf7i68jkx+Dv63jnDl
Kl/KGZmLgVNIZ0wSYpk5tRgcFtVmMl84mTGsD710VJloiSkUg9omssDNh8/FwTuS
DlDuzZTKAvHccZ0vUdgNyMc3sv6Y4p6SRzcOrarvNfAdp1GOEsnAbMBXDVErwSlz
/uoI8sVPl5RFWbQeLyn297aKReJTShqiKMARl/PdSwCTv/3Q1fBZ9ih5oo7wPNxh
IJJUP+O77Sr+2QR+h0JaG5dNAf0HDJnRUnM4ilkGuUdGSq+fIbxNKhsHRc2Vay3K
Pm/1S6/r3vAFJGJGmXOmDqVC4m4tApXaww7aiwGrbT9UyggKD8ja2NNKH7fTghkH
tCDJnesvYRnYtNvOAFmPqc9NXXqQ3k6MliYOG0mLEFwNGKxUWagZ59i5+dhqs9nM
0Uhs6l0AdoVvOXIQ+l3SLf3RNYzPOtl/drTQje369QMYVfA6NifqyFwA9pXX8GDD
GH82s6vMQy412ZOHNRJzGdNp7MXQanNZPCXfj7wOTCf+G+46HqZt+7QZzkuRKH1a
Oy+EhzwtirETpagl5QXzY4gTpg6DfZdbANIVvEqHkzU27YtrSFLnREUoVzHYkISQ
pn5cAweAf88m3mEMzuMJsKiWc7oZkJm7w/Dnmf6HMU3T1Ji09UgqkQ5C1c/dgoe+
zBMl4eR3yi8+2LEsLUMSgAz5g5VB5aBdVwkLO+UliXhp6wdZ5mjRcaIOrLE+wQWD
7q/PrCRIqIF0WoQL/eDoEAT4SsEiiTFJ0d82HqVe7fFkMNh9N2AWc2psAirJxAEw
S88MFkBfnsfP85Fmwq3dNF4K159bDZgiSd0vW2QcV0/BHSwWBU6NaJ2URn9uOrt7
am9byFApDdAw8m92RBforNWhGs4zTtwTaYIveDqvm3PiG4GuYYshEPvNS8ifLG+E
64tMMjzScNajXkVCLDOkJNTvL3Y9oWM/jWKDmw4KJrDIFzaL8MA59gxxmhrEDLvi
2krpcnNbWtfLpGUyd5XC+MlxkTAvzdyjo9NOIDicnIHfP3SaB/7BOq8k3XlqRZag
V5RpMKuGNZH42R0aZxwddRJEBB13cierzsAIE1d4x03jSuSX7BYEjx3UguI63IXQ
5uB4E1ExnousCjzvMnWBEOtKtPB0lVSzFgVg6/4M0KTgHooPCqEf5OVEUllUXJce
A+xP4b/szcnn4GOc35xRuvRsbD0O/bx1mxCElN4ayUv3QQtK5mOqxeMX3HrdPYw/
Vo/29XIpX5CJGpH0TPLS5RjbypPCwqRG4uwcE14whzQ2YgEBoMSrmVLvHgnMENXS
rhCyIKO2QpINN/UOD9pHIZP1L9dJ9OYkgYI78pJFoguiHlXHAfA63epIIbgHpELp
mad0RnTsjnJyQRoFEBlHlqDC0imZGgbtgyCNWagu0hZ/Wzw0vZM75ll53b45aHP/
M9BTcfzwris1y5yPPzCp1wozCQoXBBY0mZ6MXEKcVhbEwhU+ONtWdRg2l4YE8she
8JhjFkSFOdbdCNkcbuqnNBLQTLLHvP4ibYEWrGv6Ev04tu2Vta8U87NQog4Lsa50
cJGo6FMsth4c8SJ1ViO/5duAPIfSaW+BKbNPRjFsH8qS7S4jxck+LQLQHeuWDRb0
Y8RsFSqmHXkLT/BYw/o6a0l0V6JzxjAzoOnG2pF9plY1yxOKs/+UG/vaTQcHHgV1
e58v1IQX/cGdeas+ZtSSpOF10sxuO8avtjeK9tBJ8/jCJ9Fld9lYNDt/M0cvOSBR
96/EaKZaeBVkQ3vvFpW8N0AE4CQImPDuHsBQMivzQYayXWfehXMU2IUODnpxNptF
bHispxjIbDC8GPoDA1nt7wFrk6LXl9Jrzbs5IuVZyVSTAEob0FpIWB5kTb8r+4lc
ABB81WarnufFlNrS2vxFjW286I7yTBrI9Gs9MH0/swOPVPKfJS53th5guotL/xTy
JM5zmyW9xSCbFWYJe4YSZIDCWDwSn43Rtm3hhKEQ60CJEE+ySFqyFL4DUE0GV5xa
RBvcUE4mp4tmsmKQo6fqQwtoimZl4ixw7khKVpMOfg8/+U8ioGOmpIm665Rkfeqe
irTIWiMlnnm1HYYR7PXARfiR+XCNRr3dd7iTWlbiZcE2JB5EENyn52puX8J/rdm6
X6xb49IyeBaNu2GVQKpV6jXkUXJaJ/orl17jSE0/u4zrH/IHYW6BCQeY0uyPlDmF
GN3gLmtRGoGLtQ4l31F3BKPDLk9BVj211HEksJuUO9Kio67QR6bYKulL9WT9J+2V
2zz3gDQOkjAhcvidaezyUnZktyjTHylVQyD01VbkhJUdgibyhU7JTfV/LcVepdd/
wLgN3AU6LRrsMH5UJmlYgc2TC4yEbmUm/YLPkh+WM48+xMBu5SsImmmVRq4G0lKp
2FrloZ8T/gBwegQ4eSJ27ROLe7sgOOY3YLs2OwmqPGr+28BZZCDlXJ9jzb+hKe7T
ttL/jSgNUUq+4gx47R1TqZOSlihQnKO8hsEQswFYzBe74Q48uchTqWOUym6l3Ppb
NXVpjj/R9SEuHRLzY6GXm46d7CPg54r/hIsTLVL1TZK7QoTjcTMkSDCJF2xZIDXl
YQUQ+7x2d2wXtDvtHoMxmvKqsRc1mGFzd63WlOZHvhKmpuwZ8rvjm/XfRn3mbRci
bU4h/wet0OFXbe83CZ6cA6DfxitPpmG8bdmdCOrOhDK0N7CMGij4xL3vS6OPivV5
wceefFPWnZUyipKeqssIiiI+Bate2QkD+Lm21lSstwcVMd7sX3+DxBcnx6ti3WUj
zZ92nWjJH1ccRX8bbFqAAMTgVDO/2R7lfHJgB3RzCJFC1VPyPovbqSToH3aPPt97
u1dxUPuOYZdVfTtOMFhwsSork9h9fW4iAhgsMPbgTwEFuLFLN9pdLTNmn8vO1ujf
4j48JTHSNnxxZcrTFKeHhD389Y5MIGulrCDobOMgTuYaZyLoT/Ok5euJqR1hu76S
EUC5D2aFh5JOal4T/RJ2SAoAmrluYVZ0NfZrnd9A+Oi3mPIMOxrlVh1DECr526pa
gFr1y3A8potKvc//L7/xPTmgoZxVxglfIHAWSyBJv8tXul4NcgRV0skDsbb76n7t
b2F6IAXeAvLcJBLjWC+TjsMNDv12Y2tgtlgMcbG90UwvSoZ+hYQtyy55y34/jNtr
yGgXMsGQ0JuNpse+OV1gaQBN6NpNVZlefnAiYD9tpAT6hONET6nmSq0Y8wmOIhjl
RUickWI7WRkDARaSm2d802mwIngnzguiXn54jHhDWQzasGvQNoLJqNNnR9xfr0vb
Ubs7n1i9jgcZzhRpmpM74Yy/zbO6t2pog6DzHTY/VXhFw30Vp2tidn9W38tIvY/z
fTQfttCAyEahRNS4qQB3iJMYyAQrfbVI8EpwCDlPs38yUfOfgjSaNFrNxnTd3ZkS
t0GezhMyZhmGRWb4euPL7n3i8/ML++u2IB2JuKc/RlfLrUGuTjTXTD2avVNPoTHV
O3Ey+UB+9m68MuyN1bHlWGjpRVsXWUVXN1VbmzvO29IQkQ1iQhh5NZsCkq9ysSyq
E5AmjNZSY4xBgFskfW4WbRukUaPcVccQprPujrioSse2oyOizkj4Fw90TUujiqbj
ewqeC7rPyVjDLxQ79CKLN+f1gxPk/ZgIgn7cLlxSQjDW3Efb/aiX68peTyGDq8IZ
ckS2Pv/veu65GtclM22CmKMn65GJBhoFm7MC3X5AeyX0C3Jli44/OMUbjW67lnPO
ICPhaEDLD1OS7ODhgqUchhqEE0HmReEQicHtTPYx4LawXhNmcC8/syX/wJa3hMW4
kflktHR0RKqzx19co8qkXDXCoFBH715xGLJ1guZh1JiRu49++Aam+bxqVmpnzQTM
k5hxiux/MmSTZjsh90WrmdheIBYMJPlmfUo5kOietyA/4EDv4f+4LuqpHc+t8W7r
xpKAqMKw9RkSA2avp2jpZKf02E+XnNwQgyONWvbrtHkQnQ3mjl0BRksBw7ey64zC
NLX/rLwcBBE4XHQF7hwPOv3rvm+d/8d9n/x63Iqnu4vBxyHRf/tevxg7lc0B3Rl1
CMMHEpqoA+zBvAcdWvB4j7uZhfsEmUOSAee1sWCv+LOU3CY8NLOk9zwtsWl+UEoW
WYwSp+22y2MKyFMP/zppuEXQCtzKu2jYl/0nmup/LfpGL+RIVPQp8WHB/ga6uiRx
ElELgT2pylW0gwmFvemX4C/S69iObLKrKe/4gcRyYE62z7si9rdDRZONGc2ObsWC
SQ4mCTa3fVAIXZJQ128KS1UBMrf/ZFig6U0IZ4VY3ppeLC+RLh2uZt+Gp1y3fRqh
h1TQUE8+4nsTZyaHnipoUWsQ5AGhy7BEN3k0FTgfJqOBc8pq9wmdxvsDCuhNQQi1
8ijmtg/cf7fAt4b7rn4xla9eg5m3TUcYhp7wDTS3kxGKorY9F3wOXDENDwVzIZc8
FIE0A8TjlCQywRjfQAERpgO84TJyZHLnxlBg+DeNqDivPMQp/zhaXpZnSJ+s3I+y
ryknVUMCZU8aO7JKt+sIsr4LnG+KnA20KKUvIfVPNLBdLtNm9vfJT9UFqlumWX3P
3cV/PyacfXeBBMQlfr8n4uf9RXuGWZi8JBRfQbgIfwXstfND3QZXP3Hn6NU7I83z
nXPLl3Ds1vNTbM9a+GAg1AVoumGMg1xBB2JsRXS/vVohTg89Fbc5nx2oOLJEJAvx
M5hVaT/icusk+sbsKWJJ6y0EgjwU5qd7jAtr9ij9bhxpWtx2HcMCYuVlR7UFFIxz
kdS3mGbxZLSZCIzUUEHKD8e7jT7JGjpmyKR6tevv9sISdKmA00hVvVEIjwwLJmL8
XLst6r5MKnT43n11RYBGH9ZMrv1bs1ltMoY/lB5IpG3iE1gZ5e3qTkq+GR8iBbia
eKOowyiXwZ8iJZIEieA3yPcfsO42mH1Py4/aV90SyIavFivivV/rf295cjpqDc1g
kDWABc1GThJkHd1hYO94K96uZlucARyRpDwrwdyrtBO67LnD8TR0uC1mAIGbyTYT
VNgf9IljH7OLa9TDevc9jaAOGg3ETEEqVm7ADFdXK5culy6CqtzLi9GNpu8PBlj7
UEvxKvmbeOwQ/mGU2wIo1jgfcI8BFKKT3LH3oz1OHUUy4IK0df8qXypfQoW/vL9M
I3+wqbOLNY1zOD82Uw9hixjeN+55XNGhy9EByYLuJhFNYyajxe1Bq0QNQhcCPgRf
e7eZs+tSi182dLikrxYWkcqxapcrNcwfxmRrX4z0/o6THS1wznU8unAJVOlat1fW
verrrxidahCj+mBukcopDAvgrHS0XO0TlpjhYD+78HMWRSm/JkkZIfKAJCprduxZ
31e/eTX9rw2jJaD6J26brqJtnn/15xxbDMvw6GlYBYQXizeozJiLgKJTZ8GAM/2L
MO0tKmoUf1Jah6m3lu57joC9FiWk0FSHAot6n8/EekXp4xNAunP3T+x0zOpKiuka
oAJbvyJyMl+dy/kgIfjLlaxqAD0reT9L0fTJCn79zXINQ/NQreI+y83PKQa+931G
uO00elK8zM/CtZygdD7zReXsMOTcA+6kDUHsI2au6IBrAzluhQ6vF9Hpp1rMGtwM
MBOEPfQpBnoArzB6pAJgf8KnTyn+EzaUQAXlUz1h01m/UCRViEyrr2YUYcaMl8Tf
4UWD2IXVqTCDFSuz89rGCU/MvGAmBYL67l7mG1lDYn0LgCbisYhGPm2Rbx9Uc0lM

//pragma protect end_data_block
//pragma protect digest_block
lTCxA5Lm1/M0xA3YLb8WVojCLTM=
//pragma protect end_digest_block
//pragma protect end_protected
