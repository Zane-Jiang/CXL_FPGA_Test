// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
E84oXqJHw4l4CPXxmF0VS8zmQrfPMnYLKL4NFfAq4ScqTelfM9+NpHjuhwQd7Thpr0PQrdRWphPe
j5cJH+TwkmN3rDxLZg/KpVEr5k5HTt1MfuA1BwCeniWThVlfSnWTMhSlNcwiFBbmQ+K+R8ZfB1OL
+3VZ4BsgUvltywPbkgqKzijMhT0CTXx4+v3MwQbp8XWIIumw2UCVv2dnY6bFcIuUbSpa+YOIQoEZ
SL4lDnvirzSuNBKg/AVNy8d4Ud3CkxBXVPzVfc113xRZUkzyRHigzI6/RIb2IQnEC2Rq4OJFjNOw
mCC6q5yP6c6HYo6LKnRHUU332KXxyGB3+TFCRA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3952)
lobJYqsn1uDJfF6TLifE9zrLK0NyoQRDblffwet7OmJ/G9QOGzDCK1fPgmjLJX+08T6sbsXZYtD+
/m7o9dOdG7iS24fvUZ06D+AwadWZtccK6Bg+T4JZLp4c+oUo5bqsB/DVCiRWlZc5d/VS1TlZxHYs
IdFH8IzsJZyjlU2odUJMNM9D6aP3TWrG+5OC6xrFUmuYjuOCjVdHBx3ptWaO+l/c9p9DAjE12Qil
ce4+w+/0t+3HBces5OA9e28/fu9czxmVNZbIHea4UOxMx7aH7gAVFb2w97mWm7zO/2XCuwZDgJgS
z/Zsn+7edl3L/kSprUoW1mXclKlht/UrLWmXM+DKFO00uDOprt6H0Ob6A0yawwSbL77CXjwRqEeY
h/5dLYJf08m+/tHeV76NKQVri2nGEnKa2wSnPE2Sa6s/8ozlr6p8lVMZglu8yLUkvjC5sYAICBXY
FMll1V2iNp3XLTZ89M48Svcif880h2XbqsIGBi+rFsGNGFyQ2OvL0RPzYkS1kst7e9k+4LbPC/BB
qGCpg0u1kBlxymWNPs0edIk+Yo1yU+phzO0TPU8+nQXAGz+JNQei1blFOyDqlkZSEvUeJYGCrNRJ
ypAYAjNSNevxWQM8esaO82bt4PdodMJzIhiz8dnKgcoZ+c4BmA5xXf/HbNISMmrb2nNAStxlsPrW
mGWN1bylE3+D8QTztLRInBeLQ1CKQ8LZFGgXfsR6On3VDpkbR1yhsOYZecfvvbCMT7s8CSZQl1Mj
o5EglBM0ww6EENjSuZ8j5DeoD2emkyb5uy0lCv5tXxa0TLHAEsFkEYyPUynZ0OXBr2r8YwQGWbn2
4V0bgzArQRnFh8CXvskIvqXtzIcov1eZWnYYZgLH4OBv+boakUeHq8u+BNYnyrju23yvF4XitcGy
UKFsAAL5tZ0TZn7Qrb4s68fEueI/MkxrLPciGrbe4eHxkWRvczuouOT6LKl/8DbxgMeGZz6KO9dX
OeZjSzLk/Y0Npm2FW7Bb+XtHtFYKf2aFfv9BvN/QNq0pBoJ+vJBOQbIx6NZZ6HVeVixyjBK7AOde
aIvBq72mH0XpSk1k7A1O8/s7/IZYmpV8Fx3RPY9ajnkY4ESE4kktP9xhPVmt/TZh/iyMypi1WWM0
H2sGz6J/lcTXK+EXjun1TOwZW3Kpj07IXiP4ckros8nMqOEtoTG1Y3CgWp6gBeJfmSEM2TPcdLS5
gn96SmwvipSTfcbbqFta9jsHvryRaLHoNk6USuSAXrjFutGbXZyRPedJeyQCLovHApKJqkscZSw9
RXIpsHKQligP0hGeAGYepow4vDVq6PeI9p3VWcf2npGaw2bX52hWiHZNx21BCCFani7RQJYEwKLT
LUPnBD6RrfLI8DmF7D1XOlC2tUhOKdovlOyKO4djQLuLmLd/za1MZGc4IbV2e6dsa5U2CZD+imZO
bLJtvuQZeiRyLLHSAKxQygJZamoRz9c/C8GlvCD44w59pas12/eSzpe4rGYIT+ta1v1BP9f4Nwzy
ISfNr9CDfTbqEEUixDPONq98ni4ijFPOUVTVyn9uSMeqdgMCJU0UmV/HiWjuV7NpdeZ43PXIo06Q
sYRDXqElwYAouaeXU0a0DT3SPEwRS1yeQVs3BVre8ImjZ9HkyhWKBkiPGGiZZJ4NSLgIEXXYcpIy
wUJAmahH6huDaQEXF05l4sTkeiCFxr6SmDSuEZ7WYiGgfCVTh2devSupfzzE/4BBNSAbS+JRUUj9
wb1Zz6CRuPQbnPR3yfQijnHcbriCIptMS975QBNeH8YY5VPI8Ntu4gq14QkYS0ifMlqvWYjGF4YU
BCGgOC4umH3ebX++E4ZMaVqgxO0XPTxQDkpFmCuxfpNPxQt6iBbmBguwuNpa8rz/UPp1HkfR5wDV
onRD+jY2WsD+qNi7MLqqHvts4qbb2yFJp0sx27wYZcQ85iEg0h30sALh5JEvkaCfXxx6JjnWIn34
1/w+ezo4vffDFyW8/ZHlEPwfb9XVHYoY2qn6qUohTc3fsXKj3zwYYwkYRy9QZ6XKKkN1wZ/d9PIo
PqSGaTB7IJ8vuuC02GviuHexG1dkEm8tEt5HF4so6oIyMfNwG86PM53ZoX0w8r98OFEjX1zeth6S
jecJyj9pWxOu5qnO+hzMFSiwCo+PvJjLcXUeeGQSfp1h2xnqN6EFoI5DKYzinAMr/lf9USpcYKT9
8HeT6JiEDkliG+vUW5s3eyBxU56MRC8z+mrlyMxoy6xjCZeEy1ykwcHmx6RQsq2y90qKVlvDOk9l
zbF9SRY3bZ834p7mpGDm/cy2h7G4WRf/8V4VXv+Ou7lW243gDoLqXkoI8EhKChL+tw7PjfTl44m8
SJ12PXNupSI8dVIU4vKt3RAiv7dHLiWqJAV4dDAJM7/a0hKHM/gXeASQU0J9TiL+TgajNXeDXKph
f+0iADY91+AXC5uwP8rvaykIrDB+JzcWSShzuAoudryVjFpHEdYtGqVZivXVEwqiLOQG2Dp9iqYC
wYBASJHmemwRYFfUSNIqJOXflSi4/JAtOm3mH32+mtBzdphoHapt5xNdbQZxp3TedsqK4OAuw0g0
ZQjixO6KGl1n6BSX/MALHTDdnuaLP3Dy37q8Xj52oxdAukase2OoEUpwR3CuC+n2qQPgeowujju6
vhVJKo7KnERDKECuF3TunsBA0kjMHTlRsz3aiHjQvdOaes9FbkcLBnv1diA3nEcrGyBHOPIXOIsZ
5+Q5FZZcf0PvtXqgZpzvJFYAC2z8wYtRu1aDnP09N4wyV50OsZKCN+mwRLZPs7aXUnP0Rkly3voL
iJCV374CwDuB9ygirlfYEut8s7p8TG3EaszNiBbYiqYuTPGkBz/b+FN0pGQAzXZrPFikLZJ9J1US
Da0RTbPjpB/Idpb4Y9pcHPnfwtocj8XYVdFw1m05PaaA/MOKR8PgPLa1TmRcikbh0KGyN4nQBG0M
wYgXiFxetseNeZCQHTIzb9gctkWGoPX5KvG8yzvjY32TWJ6mYMXo1GtT+HK4QZDufygBXrjk0H5F
ExLNr8YPA3+uCi2MiX0PEYTTiJB5ET2KmdiKda6jDXILWcz2yxfUif5dZMilTTZeYq6bTmBV4mhp
O2aiJER8JsFDnbN/Av0EwVuJbboLZUR6ErxjO8vsGXqtgJkQ9CB+t0PM9ZWUCzT6dDVSg/8qtkak
g+DQdNwcwI6TvG+rzzvAVfyxKDLHVnaRMAwGBon0XSakZa2XymXXe0TFIArUA5hdWpdCiF8ePHDI
s/L0O8p6BfpCBrxdNF2+UTr/Pn8WzhT1UVfkE+CXG7+FBKp0XUYM6iRzmYXTY4t5wx2IlZvdp0Xa
DXvpG9cPg6a4rtJG/jtAM1VRiIdp8Uf0utoh6AaJgu8SLOpCJ3rUMvFvHASrKtpGiYmjfDjJx6rN
3r0uyZia9K1IW/D4yg+KXDMUO0q6mRf4OUgscMOHACECnBhSYTvRnIOWj5pqeD0+D4NizyCRwkaG
3r2urcg9pJwiNdvhsNTCzC3kXXuYnYGpxJxby4Kg200EigkCHxXFH2Fj5ehAed+diT3CXFQ2rJ8H
N+LQySd8EdHiUDvdJo6FB66kwy2j59JXbmfF7kaAQmBmoEbouHBcKYnJfRnYZRWWeiPsV/8O0AMl
dVlscVz6ho3UPv6RJF87SLaeThzdDMlC1nREiW8pjaJga9fm9CLNeiEe/ZFlsbkAuZ8JvuwO90nG
q7wQvWE3FMdj/0Wlc46Yt/D9KWX22oAP7gaYW7v18U7YzQaITXz2rmRBZIDNr1jBH0rChN0QjKvI
DrMeTe5Zo8D6hcBlOzP74mggH2OeojSqgP4ppa5AmldZc7L8Tdg02HRrczw4xyqoiTGGX4+KxbOK
6x+lG4LHzxo3aJNFQhbMs2lmP+ooMfllQgS+EpvTVPeJMW3z2rqrd3K0UlEt3rVORKvySHQsbqMI
uBQq2/pdrO6hGO05R22dVDJuPBf7nIDse9Up9oQkAgzZOLmK19DWGz3TObZiiCAFEVM1X2G05aEH
VysDC0cWrbDi2gBAaAxNW6qI7g8fbvk+9KGe9Mehazr9HTPbAhfk3oJI/FdeE/KXlD5idrtLCqwx
GP4+w/UyiQyDRM4R2aomD6UH4ymWfBSgKlNI9LPPLKli1TEdfPAFFF8v7cd5vR7Ifa+uq0iujcDl
Wr1ILfFfhCrp4VqvpvVuh6+96JcPTZlhqTS6SqIrXtdPLeT/n33/snhsAqIu+j4mrM4M5IQguYR4
XbVhykVxDgr3Kg94z3/SVcoo8hOyr+qivkx/eRnZOyx0KflNLQPC/VS9HvIfRuXarbT7W1EVj9/h
rvdi4waQvDj5Y9aT3K1yzRJq9fBnTD602GqaALnGmVExZxSiDJcdWtHG22UVYHdU/AloJJH6Rdgo
OF82ckRyhBlmKdPWdvhFDHqGkwH+97YdlalQo1AwcSfYbql1NYoel06eX/Q3hDWenz2HZ5zY1LTP
CiZbPslQbSQkCkaQvUnhvdV2/uDHO0JTuKY4eQpv//zzoEhG0qKd8zEPVXcJqpjMYuCQlG0vMVFH
Z5p0mSV66UArWb8lgUCIsIgEgKczRVQ7ki9iru+eoVBYR4udkOeZB6vl+JbYA9FQ4ANiSqqX7XO2
MWHkHIvpjM+RJRdwWQZNUDgwxHG9KDFZFE8dBi8KLKhJCGq+X/LSXyuIU4NbbmCIHiowd311wD/3
z08qd6Abu12TX95Ds9JZNwlcOZgtPUZ9IleaL9A+CQXJnADZR9SlC6EJ401cDC45CvCx+MfbH7R5
H4YCpvGYiugMnrbE7rqyGvIf/CIPUMumhF+dEIx1hrHZh6Xj6sPHKnpncfwvNVpxSXsqfPbDOgst
s4xcxGSbQKlgS2P1VfHPXzhVTyiOTnotOcv41RitKtW1gLJc5PFPfiQWHHpbh6SL0EI+q8CHL2Mn
NsvkGEnhxx8JL4BrOVewVyVdXFKfn5P2zhbGdOzcYNQrFAhwLJPgnO1EbiwnseAlOlUzytdZNxEu
VGJEADFhOiptsxdRbSnodsOMeKXGV8hEldGuhP4rlxSbRrghhai/mEI4zGha1meDCvnWCBwSpOes
p4tEFK6cmY6Tzk9aEcCYqT6vpPRwPJKtSB0/UGPxRt4tl4ibtP2dxMwbwABS9FN53YSrVXN8IZvc
Zu7d8F+zkUWDOI69f/ldFBvhTt2cyqhizIToLrb0ax0UY04A+6Hyy/Qi7IX81Szi/TrE+xWYQ8rn
hOjglU/XRdXU8ihjME9vDeyhuw==
`pragma protect end_protected
