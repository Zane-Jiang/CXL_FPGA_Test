// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
LscjbBnY48Rn/tmJpsTX++aAPL/iD2zvmCCf0QAuc1zzqBhcE9mq1ega5LsPNJdq
Oupw+xNP5sk9Npn/SbIAv86tghJuI+VGMl8pAjXKbnC6HRVk/mDoX0Vs7PA0OKSB
U5wzBSN5XBHSlLcoyf77/TnVmHCEPcHW4QgmAuW0Y4o=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 76880 )
`pragma protect data_block
Idz4cSN3r4Q9W/2GMUrefl/xtL62VW/vw2Tt10ipALuMbEsAYZkHsXzzxjvDqHJA
B4iiN84LxVXueHRNQuW50xLLUWDlvdjs66b257wN/bDfMvCehBTMygVZ8Ho7no93
2KEWRwD+U8OOGX8Tj5oA+GN7siiSTsPzsiAa05m68t24gvvpjgH0Tigbples0r9T
8+uuxnW9Ke2ynvnlc1mzzsmm2T9FTEe4/sWsncjRkg3CltA/7AwQgv07EIfoE6X2
q5xEwhkg6tuTqnlblKwDJZZ/ebft1wqHe69OOBmzgJyaazEvHngsEtZb4l6Bi0xx
LA3w1hVFRH4Nj8RP36EdrG52Trmh1eOY3Nl54XDfAE1oAaWfO/ThlAA5b+h1ibxh
wsazVGSse9S21bLdCHnGfwElF97MiLgxCgHrpcV3Ff7HgK7+3IRV6U9F7Tu5sg9u
awz8Zg4NtV67VTjt7FicTqRytRFdVcHUONIZGwPVVtjxeokq2g93RDsvtbMv7tF6
ozq0G5Nl1qclvNUSnIaUoRG/1/bM/EBZNJHvOwAL0YzVxMoFXnmCTu/kglOyZUgy
D1jrY6tSjZyMWO7fkpWBkhSmkMfCcLQ/LODf2sGKZNnRd+xGF58PaGlQWNM5XWEv
1VBVnLxZj0P62z7PTxlYWuRKwCgLg/VwS6RtmaYElt4hqowBSvb/gMuFHAYY+e28
Os8oRUzKFG0aZKAtGGjDjJNpJvPO6581sf08KeRaZI9+i8qbAyc1fzDYqLXEVSRx
3o046XHhjH2mSHiKD3OZ2oLoxY5IBCs1ItU5rxCnmQnVYwsqoH2do0j9f3ylv+Fa
3ZrqgqzlZlbCetZOmLbUs1qQ46gFXv0JpNCy0SdkLP10/zKYuU948fsMqxLtUASC
ziu3MECeE+/gfSBqmRNKgdCcn0CFWI4LOwpoZGw90hkAGrM2ZEqDQWhTYxJVQjer
DjKZpQ7Banq7O83d0x0TWSxFKyPH8yXsKF/6EMnTWweYzts/ZZz/TrIODRyWEIYE
ixdEkESL5H2o0Bs6PU4VRK5rGER/j7EZbRaiog32djfA5dRpjNeWOzl0Oh4/nJm/
bsUish7ibecXs0tmAjURMKNc7ijs0rdrlbCvyF2J8VXKNVqIAYQsu2M9YXZWUbVE
ufhzummO79DV8bjhpN6yUpC/cvxZWps5QFk89xdkkRaxOIYeLUi52IP4popU4O64
f5N6Nr4xh0CDPR51ZiVD7hewtjTxYgDmINRRaQgvIhajEmcRSehshJed6uIvC9BT
UGjiIpzMFxANOXvDcEOYkUWIcYFgnugn9zedHEAtYgs0cxZSR7L55CcpSOcvxrQO
DdiwGF81jwC6P+UPX3BC235QXQh1Pec84EXTxd1TcSXf/WzY7dw9kj7wmtiSiVGR
VewVrOqzxmqa9yniEks7ufekxqWNPBxCv5oIVZrpf4uFqmWLVM2Md+/OZwhZmxC+
iXPFkCMQT1OLGvXtAlScjMf5XetX4tKsELsgGZGO6hu68HhscGzCJ0x5kaKtdwfv
nomdFfq+gXLM4JU7cskFWy2+43c7OPJ0atPBMsngWEt2vKJSTtfbzXP57OncU1cE
LCxOjtsWsVeHSmy2qWnv2o7OCYArdHo0inHA0SgLp+4TAIdAUnz23n0iaxx7DS72
uZ/4y+kvTbO83FcfDc8rt7XzH25ZTRliat+ASVl42XlmzLxQt70YJ6KMG7960z/m
N4iRwaHJYpgXnHZ7BHEniMAUoaUVM7yLz0PfNHYUwXP2pQBm94ugYGQNE7S2lvw2
3g51p+IhR9+85/LIjrkcjC0/CAQMto+VG+KBiUJjgCD4jXtpGM2mJhBHU3KS2kOU
XSe1n0w/Pa9ov8sVZxGU+GpWfqVILvtHJjLUVYO4v5Qlc4HTfUyCZ8BlViQqsolk
YhaA8zbRj8BzRVCqJum/lFUzSKgTr9dAWSiUSwTjVdmfSe9PvIgScOmYFx2MEWmu
DxyVTylc4ZeT2+lf3O/C5eJcY1SI0YBPD42QF9qmjB2SuLBz5Y2rialq9Hp/Tc9p
au+rMDYIdgTUKjtf1uRZEW7ULTZu9WSiD2uoJgJ/N2JQ6pwWvAVGM7qQ+dhbi+n2
SGwsNw23Ez9t6tRs8+Ewi7q1RV2TOXBDiSZ9unrYTwFAr0m0Fl+EtLcm5TppuVYS
nmy9sCHwCYt/JtyzPpBAiIeoaa4EcXDwX+yn9zSuD8dKvGSeSXe2gHd/VR1EFCd8
Ryij/cMnx0GwYBA7NwJIkeh/aiqtZmkMHo5xxR8Rt16yknEk6JjB0BM1W0ndhN5D
Cwmq20i6jhvTlqaoHvafFpdtoQ+4bWUlxbpvr/LFqSvDNbuLR1F6yT8g9uc2qpwi
3DBE01JZp1iQynaFbqDImn8vAHtZRESI6bMCv4ZoeEYd909LTQZKY3aj0Yg80U+c
Dk5tyvMxohQxFsrMAZwnNfZnMrMXV+/5E/OtM0bQQpeWlU4AQnNude0Y1xx/qYef
IyJBkwyAi4WTDWt+qqb0CY7w9NY8+a9x1I+97w7IjJcHRuj/XMM3VLZFwGN/tOo2
IMQi81gRlBQ0WN6ztTwNkd6d5bJB+xOVXT4D0mtu8S77LFAn+7Qj72a0Ct5iwuvN
LMLmo9p3qW0qRFV0KiTw/2iypkdgtVHvRaCPg9mMXKs1c7Png6cvMkt1iREJVGxj
DPwIJCD6PyG3CtPbP5WUp66DUWxo2TaiutG7s+0Y0f7LYaLOFSEVEbBs/misW6O7
g145LHqpebmsKz6IkMwOiL5TP4/tlOmjuSvib/Bnd6ithTsWIo0pIPiABfP64SBe
pEodSs9W8rYwf+fu5vQtuYb9Z2vmKN0TnNcjdFXQsPoOaaIV6uTZbcY/wa2sdA03
9l42njFYYW+UF6O1rrC/NxdQ1+fqkNmhYVjzCDCzl8BS1cfGN/ps/tQ8BctJA3VF
ZqL6wK3kxYmUEOUiSNbl7o03DrKtJ6gFBZ5CDppAnu2Qak4StxA2/1FCU01Qkoxa
glR4HLSK79+W9aDlxj7uaq5rKc//BLHxjzztcoGqhG/5X8vcH4Wg86Uo3njnhI4G
vjhhz32u3hLfVjUO8Ei8d2b3rPxG9BvUn3XqvUn7+VM95GuVmI+piQeHfQY1czJ0
7XjyLuGweIWBiSF30ReIrGOFDFCWpMWWOmvsCkhQm6zEAkIV+mzOOFlMrwINa+aK
JCUPx6N67T/EGU0Wif2Lggc0bX+vCkSMnzJwQC0kNN/JuWiGi5dxTXypRnmFF8fD
GAZZU6AneXrpUl4qcWTZwDtaHGIDwPJwnToMJjuSEfeVd9/GOvvFcweipbXnMk7k
F2rORKKKBDKQ1ePSijbZOkymW3b3Nn8RGLYkRQZK9Req5WuPAXb0Kh4LX7mFiUSR
oj1IOsmrJRMNRTcMX/9I+680rNhR+wN9pCh5Hanqnw3MfSTnvQfFMugcWkiQLu/A
+nAEw2SaepRER1jCx+/VI952t7JyNAk50ubWQBBYbGgW/pR63kQw4h1qtdXZA3tp
PK0roL734wo6hVDIskv7bBkCEO0kdNoi7JUx2AcXuTrdfukR8YXDahm1GGGph+1x
x6ji4tdyTKzhIkLIL7dCm+v1iRX/Bmx8JwPpP0flHY+WqmntUkRQ3OtzH6wuUB6i
8ofRvC5HV0Kg01pKlgx4SNTgGrardKl9gI3QbsvxtJx9FREsPtAhyxuetKCpT4Wr
B29ZBchHBxzyuZah8SnkzgunCxgWtMfIWeAr2OpizLRJKmN73lBM7rMg1VW/r964
RTtOc/a+G1DKJsd6qBiKVmDvLZDKKdETzEm736Dyp0XzMN+DIXoSCGhauzpHPeYy
PsW6UnTh7SAu9tr3UOW6fsn6dy1DitFThP0XQ8Fx990m8j4w87pcshXUzFJ48wEd
rq0RCU9DPURLiWYJ8r+u93Lc0y25vPGSWC0o73L9eBRpFyhwxItA03AV4lAtDjtY
x/qQRNxaqHvDeYGr2JLCT/NAgm1lUkPOkhryXlOu6KlHz2V1kqaemtOHV1bRG3lR
odI1gZOZRnWufirV2EWY2zcc3i0P6PBBlNqlu4rGf5M4w5EpbGaPDXR143VmagtL
TN4BdhyU0B5PTxSMEMCc/2MYflGKXO2eQB4Azzux8+7XoluLmuJVhwJerG1Z5Rgw
v3YWQMvJvakcWTVbPdxYk9Q0MayL64X4JGqiolYDPN5f6qKLxLSuZMGGXpcCP6VZ
qDz9360jz00eGdIFSEVOZhu3QLwGJq9GOuIaAnlCQvTiz7DCxDXbHALvKMfcWrrq
Zl7cRVJLJ+bKR77XZW0q+v8NvLZtIFBeQsCZjFkYPPmjeQZO9HS5VegxndeZnh2H
MxUQTAf8QpfRQSwYUoZYx5JC0XBLLoItxdiAcGMN2s2VVFzXmHGND/E91jkRDgud
NvI1lGXWK28DKXhK+4IP4YfRVipgkwK0E6Y7ZmBaPVVj7VimjK75SjukG/6WOr+g
HdK+8w+F/RP9jNFfNW39RzNFAlUxWd1OeilOTLzg4qzg6R3z2QNc9d5cCUUcR5Mt
ZnE3BpEYraRM0x3pB33bnQqoDMkGX0dDm+utdIqBbYgzb7BytbI4G7MY29PKMBo4
rumGxYbkg5tLDQK1n+OVXlvYSZV2Qrc3TIZLRqG8WyxEQXA9ldBjNBDk5SLZHUIR
Xa7aGOlDz5ghLTPJ7/5rwAhX/+I6y2KBnEJme3Tl/MdD9ZQyUzGmFOJ3v6dOHqfO
EWhZP9c/0XT9ttFqu3B29iVnS5w+BxI7FobZZxXB1paqKUv6+1TfZ/QyiyWhjKN6
yMInz1CF9tcNb9FfPtuYmq8iGdrsuaJGVklwGfFaQxLY5oJ+2zDvqPPb1H7meXcO
bcrXJ3Oc0unrdxxAn6WgcTpsLhR10JfzeWoN/PTNKF0g68MeRnUSJb583qwAHL45
wXMw4Vv1pc31lvFq/oY6/BipKTFs9rvU5PyJQD7qqlrMJFUiBI1cAK1jM3fkCcyO
DJCGL+jQ8oKndQm71WELsDTchkdAWhM8l5QWkmNds4XauszETWvfI1VWAMx579BZ
c5XLtpHqWtWJ8lQzISZZJ/EmKii1eSVPOtcADitAHuLQSISxgMdx4u9yEyNxgmc1
ymV4c0CCwlIRomOIYtnsrrQYH8qtH/34hdRUwxrDk0p+RMkrO0U1J0bRuTDWiLOc
Jyhw/O3Kn1GsgBnwsj4ystrX7RLOdfbF2hD50mlijamBkHDoJMTthOAZ/wFedhF5
GGRU5hwUrBhD5Yz4s81Y80ZzUVcPQsEc6UnuxeDpvHVeg0vEnzbIcz8Spc5qwZmT
gKU0is9aY4XDql5hnSZD+ZmS7tfmK987j3WHJusJqzLTkmlakypPJ3D74pxWQAnT
Xtd3siTTcd8J0XoRMlcsakDeJ4ItXHuckWX1LQrE/7fqAJa/u4FvUjY8rfdb/WZg
kSK5LKdjwBd101Mhom+VqJ1h/fruf2CWqbIiukml/F3mlWPblHZ2Z2kJCg7UCcDT
R3Ku2x+2kWmsNPZ2pwmrLtX32BKbgpeMt5na6xvagD7jk/dnt3WdEoS6LfYqU8NS
BqZIuN4aMfnzuenW/cnIT/bS+bzj1JAlCwtlW9zcJ3X083GLy1o57twqtphLwh0z
fanzEjlEWRacXO/NBSz80StLh6GwAo9XbRnEWqpeqY692FQ2jOIUZmc0/lw1VHZJ
soqCW7kX+hFCGu+PJSfjBC4YrI79zUzyRivzKF+WQGNzS8G+Svt4x2amqZdvcJi9
rH5gqaxd3MvmxGlfOMvPF4OWAyVhmzGKm3Sq9Tj+lRZqLATNcjv3m19y3e+OJPeP
AEJPp/bOAMRarkjDI7FwvDXK2qN5L1uMy6LbT4ixoLRsKJ3pxsnNho1u3X7Aeymb
kR3crkz6Ann0NUFqVxucptcuhbJP/Eifu69iL5hdPFoy4gGy9GGZL7CszObbd7uC
E1BPZqw0mMVKh7DlPdkJWZTr7I5c4gZbS9/DnXrMhVymV7fp4A0hX+0ZabGvafD9
sARyJ6kkP6Mnstmg4NuC+culgri2jQhbGYDNm15JsYLDqmaTBIwAKd4UauifiY9H
JLq22Pi/ABlMoJZ4Vch002O3AZUqjUGUwqwRa+qT34XeamnjjLjWVwaTr+WNKeqi
EgCaHAFaoN8FZOi1W5bxXxn1yk8Z7oKDBMlhcBaoC2GFxHOJXUa0ip7E914uwKcD
crsGaW9bESzpMc3G3MbL/09/TTbNhGwUCF1eNiGpiVBTtT4tnJmdysDVInPLMNzC
vyfDG6KyXItAy+IRgx3Xx0K0YOtCjJdfnTNLQuxdtatnrMqitMLxv8mxKwWV74FZ
qYHiB+Thn9cZJ9x/LlO7oj9iQT5sTz8a2f1Pu3u3Y9E5pp4YtMiydzMdW8z+68eG
9Cde8VF4UUS71ZlEFNaPg3L22jW68AvhCWmzC5RZMew9BYaqXg/x+Iy0PvmGHznN
87JSJrlfs8lJ52ktwa7b7erDbS7kbVo64zVk4wumylKKqYSorvsgpx3Y4kiscW7n
B4LCnXIFto9jKXB7UM9yVGOWbQAOsO9llCvZUsQgunCFBVg3mc3IdwSxnxzAPtFJ
YWI4PnPOrZItB2XhbTVI4y6/TvRRUICK+E8SIDjIQEZ+0gJt3l9SnjPBKTLtxDSF
Z9rawzpNBpG7BgeZUa2045+CAIm7+RTxS7n98Nxi6rgi1n60TBHDrShI6HRRxcE+
3MveFRZom7okDgPtreJmqm2MeulAtjQ4zoBbMPwRre3xygA1Old25F3Zo34lU0Ky
56I5g7kPK33acUxs+qDRcZNEq4O0irSlT7/+YJ6gKH3JUB/97sZgJWMDJN+8ZXjo
OnltOs/oABuhxynlAvvPFQ/5hw01U+fFg7iIvKervryyU/zTACdrYTdNLklHYHCg
q1Pp7B/WxN/uouVDyIcdkkHBfZ9UqNnxEhBJ3f/C6776jIDOJswmRY/iSWiRJA4L
ffYdMqG5KQzLUddGM9CKyLV9OdSM33QUpjeqQys7uEttOU57n0dOrbea7/Qe4DTK
Pu1hTqqJhbyxeIpDk/NiznDkDhcwx2sEq569cBb2u9pAeiFM1aFRBHt9I+M9XyZ8
4NHTZG42kWo9NFiksE0uBuDu9NytyonkDkAO3t4AJFAJ0oeKMMUo9ND8ySOlVbyI
v2SjzYrt+9A4/MSErMTYgt528Pm9UO6mWyRLhksD/DTTXUnAK6fqgDi0rdbVu0vY
U+HfHYE3rXi36jZ5cvfi455C5B3/4/LLJBn8nmjjgepJ+fJ4ffN1Vg7c9e4lucm4
wgkSMin+fdVHD7pLqCbzB1OcUZYe+RQ7qI+7nX5m0rdWFEC+l6Meya2oMmpo3LjT
t7ogNflT82/Sigc1eUfNVKT7bgSxN2QFiG9X486oZo6rw+I0e2/Zrcl0GC7DU6qJ
5W6FkImiWm8xwdlcrOxim/fKdp22V8DSKkPQkJm7r+f64gj1iM8w/3sA6+d1rp18
845QodO3lC6g3bjT5i0gkdsGbqAaBTIQ6/kCmEmufipO7zjwMP7rou6Z2DUsATbe
W2c4UBnby7NjDWb9VHIadzD2HkRqJhIvD/uHqMBm5jwqj7d0UQg5RBDrfgED1Fhy
vsoqppWYCeOHysfU5HPlcLADqT17TMKXAKkLtH9TOJkKApUzPjERbb6igmmUg+cR
T/9c6KH6FVI9caKgmZ09pmUfIwjCZmWcNhZvbAixUzmko77ymBP43KgMVJ57sYGp
TtGEIYETteYq5Xz0podvZit7c9OZVIIurS/yd7cJDBkhBB6hhCuUxRMj/GuqgyGT
a3l51JaS7sB94+T26hjhe63kzKJwP8nSz2gWCFSoowoiB5Bv6mbA5s9YVTmQI4WS
E0D3wExyASsBa9v/WTHf41kFjkb2zixA0++NBXNHyP29d+aN+VLwpgQ0MrxDtr6R
wPTbwnvAxjABnxuA0onLJvOXGZxopwOHEHdz6VSDYIhJXxaqjvu8CpFaMENLIjcl
JbgDZDR1BiLkmmopp8LfLwc48PoKFGt50hZYtGzHU8nz5qrS6ywFKKBrQC/K4nuz
+I9n6XTw1A+44j+0zo4/ShsMocAP753MIked3ot7ezsnkGjXmQW44Q1Zl/NgfKO3
BQ0MiJp2HiVzaEijCa78hDemEkDQYTT+KfQo9cmHi7OViQpRI8tkJxgqFKu0Zs7G
XEFICm/2+mX8v3ZAo5nc+zN5z3jjota8LHDa9KlS30lsMn1APCHcEQk/hFErb6y2
j1pouaDHLnWseewySVlLm9cN/7kMWKSEF5y/YJxIEIFg3KDrficNuG3WyP2FFUUe
5aBeukWGPMaEq7jW9CFWTrmYWYQcvp6hWrY8A14yH7N02TvVIb7+wTByiwtTkSrD
f4rNDd9VYU96AK+C3kawMyP3QN4aUOfafVWdKdiiU7cRfsVXB+BCQsFf242lpEOb
U2Lfiw2GbSwTyU0wh26Zilxsa85KUOVDFyw9fnYPnKBssN6w9y+yvuCiiwYwmD6l
cHeMTCIvS00JwPM5dlOSEggu6J4bJmUBJvIakudBzUAxrxpaVYKlGB7BPae7Uv4S
OzaqVWNDW4IJ37fWpx0VnoK6925FmuQ1N7UE1YF6zyhb5e5pT4CW4m4bDg/+DVBM
wuvqGfe3C0xQZGdJY8yzd3+i276zSn/oncW7KHUom+Pr6uETNLkjOYxFGwEX1Jsu
rya7ZaPosUr+p3gmwUhd50JCNJyUStNjciPJZFMrZPQmB4v+ni2YJyNoBdsOvF8E
/+nEBEoGBzD/ZplHAKLxq4D8Ty3USece9yGRp6JTTPuzV+Jjf+ukWIUavAVKq1Pn
Z3DcbXlnLBJlVmwYj0TPFPisXuEEDlT4UBrzLjPvvzYUSA6Og2tzb212T/e8OAAK
BfRrrHQKB/WrDREaHyKm1j/m0U5lkS2SYi1wIslS+KcfDe+Cs94OUFmdt6j3gSsT
xBXleUOFRyD8G+IZeQAjbCTYFWHooTBwxv4zUN8wOQGupmNal/NpHiWxS0zrh38k
xQvuTtpw5g+ImPPLysrcjGLzBwFdalQGzMjS3MXndwTqzoiNo0Oxsb5WXxBE9ixZ
uROmVzYLu2zmSlws5t21A4MLwFIkBdHH0E2gNAj30TMYWA0um7Vz//xc6UhitXIS
7nQJ/4dNut1rk2hD7B3ITKtg/Hvln/ZLrrITYMKEa6RnY1cpe8607YipUe5+20YK
ckX9kSLeWUdx85vIJjU89dUgdGeIol5GA2ASDw4d0Vie9z4DnNkes10KH/rnArlh
T7kRoGKxBNocNRptPtplclHs4RzjoYyuEXfjuhwnTvZfImcFB20tX2yBPWujWvIT
0oej465QtgKgPAR2GvIw8psQ+HKqvON90dp5IGADbAQrOXR8ki1g1U9Q1tYy+ysM
p7eiaTpzeMuj6JkG/3ZRO5HqgCB7v1J0ZzigdWDPHu7gHcrBKA7xcEq75Uc3qM/Y
GaaO2ER6RE8+17j0WLZdMym0E3uylE74C6KabH+5OtANSAlylmrmhmxUr9bAzHjL
+9XgGIqfP81EZIYMOuZtd7+bEZEIu1R95sEQQXWxJbUnhsEsJvcFsUPxEZGD/lNB
bL89T4nHjy+WRPUG9Jpm9PUPuTOyHSpkollIYbUG15MewpHm/nNkRSaMwIqBi8JK
ONeeJfFr6Qibk7I4CHtC46KGiqnrqI2HG4Mndg/Oi3DePiS5aC32aoXTwdXMExxd
f65BY51aecGsWSPDqLe0r0WP0z5/aVfKBiQxVoalSNPPjrnaGGUyzFuRCEt4bL0y
Fs1D4gFj1JsWHgqISXvpVS8hyLXL483RAOoWBzkaF/cdBeyFGmLqbNOEIyeVrMgP
1h170FWm8TBjASb/q3UvhECJwso+cKRpK9msNEDP1kqpTmoT5F6676m8OlOcVzju
GEjSo8CC+2pu4GHKKJJTb/qj8gkMOfNVnN+6m9n0KYyTcQxODUEMT50CYnHgscH5
UBXgkdXJDmhzD6OBj1pN/Ro9/qromtOyemzFlpcFQKIl8mll5MhfYAgldxR2xGz+
01SlYLdZ9dJH2CN5jdxi0oPdFEuy4DMC7Ze68jFlzS/UffySYJ/1wdwvyojtrvRx
otafwF8B+ws8bXWSozCZ6PR/MNKkCYmTpFdbSbb+sqARnkZH9eUSXIw/DNjFBtiW
3inLasiBpIEcK5+F7YsooAdmFJEwFyh1U2uIVtUDr6hyltqlZP1JHgjT5c0zroJ1
2KH+OBtFKZyMDWQ5uEvEhVio98A1QSPFBU3E3oI6lwiscfy/sPcmVwRgNbMfjfko
rrKKSn29PXPJISk/2gfvzSzX9BqCEBVKRkv2aRNKEYXxbaIMQrQ7WXXCtouXsPZN
eYICumqIEaa2Oeaf4DQ3qiNMt2kp3pa5ya7ooiQLf+KEiKMU3cimxMoT/Y7F4cGJ
irHV4RvLFmg6gNyrwTM8y196S8NvdRml9k24+7fI5yh1OFHA0v3IeIgvf2CwmadR
K18veDRySUdsGJtVV/9tos6q1kd/GVL5ox8NV97W0VANiQeoxgs6udf9ayEaKlkP
VTHoo9LT6GWBl+ntYejWgdIrZJv/lHIU694nQBuxv8OcBzr90pdvct7rIEPR53pO
mOa1oyI6lskD2xKfI61CAoWSwvfv5qZSTLaoC1yTpymAXQQHqxRIoePJJXteXq9U
4zBIL8sPOpgfcR+dU8GQ2D7TPy11hxdP1AZceIkzPGvvHPTPVb2/3XmYQOLF5JFh
VxP/i6Q1OqOxsyYBSWELqZV+UI1Ok/1c7iVawdwOGQdL950m5RV+a+WO3rJpzFQj
Sdjd359Y0w0Lk2aTMKs5+rgSKOcMsdWgW7ttweNwT+XXTcvj6RanfJ5zCfB72uqx
bIUWQXTM+4pwuViiInVZ0XiI52cUzN8AcD0ULy7A0HNG4AOp8SO5Mu85+RVve4DP
RQEj1/9VzgrRTPCwbhNqVLBoxFYb216V7b97yyYOAwNbscenoD5o7oTEC/gCeKZL
PIQbvtfTfkHtQJ+uJIG52YgK0FkxgUWDXjTsCw/PBG635JK7ILey+uhBCcivdor4
wwLhCPqiikuv1CbBldWIWJoZvBf095G03bflLsgD1PachRQaBkvJ6pkFyzCUnYtg
djlcctR+Ks6dKBIXrwgwnXyme7qur78g52r9rAnxP8H3Vu9GaHWY99e8GI5KZhBa
YK5Vfn+6WIZ7VIiBt1wxdVAsILovE5iLFsYxK9UYSNXiF5QJP677LMpNt6X2xVR+
NgSv+FHGfg9e3cdqn3DptvNIrQWPfAxYLOBxB0R2xX2F5ZIWVm4yy6eUUujccdQn
WOTKJFvhwAUK47F941cIN/TgU14DSdGC1M2aDQSvMOEGcKHokCW9MGKZn8vC7lkX
eq8UxdkD/AU9KtuDs3LW/Hi/CQfiAq5+WtN7B6QBaDydNg1WhwNQT0pXWhCCNpJh
gpFSJe1fRl4HvkJSY69uinbZN76n0RegLRlCoAvd3lwDWn2kK5iaiIl5ofugV/4R
9qN72SYJyIa/1D8ntL/yTso59Mviw3nVhksTxZtBmQZBKuN8nzxvmcC59eDcOF+T
9qbCTswZbcdSJFuD/IflXMWfLrvSN9/WGyfjdEk68SsX35rPbMH7Rmo00RALwMqB
qMA1ag3fH+vNUVsvM+01o0eGb9jOzWGVjAAOxu4u97Ey39PPBA+mZ2GGIQv+IvDe
eSXpPX/mwrVC9Fo7rHGkcg5wobQKpZ4Oce5yZizlP5WGv9JIEfksVLTNSUu7W5il
nskWxbhqY17QK0b3ky5EFOAD7iMUDLz8EdEs6ts4TaTO6SiU2mjQNdSGa53/AaTo
6OFANbLHUlO2NREMPYivIiRkmn1400jOAYnZUgjeWNvkZjHS//hGnmMJ/k2MPSTv
18lWgIKQuePk21EIDx0ryLrNi6G+9/6VF3+6DVwPWhEkCdJbYI+qn5alJhwBuRh6
+Yg/Ex0tv0dhV04ORauf1UoeLy4x2Hn3+jeLS/2O5ihcaZcad3FMYjwfpfdbA4cR
nx6iUcgzkD5MOkcgukgxeKwhXQlNnYaVY8rekd6ILJ8qhfRINsL6DYWxcID7cDI4
W5RFYaiyaTYXqhVANGSBDb4RDZQZBzuP0rY8wLCEmXrJE2V+BbmJ0BotVYA1BHsj
HpYG2Mk0xvNyi05BFSGgFs4JWvAj2K4RVH0mPJg0jKzggdEFgrPjVpTGc1cbt/qs
UB0iQQg/6QYV9mzySu6I2mVarIRrWuR2tk4T75/0kxkzBR/4OX9v9hokxVOYuJAm
uqnLJa96cJuqhp+GAPBV0q2O2UjOKPZfCmRqiexR44My124tzX6VD9F/4a7EOxur
gUTkfX7InU07tzxe/EmLUHRaCWwEgez/IRdP2YCarkrJVRiX+gFJAwKM4Ga4zwzC
5Op54iVD+sJStHoi3i3PZd9hbiR7ZPCsCpbRPuL3gpPitRQTpGE7AWepT2DNJa6V
4o9Eq5dTjkLzOBOU6pgEDMxtHZV+oWzdM7a1mvVQxP8EPrxJ39BG+qHvL+cJQvar
4lCwgYKHvdv2buJIKTikmuXiyam7YUuFmS+Ne2jZflp2g3/KW/C3WKbjTrqfZ7vX
oTDxLISvDauKALAc3oCiHxikYOcop+Xfhd0NU3ryUZBdN0XcOV5CoR6sDSyvaBMY
W/S7Qpxb0zakLS0W6434vHqEssrAIH/3c9JhtUfkEL0m7euSIVe2oXZ4AiSjUtn/
AlB8ChSKuGKBZjqSMT+X3VsWpvTM3K1DZEd44nfYuo+3vrgsJ0se6HULRMIe8af0
yzIQmq6FhD5E1dP06CprlTsY5M8AYJ7mSdavLwRifvzJMPml2LE8VcEJe5vzuORK
wywS+gAnD7vXxYBpPrv1+BlOkJ0ToyI9/a2mXOfUDBqboCSNkBoUYAcRIHTR7HO9
22BRQqllv8liSTEg1HuNibZm0A33OANzQh+mPFCvOdj8oA+dsnWXuqH/wNbPO9yr
nD/yqwt5lcciogokJGyPtFjbzKYslgYJOHC6O4ZgCiSz5TVp5KGUz16oQjxbYMMC
RH2YlOeDzuZcgZRU4jbFfizIYlWWlkd4fcv8KvjKF//VEU1h8rC9mO4sqSZyEjld
z3kbJ5rHQq14l0I/DTjSzZWlA76ggngFXSNO4dHiVYdmM2B379HlA3bKPSbewLeL
CcllVjoeG64QSePQlwpzuJW6m6eKLz8cbTekPLUCH9Xe4CUj9IAu7jBV0UUmGjiB
2Qle+EMPWLl/xA4qZMktNg/tRvdAa4xcrnuKpukByhb/BfDyojF3QomT8WOFrB35
RnVMMOxNKNexhFuZVDOQNav9fB867i3BlYIaXkVcfNQzpsyLcHhwU08vIj6m89/2
8vnu+TrgcjCgD4Z+r7jrta5wBq+LIuvRFB08IIfeo61TGdVoHVKIN/7UKWk85mQG
xgzGi0K2d+oKyzfszoW5lNVA2HJ3grIBldbFBlOM6pRktBO2Fnr+hUmwBbrDSHBh
xH4VOHc2B7GhA6xLrFbsCS6VHIUFxzQc2uCo9RrOTbapHrKm0f08OWQ+F/0XKp8Z
0P3Ml8AxqSEApFvxEMD6OYL5k3KyyrmDiY9zrRzOWrQ3C0l1jyLhZ7Sw3y8svlfO
jFupN7eh/8Wv0r9VORMw79OizjlCFhLLy+BnSkay7BZU1tEUuT0LIQCApljqVnBl
O3IPvwldZXdHubodkQvedPotJdMgNKeUmwcFb5acaC0uGyFpylJb/h3mofeWZ2sj
b8J/JqCDFpwVa0Le5wzZdjd6nTv1ZIDYuiOMQrVtA9yzNgvLlCm7rTpXwrt+ZP9U
grwMMurFAkjkNjnijLQUNYeZEfTXfkKj4rHapk10iqKQxgqs+yCLhaok6bHLGK7I
U9mwhiaiBN41XmCukV+FxC3zwv44n37L45YWczfrzShvBVq7cSBJe8ZzOdHt3R4z
4AGwC/c78lAwLzCs30APiDi65A4V+lf7/Dak06mPyp/9NvzjZOkAWSHr6IV3xifU
m0JUDrNh5N9SbAzOV1Vkdc+bV/frMfjlSGZF06LKCsc+6wDkFG2nxYqD9OjvaPRl
CHUTH19btVpLGAdVewWLqt5OMakYOD/SJeF9zM9zvscWlFzxcsJZUX4lf6hky1hl
on0sMnH4IOrNmujTztDdzo1NpnYFKIUwSf5YV0w+CETLBKA8lM+YGlErSCZ31rfa
8/W+M0gN8JVuvpBsr7OoHtex3HtEFTF/caXhBJxXcq1DWM7Z4220JO0Iyig6IaYz
g+W2MMbzBZS78YSxVTUywKqPvx9U1pyGmLXmMsj3Y6G1WPtFLPsqaHPNRCtnzAVX
ONJrBStP+OWxuCDdNhEgWys3tzvDu6WkRHpYfYOI7wTOGywz8NzEYuGXHm90jRLK
BbWMIQfxBY2mtA1Acwmn7CbBoU1pr3Hupi1v2ip3ymH8iifKI2IhjbxLlcggK3o4
0TTqO5lu22B5rBIjAsiRV5FSq5+SyzcTLYiPhp2wyqVaCXfBGGmc8/Pf0+A7mjGg
Xs1UtCDZ2y4mHDvE4ZiFUDW8pSP4OOInbpjVjL4eUlRA8KgU7BNf2f0Q7DrZoP5+
AKxIF8aXBLuXoxRLhC/rcxyvxXh2NkBGqdPjY0eb9mNX3CvSIyVSpaxbh6KC6EgK
/VuyLB573Pi4TqF/QnLqygf+JlPv7z2qOWCCNyCioEq742v4ffpbVtwcYTrlrhxz
ChDmKEvX3GWkypW3KbJGCwE253bVmZNCHGlcpVvN6nQZFnBS4LZMm7pFiR1wGqMD
AEGVisl8g9eSvX4ZACpewmLucdk+Mkkm0QZkgoa6jsvtPnLZ8z6+KqFkAV+FjXqw
CZCwk7CcVDmgSixjNjZrIOokhYNWAOLY4nAPUbXodWcaiQjrFDLFsfbS5wMHauAS
/zOg9qbgpMUZQVKez9hIi3e/+do+ITnXtzgX/WKyUoaRLbqgIIuV6plpR2IKiGro
UqgwOoUTpGI1AMhDmazBjRZbKM0UBWtWdK0HlatWCkiTVQxG9GOC33WLL5nAUtw0
xS0HTLUL4ZEgFawaUDbHDKA7evUOkqQqaPIZGqYPap2dVDXuAP2QK4Kq5MeLDP4c
Wuk1Hi0DiLzU0tINLWJtziuHxqjzYPrk9y6K8UdrsOSami4V1trWUEIXjKIUHbyQ
QgK4QP8qG1avngRqsFwNunIBEt+UcOZTw718HGwtbttA6DPwaUE/FEnZbM4SaQ/U
cBsTkBPjQjH0Hihh6K7mIvEbDW6OfzMB/qkebEAPTrqQV9mcXOXAaSCc5N3EFDnf
QbPReqZbkVZSsrlBvXiFl7EnapjMTCArMXBFeeRZ9PqHAJaRO+1CPuluudn0sZYf
QCbfm1QsMqrTU8EN2T8P0aCOMjuTlRB68Kbc2VKVUKgjKqgMj9Sfd/3Lvy9JoxPd
OCVkpmESeyIED5zc9RSABBZQLhGMxKsplsGBVYb4eNkd/tGtcW4yzNG6JAhSsiIa
AOUTvDfNmLIT3XCGMAOCQp9E/lHBn2+ozAfFQ/JjinET9jsp3zZ2ExtB6ZeQqFXH
6T9Xr4GmyMcCyXz8/BcauwgBTnWwyeoRug2/1T9W3LVSKYOKjF2hk3Xaz2srclDS
Kg7WfDlsOkbE+MureB4U7/HC3l7Wv5fV9HcPK0YjQ1jAqGQeud/K43xEtaMgSHVt
c7ELJuJkN5lmqw7UT9pqWmLoplcz3ccgSX1zB4CmKGuwke8cX/91gfmC/Uj5yezi
9V3VVoZ7drG2/CsUwWqiPWNSe6A7/OnlVw8U1tjBp495/2y9jn3VgoUxbljM+W1l
6H5ZHwQjAq/kW4uxgoJLQ3k84jqq6FWavnszf5aDBMciY5xtkPVgyrTSEglaXEgi
KvN5Zf6ZcTjm+Vj2k219D6IBkbq8c1SX6y0MMC7zmqbs/z/jANgdtiEYJJb1Ylqg
H9avS/26EYRHlleqwQZ/HVvVn6af5PJM/sCW1mNuHL3nru/xtg2yer9bpe1KMnFZ
3s7aTI84jA9FimoYgzI1yHUajKYYLk2TOqBU4AZfrCvguKaP++QhOQAOFL7QkMKg
u+hIuus0oYRTn+o0WtKnzka2yZzouK8S2wD/hhp0omlh4c6rD4tkh9lXdO41aLk9
H6tb6RTQHBI2wD7OAAf7Y8YYRzwYaxSVjzTzvvPHQ+i3PkaMnF1U0FtGr4XhK0m2
HdvEdr07OpIG+nEVBpegfuu0wBGbYMIOgVulRKMQ/pQ49Y7E60JSQZ0NCQ6lus1l
+Xwvia/eufmY8cNlSf93NV3cBn7V/uJaVwldVNDuByd+V+sDNhHUdWQSkHk7m0oY
gDkR0YclTfBN5AwW6WwMhKle/QzL2F8hRiAr+4vNSpwGZZf3zTuiPy+P9Ip3HCjj
71g946KhCJcEbjMjLpkNSvxApUbCo2J2U48V3aYxm3yKa1iVHaBtsdxahL8lblPJ
uNBSr/Omk17fS8L/p5lUwZchtQggQXej9IRUK8x63s6UtslcLg8Aq22WVsrzMmC6
hbvYi7PIagq9HQwBsiUasOnDA00uyUmiVIFjOsj22RN0yKZNWe4s1W+sADYh2SQW
HTHXJ/5ZB+c4EoLkhd8RdwgGUKVL00f+mbc4vs74ujOFCkZZMU7p7RmMz8XdFh9w
ajDUtdDBAkZt6B0igUqKiVw4EDAxacP22RoNxejy8CZoqS9sT7FPBd6teskkfFAc
jklJcriTjk4No9c2leJhaxZiRuiWo42KvKPRLF0JsWKcVwcbahRfvxNAhDzkN188
/PRw6MwwEY8xrCHooo154oY4bnyXGMVrKRToI52O2x2ggT1WHzzjWqDkHo1cIfFU
B5G4nENpe7bXzDW/41NNEyS2W+fGmLBv6CdgFKA1IplV7wcEg8+BZJyhKkJLlJrk
WCG8Q66Fi+tQvw3FCo1GSIR5lDu56xcMqdUc4jUD2LWcEYqK4zvbX9Q+94i2AaFm
qKsf+jIuLT5mAi85jacSHUzIex7j5cJZAepU2nCEZjWVHekBfsRQl/agSOGoYjg3
WnFS6nTcUTZ9/fPi0FEICLz+Xhu6W44m22woNqwKMjXDEz8NqP/JCQZyt4ClNTMv
bod/wv9NxuDGAU23M3GDo39bFIslZMXpjLQp7ctLIeGRGSMAWfDcul1zjZzhHQAo
6n8DtxHgMJO7qSDHR1jdy2a0N7aLP9QrLGqiObMKkINAOnEJSFfxXdXfU1QFX637
GtGb+auZ79cIJv+pfc7Phw0jg9UBZCdAWZkbma8wUgpKduBVRJ/K2OwQTYYUrvxw
r99956/rkPJ4aEmI/pqbC2UR+/jD7aoK0fmGqj9P61DIhMzv5g2CUU4LuqBIu+hS
cg1lohfR/WLOmZmQ2jPrLfBBUse0VCTZR9SFC0VrAYofltA/3l9TY+AdYCYrkqXJ
Pv724gFXvkEGFWKvPZzw+hEAua3etAL6Ki3aCPwtaHw9NVtKWO7KlDGcbQphd+eL
HDzj9BJ8gdpI25HdQguIGEtBfaPcSxgxVVHtdhx7i/qSs63zHGDPOhobSUc3WZfp
gNFqZqe2B+UlEIpBhNJiR/8CIMv4i36m8T/XchJYO6kqSUE/ZfWKuUsxVMZ6lh1+
hvIaHrdbIWLayiMpc7kIhy5Fp6q5N+N3dyJyJJMVG2aapLus0UER49SASBD3hwG0
6v5zRKcoHP/XS6+WanImwE20NCkQW6+IW2bUIXluGlt1GpvLIRfEWPpDmSL5EbMJ
4YuBBeI5+BAUyl+2obKSflK5LicB1HzWErWgQrDpIl7syHgaZHB+LyOEEt+Qy97w
NtKoeYic/LuX++k0BYG/vHDZQoCon/IsdMABN+hrUhewRGqBrOhVx9pZgI7C+dbP
4FJP6Iym3D+BbnQt2p7cPwdHgQTe39NGLBEzl6UGhkl9PBMNGc8fmDAiy3n9StBj
N+fVNOT1492dUrdrFZdhXonlLpjNAez/X5JzN1ZzXsJgyIbnFHY0cg7QYmKQyOjJ
vRxwn7P+vn8JaZSDcq8yUOqPcR1PklzpXO8LKj35anaikHdMwC1OwI793h5NDHEX
NiON5lsDS7wBmXIWdkO2IDMqC/7XLN1hQBvwcmDPAGSRxd8OYS7NnHm/sgpKjmbW
/+fCdCsYwKbmoURt3aGjQeTEAROmVG/6QvDhWeT9JtxjBL5EDAWWzrFSqMtqYEB+
4QIuetw2LWk5mmu3udyIUHOx+AV1hXw5yRkRuf37K9+IiVQM3qaRIeSRXp+qyG5m
x4qY7Wp1Qx7vBfvv2RSlirq7muNUveOFWT/p6VDvFbKM4oad/w9FgxID5anJ6ema
CgLY0sOWxv1ZPAVMCu4NqBGDmzg+KLve7xfwPWyH31Gd9uH/ZaNJkuCwZdnBoVu2
Zvhch/PrwEcfat2/fuprjGxjsO74/esCf7nAiyz8Sevm0uHpD1pAkeSAJZBFOOlr
o36YYF8HfeqDqNoi5qCKtW6ZeHXKwCJ/5wOifWr0h3TwAg1ziLOP8Aet/DLpEviq
/DTKybKlzR676jW9MkoRmwtdV87l6hMlpr8NOr3oKQitk/+ruL1FZYogbX/hgDI5
8u7spdqzkZNIKwKH0QK2+aivHOttYqiGUNMkEhZuq+px2Whk82Y9G0zVvRBYk7QH
QNZMruL2VAJBXiU/Vk6NPRiqKK3NgilK5LUSEWszLppf9wsJb9zt4+9JafcunAIM
dYa9OeyigroGTMUMCZfePbYqcSjJEWjNSg9HL3XxWTDLsFZh0YmBy9D/vV8CW3mR
J0Bf2UdGy14OB7b0jH+c3HMVnjI8/dt5/6gHylmqyaOHXcrItH2bIInZafV+c59Q
RL8LUEr+FkmDC9rPOZim6qezDegSIY9vCVdxKsKgJKlgKKjhhfZSrQWFqbBgR0Mp
rZCTQd9Yh4VZJMlDCqrhhP3Cn49ntUqT4mhurQw3nmGdFv9MxIDUE1bLKLQLItuf
//Ehhyk/UPUL/6iHeV+TtJdDppB1PwBTYhzY6lEHGO8/quOQUHYY9GCLtjGLqK36
ZFlnm8XoPGbN/Mkt0me5tE9uKMfmZhesMjgG6oIk/Vgd0bQe9dUE6Gx94K7bAU2/
UE8in/GlFGoP/6IaZdsjGv6p34iD7mKaHIuY+sNL27LgdPCJ5cTRIdnfAiu3v93f
bLHP266pdp4Bl/3W1cVdhcixI1pTaC25A1dbUeKZR7DlxxQGvN+P3bVwdhvM6EBO
ZE4bma7j05OCve2Lnm8aLbcJy2He2x+jd7uVX1BSkhd3mjAR5ME9cyvvnGnHTPbK
zTJAIFzY2CxIX8/rISFV0h0iQQsaZggAZY29C5rx/D44iZNP4QYHPGxpy1QR4Im9
vW2XMsc2RUrHIpVBQW52VQYL1FsCCzDWyobsg5y0VYPglv5c+0goXf/1wnfZrAl0
gWt6tKv2HOyoKD8Y7hqza7GLi3JIOYoW8+o33g2whdW190Th1tpDoKYEWmt5GMnP
rkdvE2wS7K2nPRuSL/FKqf5xcBjhbZ/7Gh0Wt5Z2QOtqA60hL8gI2Uai0OiXnEsJ
bCGbWiWKBw/LiYAhRm5Gy+yEyvaOQai1zfKLVw87JmORCOwZgK1RMGhKclX60RUc
xRXctQvSQzk6IDwYEcEWgOptjEqoV/5RSCCOdlgzxIWZ/JDr6BYM9cmORspxsK1H
ol++4Vod2unLyspoZVwtSE2XlAiT1H968wFfyrTxDcHEI0bYAPTjnJ6QAG+YNQQI
YEzIjeRMGgvGBV9ZywXt2wI2kCDi5F3zhXy7MWXELfwgX8kn7hmM6HCFyAyB2oi/
fmkQ5eETN2ePA/EwN+Q4BY3CQ7X008ibQfSAbxdHPNQGIXXbw+7Jlvk4S0kVv3Vq
61RmnVkXLjv298NET/3Fmt79lIeo9LCYeFicsBSA1m9mffSwcTJo6AkyPhr3el7s
Tmt3fyNoSdModCut/dGNnJGLWjxJZ1ityNPNZn7mHwEzZ7FNqhPB867Ov2heOoIb
vwysEcBLr5ee7xCOcTf+X1cXnC1MdCeyjBzutaoQJJxNjYnCHl78uwNAPdcsGZtX
T3lGZTN7ni2c+DZuNp6ARv95YMNoUe9l9CXkM/cTVCB05mSZUHQ+YAoPicOYAc+Y
Pd4fP2M36m9+XxZbUezopsTeOjlMoacKl8/0sznG2Hs3zZUaFC27p7mHMnJ407HU
DHO8MrgvHMDmdq/5JZaMXV1xEFL9av51n3V0O1u2tI6KugYVcOXuMW1p5+XI5GmR
wjA6ipqNok5svuC6bved/MEuMCV3eeVZeyb7Cf7RvLRBZXlKU0XscytIaZPXGGkZ
cfuN8iyN9Vs6Y9BnpQoM9d2J2EWMDolXSGFlsiF1mDHqr5PqKlQKsiMXsW+2y6aE
m57dd8GGxvuS8SoRb9xReFnweCXCngOKFeyPrDvTNewf8sJLfXCeMLjWvJt1Gleo
HrS/XSJpem7oOA6ZHkgiYZ2X5XeOH8avJ/tSvhU5sfKN7mGEQHIhI4o2RysuZRsn
VAVmarrjx5yI8wCC5LeO9rVM4OtR6MtxVR6lIbIyXaAQzV1aP0h1TXJKn8YFe29C
yf79VuEo/6aDS6I75FuzcVpQG3SK93HxiVGIDYPGGPDYxO/ZsUKRpxHX8Nb+NE+F
WBqGS8IPJzVs7a4triqsQdsngyuP8LpagQre4VL3DZG70BeAaM6IBR1F4HAZEWeG
dFPURGAfAm6q9c1xnlRwzlkFG0O/L+K3FadHHlhck7wtlvcxnZyy6O3PuS/bGZJS
PSeLUGHuqP/v43cbVChnCPK6SCJNL+Krb1mCrR9c4fEyqQeBEOZQTGRF53Q7jyVL
6poS7uyhe3CbXHF8rTG6rHO/6By6W6+A4isDRXlnRrU0TXKnemqWFO1Am6T2ncv1
tIITqhRvCaSWEgq89HmyTSVTOP8ELlJxBCIWdl14vk/yhkR8rG3VnNPCoZeAtqwL
ospxjmJRpWKAsrotBi5UuZ5tgNMmkL4KghcHFk0TPtMDRAaxH6U76k0eFy/M+Jts
XcpVGcvbtD/8T8/KJukT5PbR22HoZy3ZljOyj3dKc0UFSxzmkcQlOrrAXRtgyiVd
RfsWKCc7vwD+N/s2wRnuEWEEuSFMYoXFEedUbcJGqSh81XxnJmZlhyjerquOicWV
nhDDuqtmQTwGU8XsfLkon+Rq2oOsyxshYqav/aY74QPXPyZrDlWkk9Jn2HIlMKcg
hVEe39cuGAayHfvvKa9dQs37gEC2demCQwd9xHiR5RKU3Od5v6zHQFilqvjZCO/t
w5Z492MXbxvBeQVHPMNgGkR7rPlENX2bjHnkE+Jo5R8IDFNppHGqRiTFHSASERmn
T3KTM96XSDLO58YfhJt6cIqO15f6c2wUC19X4pac+a7HkiMsWt1/h5sa2O9ND/Y+
0i9xQwfOUHPdXL2e0S1gaT0IRpOIxgdiPxBtGRmkf547J6hDqhN9At6PQ5uNsXJ4
heksvaVYeITPMrvFA8H/a/xdKUkU5LQ9Bq6dKST/uwJ5mrU8kx7ImxWWUyl+8xX/
4HTTtUktZDJ2mUa0wuw81uaKXY49kji/nXlldMkFU1x1Hb9RM0wxq/bWyxCiomqQ
SG59dcSqkVWLs+c8mgwabZ3m0xUEFBnobi28wUlYi8heJGawADUTmZpJ8/Dvw0/4
XnmrQ80SdBcX4ull8tVA4Q3or3JZJySdJ6ixtr2D0dUh8LVO77O/A5j5qjZCAmsw
HyRYchCXbCytbtZxF/sgg50AkDEmCjw2CDKbXWJm85n/86DYoIHPGIBLjQqUbQFW
D4l9cRlHshDoqT1Z/rkLT1NopH5C32mesQEy3SmiQp3iVtbH1aInCa80JDXzeg2n
h1OHgTW53VqqTJHYEYH9LrXA/VqWl8xDmTIkhCLPc+dbDZnPP3kCTXYPvyhUMlzJ
jNiQf9czr3Kg79HDrK1HWpQ+IZ+AsM24W8z0m//60cj/KUu17xtiFgEtN8XF82fC
TWyo16nEpmP1E9+8rM9TEHSRdPUCjBkDWVFuIzkKfKCgO97FNTeUjim42SaUuG6z
WZtjrMyrKLy5eH4leu/zqWwDxJiE6vRk4l+qpTNF1g4op6mlVX7vKS6kN2X+1Fo2
iF7Fhfnuaci8mweX+QsaPtTI5J/we1mwONEd5Uws4cu2yc7VcbwVjQ6cvezgYWUF
j3SxUlcP+zIqc24GP3SdaVhfiLL/OR36ahR54Qz9lQPicP6RZKBjCiQLyc5g3JLr
ToI+dS6tgmuPpUg4BrNw4vcWJ7B3Sx8UREmeS+DrN3kOyHo5v3PNhMXY38qU8MBI
turAhMGRAhSASsGNGnwGBNyWDxqjl8WikNrhmoVIU/GQtj65bYRLzRr1rkU+mcOH
ogOgj2k2hRv1sexFOIYOf7wFryeWpNmJs8ardQqC2ACKMgAk5BEwBy7rM/KfNCTO
Z+IVoygLEnfVlUmhtxPXFs8vqqPbfLfkHq4SbUsZy7hHWegI+9n2LCWK71PSu+CT
ENvxkZonLx/xaKfMrglDfAACQoM7Dr0+iA/qXCec6kZt1sL0HOPWZ9E2UDlw048t
EZGc9sguRlAY1+1hP7zZDH03zMfqmjirxPVu63HeX2WSslchK2IhC01MTcM1n9iX
hN9xGxoTwpLwstGNiQy8U7CVQ7ID7lqhhxwi5Ww61hUxHu4mYVPm3vp90BBKyZ/m
mNLP5fYXnArL+FQQArEMiIn5lE1t3cOJJ0+6prOHsyHTH8bJ8GRDkmoumkGxqvEF
S7aEDtHQoScjXsh+8WmsYcVcdoWEiyiU4FOLfkm0Lg5STa9OiKS9d7YnQwQguMcu
EO+JvkaRIHY5DXI5euOu42IkFm6OWrWrfw7JckndHWQ3mbTunoDunDqUb53zgJDs
x2sFZp2PpC3ODcb6slMum0qWyf8Mi9Mnt+ntqNJsJ9syBDiF2AaaXYW8FE+9qCeM
XrLgQ8R2kDUdE4cRAhFrQjsZeqHX4o38OXXFofJ4svCSb2AP6sUTK1ThEWw02FPI
B3PqczC8zDosbGsq9vki4MGd7FEzNKCDGvY/P7tOquGV3JbcovTcSCWN8bZyWDYR
ZZ0CnnRucYjEmCSj88vk9dwquviUF8IcTNnU2hmca6RB/B5TwTtbGHQjVVi5Fs4b
43iCsjsGL1iMBhCm614HXi8+naav/8196oU4LfR9is1KskYAncuEXx88qSHmwZ3B
4r+NE9TngWErpWEqmjgFBSWoB8zR7/h5NcTIuUVBKHpgzL30wffEVBMhcIyzeyKD
Js7MEzl2IL87utI/h/RdOYr4we3PcIJP2429Gzx/SDPEFaZpyaz4zarsrVDXWw19
gYWli/M2ctjNIRdj3mF/Q3sbt7TNXztgz/QWbTpZaCtZCPH4GsRbZJ2L7u9PiRSZ
gmXR4HnLwp+gqFjNEfQc4xGqkzQpEfFrzWKABK9ROjGv/XFWE9EzuuUp5wao426z
XIGywM11dUHkn0yS3WeyNALYUhE5f4rQeBfTevQo+sJJF2rbdC+UEPbvgGAYv+8q
bPRYTmADMcfYWyFa/aXLuJsZhE32S1SvHoVJ/BphfDdpSz2Lmug8c+WjZKDgkfLz
u3D+dos1M3dooCg8u+M43Q9wZR13/+w0Z8FXO5cx1jKChAZdABdL1xvfT8WKdLJm
FQZXrOKD149Attp2iYzpmiHEstUbalCs99/w/7lSIJ43pk5Pa2wRdng24WmOuBPh
Qc+W4WP2UDwwGB2kGh+RLS6EBtTkV23bM1fwsS770CFAQUx11ydf+FXwjnJYeYbV
4sLlx2HJlZUzQG4JZbFigu6lk1maAtg20oZycRfOFyjKn2rk+h8uFNuosHC+8QIv
LR4OftPfjia1CeXRKzhj2c4RYxWCLPhblt/RLLOM2U6azxwvJrXweN0RUhqWLFT0
Eu6oHH0Wknz7Wh74I+PoSwvL/sIpdGB6+wNTE5PUhCkluFWYDsUsJ2AJ0fsOGVgS
G47p7Fc1gI6XTktQ4/qbAXkcH7QF99YPboxcSOL6ROeYh3zZLE/RzsBKcydyrxvG
7XcwMVfSR+uIY0Zirz3c5AQGFAopbIaPiwXymIveMbEneDT3T36mFrtEV9fy0vRv
hwfv94GHMCfgj7O8rE02V+avhtf9JbQcgCbRiiLQF3zYJamXMxHQIavHnsOGDoDQ
Gs1HjxpLV6V0bksfcN+kXzOIPxb7AozPjyE8S0qBO4nk8mEs7LyR0KAZfCHtaWsf
CCD4TNWqFVGk6i+WqMazfww1M0xZTSAv0ExxRckrr0hc8Q1mTZ80sa2Qkgr5N/cq
kD4swmUFo9YlcoOwgNb0c/3GFKHuRts0iUqvffXfjChWB0BJkmhn0dKwtB4qG7BH
w+Jjbb2dckv7Ay9LSRan5D6tTm28tvGYndfPwbTElGsNtbB0WSSuHVBFnVjoCFbm
Sg9gN3mshGPsaeNUotMvDWUaq5WOpqQr+qJQXL+IGE85XwMlV0u1NOXFfoLZbsat
HoZZbibjON6hteSCwH1rG9lSFim+5uUnAG/xUEp3eJNv/ZSvgThG3olqgqKcEDgp
x61xTe9IvElfxPQ1pAvEvXWq/Wm/WsjQIZO+Y9VWSgujlypkr9fu43NtUQ4UJd2j
Bo632oP1ppy3viffxLw98Pmcm6umMMx/TKodDnvw6bQX96SKqVGXXp65qJx1fm6g
N9UHnVPQkM/UYyFhucJ5nOVTWzZkl6avkEayDxfKL65sHuQEX9vMluxHJEV5UGbu
EzhafYxXJwGGwBCrUG9+JDPme6p17tM7npENn2TEqZo8YwFoYrROA+kfDPXCHzwa
t6AxdYwfs8Ln5TmD/1dA61rMykmqbDRHsaY2OiY2VcHhhvJHGBN7W7yuTAPgoGhf
7/7sdNkkOiMNnnkinbd1D25gz+Xgoz1uKhbpVae4UOlvDsLK5S2yksbJMXxKa3C2
/MkUk3FQVIK4nktouc+J8YbJEUz8E4zv7SdUmRMmRXN8rHWucPYLWpBJnCGVukma
Sfi/3p3CiAyelsDzFf31BWsMjoWis331t30h6uSAZRUSWzuujjz2GDkUHrNBZsJh
ffnzBIV05Zu2eF9+JkOhi+qIQpEFx3ZWHAsVlIQtN0yqAlPKSMZmE+DDEtV2+nA4
7twNBS9FkS4/maM/GFedorsRB39gJVfjKJdEELj1ADe5BnNC3pi3zHPiPsM7N/eS
7j2bojhDH7HJO5vv4QfjAOvzvGScG0WmShz5orQFjDy7BvArzC2WEr2MjmC7e3Sw
EsIDLhNsIfhOuYO40LMmrRAurTa6JnYjqCkX0nsQajNRaOznjekAtyOn7CzH+YeN
XPEowuy4XMrnpLYyr/1LEiCnSq5xR7ewak6pKpKkx4nQgaZGR7lvyou4/JmPCoGP
SZS+hay2vqByjoC/1HR+IJ/qtUkPwwu5jLJeOE2Z8Jle/ayHG7FPV8IBpKleN5I1
+TWq9otzauSJ0wUObLg0mLU9IRYnPKWBWftPAEjm5oVM76BRJsWdUHE414dbJaRm
EFFrJmrvoJrC3jK8+tyVuTC5Ozj5CTjSjzstdeU/8Jzb3C7B2CQgLg9D8S9TZbRS
ABGxYy6iufs7TqyT9xXCqba3+sh0BqM7L7XcnmyFj/8n6rx0AYC8pAmhUL0v2PPw
2glKeWrXK1sEuDu5LNq5//TfVGDDmX0Pv/pbGzVnkDw4yH473mhVZ4qqZj8ZjaV9
wYuZmz6Y387emTi+pEvZytv/izJOi0VQGYZtDFwXsldYC0lQc7jwnnnIuPhV5YvK
aorFGt7ac/WgShAYPok+HmwjfYsWOlJoxfApizDu7tX6J4+Jj1fNdzFBhl1DV653
PFVzUokf+VlfB7nQUaUkQmzmwTUSao365NHI13PuXxN0WT0ajqQmDO7qPpZraizZ
HB0Dz1KWZgPdG061cTlc5jur5ngO60MJH50d8DHY9p9uK1Xf5E6yOo48+QGTnXrh
JoFnWYe7zIZdkpPVADV7orGPmVZvcml+mfb4rg9F0sbvVupkkKH1VHR2cT5yZyHo
WVE/zhF2oQ0JTxbbCEjdvpTJUMdexGpud7xUClXrUVq25Iravo3oIW//xl5PR8Yq
wM3inNKDREdbTF1r/mU1AMeTMnvFAGmlpieUZ30mZcccZXEQCzoq46GGPcH6XVtG
8oLksN8nWEnWHAIbEHf7+I6Ul2/cCPF6FAyN7VnY8TMt7FHk5GCIejA5R5Oi87A+
SbE7cAPK9SlGc8+tqGP7bO6mNSJy5mFqgMR4JDgphWwR4JvOKZGRFAf8y5UnwsTM
B7TSieGA78jL0JijHDNqhXZasqeigpf0s0L6rXgghyonxl1YMbJGhG3wBy5E9HQf
5X0wPCjMZeiUh8ZrmyBh8RaiQsBhPPlxTfFysNqyg6SEELnSRRa4m4Yz1tV1rI9E
4rwzHO7HQ5hPqcrk97bfmolgo1ZRH3+NexDuZlwcXzzWitkv1pzuHdhZui186brU
Hjj4VP4RannqDu3zclE0J443ZgcDYH2gyf/Vr9fk25VwYtmZz9H2CcHOnO0KIBD4
0fQ2lhtGsRUByPhmeIbU3Dtz+oS+AHDPrP72BDBowHOkYbm9Xk2CGy1TKij5Vq7q
+9uECiufdbZALPYBLHAiIihCux37bERBTNnz6oShyMUa4beMuVOqeNevxs2Mkxi6
7K/h5s4PFWJk1AaYK63UA6fxGLETsHulK6XZVkMdGNPCpZyb5XUE91buoga9iAtu
GMK7yY+pOeoMhykWkelD+iduhZWPkta/j8VC3w23eqMyVwwn2XL6t1QGNfwaxpXw
lLvMqtB+JJiss+PIDfBaHVMwxu/hfGe3jDH1dT1077Gs5x9SJEYDvCDSyVHD7NBn
RuRCju37alcB8lwoSolfl0J8ymEjw2ska8KCSBMCGOsa+LfaPwfZphw2gCBrnmZt
iTn3U0qES1t/ZU+lnKJkNyqZ7hXbKKumZg1pdyus4SLQ6iQBtNhhWLSAJVigd6r2
jeJID0np5NfG+zKVoS3Vj6ktDzOUIhTkqrRn5ZUrK2du4UfozA0gZWZwrJFArGYW
OhtbQfl9U0G6D6Je1zERXHfoyGnqbFkpuIE+nyn7MuuZ38QaHINBar+4/x193tLu
jMv1tA2j8FBOXhe9r+BMwq6hp7xccf3M/MuzzchqlS3hiY6Cx2FOcPaN1OgKXF1j
aplL27VY4OoWTNZ7BGyXwymCFit41utFrdA6TdG0inxWHtvu/8WloQ5vSeI6ZZOY
49UeozVtnS5vYMPjexpSrc4fkf58i7UYHokiQP+pDVWLCrE+Ay6uu/13nPMxrNu1
vrUWvMbwoOGfNDVEK64L7rTAGSd9Jcfn0HBiJudNannPPvjPz1i2FQzuLavr6Caf
o3m3hPfWZwGoNN7NC43Hg2cHWu9o5s9IJ4b1bixiCqVeAT1dMxY6FgSrnNzvba/j
JUv+gn25kb/k8gMkDfYPF7GHlyTStb/BBBG1yCJVursjTqZ8dhAvKxLQPxrOQeCq
FCC+Y/kzX8YoIi5HfER0cT8GKKlluZNxPrKGHF1TuGp4vV2dK2xWnpDtYa/YeegO
jGyeGFopK+W785HxzIVhD+Rc/q0FlZ3W0muzVnVlCkWMGkmRHkHfVxpy7SteRglz
MBLTPwfvGoOMkURCJvtabI6nqXmjss2XQvEyQ8Y4CHxJ50BxdwpJXj2/hkmgGtpg
GlpU9EUJWvOiTKcEeHeffcR/6P24z8G/aAq6OREcGkD3CFk5ZlRrawX7YZG/Ieh2
Om1Di3APS5FUWw7F0WxLsPeDy7YrBqckszVSvM4Hc3UKinNDNkTsTQLRGHi4QDtC
Ct83oGhqPDmDabcheO/qCcUyJh5SixRXLagqgrE2Sc6E7bDe3j8LSRCTZ6k45YPP
vPP8ltZKI3JJ53tJ38TQaZLR+r6YKjrCZc9yeClw9oHAp37AwSzBPoplNyYB+wsk
JX6WkWLQpwYr3PQ1FgOvRlNO+D0Rb7VU5KfT4x2xpGrVPIL/EzXTEpqHhgdwAJUt
MdL1qGAnSZcNQHicrN7b16XIkloTVsA/5Xd7uZyl+yWVSczJUofzUOEwcu2+t6fQ
gp9N8SQaVi4pb8S/qJSEEgcbamB3/h+dY+bdQroTsX5a5jF2Fz9k0mRyd0eZipmq
KeiPdHylVf35HYhnu0/UmNFmgTt4Ab0lB4GjieJC1G9sz2imhzUYZRIJlG6tMoWi
d7snOug9QiAhxYsC8xzmqFbJsA5ghH35Kn6gjT1ZaCgioAYpwjA85onoaOU+HJ+s
YUkXqEHM5FVTxRoB/Cfjh5Yg885leSckUeYYz81YqzGXmi4LyvZgi49u4J70jrnt
Ca8u/tydE5L7aFoJAaK/acZ011jruhhIdjiYSa0sM3+ugnQFg7L8/0RJdyRtaXNd
CmWBJ+r/tXXyVPGO543lSWRNJaM1/oGUt+wvvwgd/aVI4HmqcPz6wAfH/wYR1Q9e
a2bb5e2IVzzNI4VNSBrAmqJaIQKlzIxw0g4se59HR4yhGAy0WiNAYd/45mBqC/C+
tjrK9lSoye+gmfWHLVjA2sEuleq+vV+tigQ83U3oaiL1x218pHPoia93JwR74lEz
TAwYjEOZHbpiAir2rUvkMhv24ZygR/JnPruvM7BsJZjx5M2i3T8ys8uxihKu/zlH
ge7U8d5wylgMl8X/JXgrP/0L2iFcKCy2JTgNslZMDzzzq5b7cVNIZsI5372EGKBc
6n0SqsVT93+rLXnSV8wdx2qAv+EwiK/HVTQFUX+nYYvfHcZGyRJOJY2KQlzEQmx5
6J11/2D1KlHXRMb8/mmDhmWwWrCvgyhSa3TNRmjwpoKNMYwzZRu4WLuW6vTn1N5Q
V9J856pzA/Q7vWRtL5RbjYdPf3xcL4jhVJXy/JO6t+CTZvEEhXMvJvelmG2v6qxh
F+Z6thiKdsH+5E3F12sYgoWN+0BOveFklncW5RLMW+Eb4urLM+h0ZfeQ2p1lJdOM
5Iabxr/fUhqaRIaCekR8Vdcid3X3f5a3uq2VVEgV00IQpA8u6L8kTPix9FNkrGO3
b92kTBy56COVvgfk733lFzpdcdk+7RaL3YwWWnQNJBnVbvdVCLWJmslZHdp+zJeJ
u5gqwwLha4OBSgXLPnfSNBk8y5IE5pW4jDcdT6NlEnSSou5iEVtFUDGQEWF2v1oM
QDzpDMAQWMKcthhlsBQB3XuTkCLyYHk9RderRQXvifeFcqh4UlTakHTzzowCPCZm
CxaOGk+Q7izsMZBHXaRvDc5taLwxDEFecMJgehR9OV0zqbvXq4aamvTypMpSXw2I
RhycpXYlLg7ii/wIAPe+aXFj/VrosOElwhrwnt4+54Ch1j0SRlaN0cRSKJigOpTd
c/qCpPceJihTwhFImPufp/WYViZEdBT0imPG6+VnwW/9zVipSLIR6ma4jRYdHrw0
QZPyHvlYFjtV/bMWWtk/lBEnNQgdkHSzCsFODjH7pYeyzTblBP1i1Aghbsl/fVwf
ajbP0NOc89Qx9VU+wNxwwlB40HDrRSjN0p93Ba0yLZZWO/qh+ViJywMqa93Ir35h
h92Si7lscW2xkXgOO6XLoApjiJUhOZ7rjvKavYdrl9lmDAnnhqZCCroOdzUbh05Y
lBGtEJUoUKE8HkLczg0I/8X9tURYHX418kkW5iOUgOaN3j8Hsg1VKZbDMI+sivIL
VrFT9EF4jbcRvg5vaNXT6FdRtU5dCaFkVrumzGxJw0aD36I5wqAn+jL/nAtUsUXW
EBxWt7vKBfry1EFWFWDhFQ/lQ4j/tbIj/5pCgfPkIDAlMEhBUskSE2R6sbdFOH9Q
VQ/73AzP7D2Ribhk8sSsoZXWo3ZK1qBOgnNtTYBI/JtF/R4PTCar2LW7MXpZDSiW
lN3SARIuYhrriUL/6+t/2sTgWcdhpdD833yu9AWW+N/IoCUlV50MWTySXCTw2crn
q2Q+SPaGLHdOKfl/GG7iI6aCtrMBmxGgYTROSAuhrQB4c4syyBn7FiJD2U3CNC5Q
w1R5mueklhTScQrbgLan90s7me7eYnUY1tvviPXMp+I4lHKhNvyjnetJv0Q6wXgy
GZKgY0wkkl7HtNX9LVeXvyW+jSG9/H2e11RlZcQXdjewcO3xgzCyWccwEXsbiR8/
g80/oafCUaXwQQFU6jWw19s1nWqa3fBhi2HEw0LSxqtghgn83vxQSR3rwhLzeiHW
JUw81yIdkZ4o1DJaiUgOq9XVuQF4TV5kj3pmyTiE35DnhbgWecASwuZSIguL7awM
4yQ+RKpHE8RzmRqAllfieqGkqTnU6G41tOqZjs3kOxiea9VnxZDtfmBsScazRiX9
KzVs8bBrjw6QGgmJGno00cZoTJi3yYD+0Qpa84W/WZDi45L9g7Q3TnKuSbHWACFT
qOLzQ/NvFnlmYaFzxU8r20ThsDWtx2JnXO0hHN5h8gFGyMN0VOa3QHzNYAeicvqM
uSRZJsnXKXpyGVbkfOXZIzqxtBpq72t3fxsf7tbyJLhpU9GGcAwN1x9ibtr7Li0m
8UCshknzZmaTT7gi5lYUvnCiSMQ1VIVOEmhiKKdy0hEiFVlKEHaBX/gxA13Ykq6D
KCUYBSSGcqhwz2Hl6b8nXH9gNdua0gSOvo+hYAwpRtN6U08shhmXCyBsvYQ1PBRH
asu41PYOrA6kv9TeXvKVYVijFNwHY0pt9S0yW9WDPEd4wK1cu7+twpB+Q3DsJa26
p5bkPbjzfDJ1O79RTt8EWZy6lgIXqY7vzbD9i53m3F3kcKVez3FDUzS5iOtRQJZG
XMRTvYqUaNGXK/5Dxs4eBwFmwGekmfrJH5Gm5RZIqANEXs+KQqwjR7ejadAGkTVM
VRdwN227vbvkDu+p+poHKW0vzyuG6giUqjX0o1Q+6EflGBaaHOohBPZfY0QRxluh
yp6C7N1TKJwljvu8PTf9jzknKhNQdrWIg+saop81gsuwTQRDeTyyeOjsfREBIsLe
6oxTDs4wagqIVSup4SyetOt3B7EUw9g9UjWE0RLW0UQtc6C7RzYRq8DE2O1OeXk5
QLW1xXed4ss5BMHjgU6bASuvfyJX2LHRPXrqz2+VwrJA1FSKuhvM3SdY4zKHu63v
ftbBsyL/KV9xu0vfgPQByV5VtVG2IuTJyWTGOGKt+HX980BSQb1pa+gY9/Msq/8N
VPyGaXLHyk5stfYoDWfEwuZZfoX/j917ixiVbbeOKDV81UT6jHLCtuaulbpSvhgd
LSFeeuk1K3FHgSzwHeFqII77FNd/6LI0sSbumVmW8/BBQsR/VM0r5nmaV7lT/6dE
m/Tkz/RGvC9C4XCePQcTeECW2orrjFhjnaToS4PXDKHQf/Wnn7s9sZqPDG808gaJ
IxLbE09ezPREdcBR5FVawtyvIrodgIChi811GmGQeBsYCTaKLGGxZ+GoBAEHUXd1
ZTSBHMpJdRx145vWz0BJ0GdRazpOoH0Ej5jThMhF6lkkHTgywZLBbhaA7DWUSvty
Y2jodCc39UfqWjeze45+6uISMB3mU1fWRrb50G2OKIqHrUbt9D2bQW4/gHD/QT6A
MxqsAkirpHZ+zL8DB8mVMAySXLiWpZdp7Yn8wsggmOHjvK5mxFdXrpsozvp2Xbw0
wcPLgptOHzcMeQfQ1iuCxUCRnxS2mFuFCTKruXsi6LEEFMIrVsNi2EvHq8MHG7yL
EAFp1K6q31ml1fd6nKUWTFqCOMCBHiQ/WuuhuoYnlq7d35z5tHGMBbbblhCG0RP1
vE5hWceMmme1TUD84Sp1EBVQcf0wYzBkd5pvoPwJ1nImCaVaSh8PqCxvnODA4E89
dr9t/jq/O/IyxBXN9OR7oSW8nDvOwSdVSb3Cit11lxGz1LmFLFy0/srCGJ6PoR0D
kBZymkxH9Lb+qRVezXiq0uRd/F4VWWsxsToc9iUTA3eM93PzKwU5ANcNPg4sdaOz
Gt4VefRsXuzv+8j3zJmcldXD3YakABZCyAglr+J9lI8hwapkztEyeKx/v0vaJJnQ
/UDW132IK7xrfKUVOdZKDARBJlmUSFKvJx/yBCv8OXZXA/zFkfMdsWhAbquYtMTC
sGiJvTT40isy6bNBhFyXTw+vZkokukOCl4rG3u13vxru16Jgh9pBxDL4siy+tMgD
pyGg4HJmZLhp87i9sazWPV+okR+uOmRD4tc/F03VQoWUjM7Kgb2L0K3x4oAUlFUz
5BZMV4ndBps/N7GMrLa8awVN+VlDsytRPcEc8BAseHNUK2PEb0gVw3kanfqt/43V
V/aloa2YhQtxVMb1rKPx+9lRcbM8Nux3g+J1EwwBwdTvL6Lx59TaF72usyAhS86F
SnDYFOapfuLoS3x9PeZUh/A/nxyqVSR5BHDGBYfBHhZW2fTbhADuezxy/nH7J9C9
ivmMUaZZ0QkWGScwKdJg5BPRtfDkGmwIwBJgKwl0P/uy4sOTENvI8j7ppQsq+8Q4
u6fOGo6G7N2txdle4ML0BC43XfQvaj36ZHoS9wEbDDr3YdgPUH/OiqR9rOrWezaP
Ssq6k+37K41BnvD1R2A5MyxKkcoQ23xW9MK7Fg4hp8jCH7Y8tjDpUsHS883QgarD
khC7PErL5qw8fV0IqH/yj+WqMwg5cy4AcH6oSTBH+Nkaj02IL7SRGbXKchgK/Dc3
b9ULS4sxecwo2dX1s/YBXcJwS5XTvZRl0sLXCqu6vKIeb4P2vLTKyBovxJbGsD7P
3rC1dcRM7v9PY/8sW0A/owN+4FLD9NvnwEUO5lLU7ryAB16ORaELXBgyJfpTPv+T
UsWN/y6S+LovJD23AO/tkzZA9lg+mINTNGba1cEjJorgm7FZvYm+utRCP2pQ9sou
3lMVUDuKndZuhsYCvkO7xhJ7WdGMbITelDouwREUKZSwXutqh5rM7eYjeBp6RnOo
hUGnQwjfH4lYFoURlt1mqslkRckVEhmiuqdlFVcVeqD8jIyEqCKaMG8y5d6mmzuk
pmTCWS2sBGA68KWOjtQOrQPrg3EDAc4ttN6uHPRz4qFGf+WrdddYCRZD3KfxNzzR
/4gQ0b75kv6wHx9V/gtxHlv+e7garjZ7i1aHjeDKjorDJhxZWshpIeeBThleWD+V
giMStKIm1EX5YEds/DM08n8/Sbrm3HGQ3bVMwaWcegTrjVKsihc5S8N2YdI2zFrs
CW3DOuP5hlOkRzdMxHSKmNoOocdWbrTt+1DbVqvtreMJz+m6+t8W+LQORksMIgTB
7NTgvnHeQ+oeBZ/377B6TBLnDwuvFOGuGWl7fprTcG6VWbUVo67wF342TEApcllN
U1IhUjDsyDBqf98ZzyYbE9PMYct3/Gw+pQnnxitlKbVBBgGjsUUsR4bxMf3bkxE8
3bvur/oplnO4h0gVC/i/UjxwGLyYUHOjsRbtudVYswGZZsmdKVJitTPwI3Z7LHWm
JMPnu8gGwol+drLbqqZhPUHsSqsdrJB7W37HMGHsmG4zFTPhbt673/UXk4mTjWQ3
RxoLdwbTZNVX8/Q12Cae4vDfMeDMeagMZMhqMflfeGaUtsSmk8UXJb5oo/8ZTuNC
ln2F5WFVovc/QUB84Bczpf7hlkjmtY4g1w3j4fpvUo2LmzbqmvPvNlobJEtedR8Q
jjzs2qsd5xGONiyzGV9h/598cG5SnOQzh7n5Y/hL60WO0AhKskVSAe2uV2TYgSDM
rSp2JknMOiDRYi/ww41T80Qqc+mfHvFguNoPj3VrUj8zfPTaQeRb+4vk4oERujaY
r7rJrnwiJ2EgM2VGd2lcML4W5Bg78zsv521CwnOoouz9Ea8MelQSl8QlIswd2RcV
kXqtSIAjksct8CsRlgaWvRv5XemObbDpNguHJ2yXrdc4TzAF9sJX9PW3IgY35UWT
/n/YaNK7AAfkN6/zgMFnderxvyCw+cN7XAYnYOQusfiu61D0JGpTOzyAIpx6TdJn
XEf/xGPtuyaz3ZfYT0DOdVY8AFTguy+/KXMnoCmZkG85asGeYp8AbrLxYR95POjb
ZwTT/fJ+w+emTyCN98LNjhzuc75fCs4tO2ecApxsMhus8Qx9bEG4KajmoQLpCSrs
unuTRrOD91RuBnio7jgRvD1DBWdvOqvL/mmRkjGFUNUCCoTlPS5hYgcAo0PTCg8S
ODMulHz8rCZW21N7iMTjd2rUBP6soZDDcX4TZ+XSMJC/e/4kRP749nVbJeQn/pmd
wT9XiFnLhpvMz2VFv6n7hRoIL1PhzZiiG1hp73xxxdq+CoGXnRWksiB2MKiiLZ1I
r4mFkAZQlkFPEQ1ERHRrq8IIb1GQ0FK5uwgfOEXf42Lch9aWaqA3aC+hQx5da3ez
7RUDhM1HslvEeydzTKUeVatB/CDXiLtCXWuEVAahtABiSUq1oIqQ325ABjjwFUgV
EsNxDe+8NxqZfTU97FP+CfkTTXrqRAVVtcZGkgiBXRFg4afCoX484QtLFq096Cni
SuRCClNH7EO6Ly0/ZysBqJK8RNRabSESacAAufurSInzXqQEUmuSRns0Ff8EZ1Af
CeyFuoUAbNULqi1yKBov3m9vvsvA6UVlzyvKVf6TJFBWmA5FT9hQ8qyQvwSPEZFf
sPBWmiWg08Br/25GawFMaagmTfI1ThvAzBNqP7n6dVPMiDPnL91tjLh9xWzssN2P
lAxG2BgGX8Jg8QG20+0MmqyvCkzRaDPp2jcmo9fQK3hMV0aj1l1web967PsgLuLL
nxV4ALDF7yPK2EQfBuQ4YvXNvePg08kCsfZuUhGvCecR8DaB7Ut/XmM0S1LxSIxb
A0G2jpOSwNy0Lw/d+IP2MIopatKRthUqaAxJXKuB70kRY2UKq3wcwwmyImgnL25X
SJ0shQIQG4pE1PdDXGu45zsiZVwbeJ9HZnWb6cVRxkJZiaucbQeUs/Nq30G/1fB1
xpi0jabdV05F+9tjnDzmjlPC6zE5pjajjHm3MPKq9kczXrK1IY9uUMSCm012SoW1
2F0exe1PwkKBe0nmTdHA6sCes/MY+lM0x2eAxWle9D/P4YMDUfYmqt8dd14T2qYe
6iIe1Dnn2LmxlFWiXTiex46hA5/QvZeh0ecE2cgUExTieG54cOY2C2Qf0SaiYGj8
PkouBfvQiIUaRLczLYiye54+qwV2n/z6KiW70maVnnpg4/O1HfqT4xPw0M54lCWG
MhjnLviN9z6N3recdYj/vQ92BaSAEJqcgMVQ+gkk7Jlb/BrDIueqFNKakzRaeY/e
dL4sIWvVgV+cx35cpRDzvNlKaM3a/5Fada3O5AhgOvTgSXCtpDiBaCP99PiATTvq
3bHTkfGxWshV8VoF4odAOE61KkAckLW/s+yj/KgTiOT89jS38v048BznXeWPa1kk
wfuFqmHhmbYaLWYu8LuUG8RjWCOy3kOslYnDTUuhRmGSqEGhrz8MDNc5P1hGGlkG
hNUYjKPGAnht1o0E4vvOfFjlNKbUOaGTSMbqiblM4YIpTBctFJoRqRlFLMMaSA0I
9rzJgx8PCqtE5w00k8IUVcuwM9/FQeMS7/IiwztHdcvXO/c5wjNJYbQ4h2qokoUS
eD+jQDnBw057w/wbpVd2cySr9VTmhCxf1N+F0439A1i6oHavwhUXVBZpqk8LBqtT
5ib2CEcua3/5+gGGWlOcFeOjFDMkwzBp+falkdI1dhakcPq/VffUalv+oPRaW7ye
5ipTguClEYIULO2RtfmY6Txf2U6C1eYw+EO9jzfOogSvGma6Jpz3m3Gchx7LWW8o
DYRAoFAmKS6+TRTFked4dsFSEuYl+juIoqPSMBZlVW5ecYWBfP7Iyx7VmmARQmfJ
9DkU4u1pU5NLP4EB4NKOv32ZWffd5b04ASZbm/yeBaVTJbO8N0Lb4O6gkE2MxYiI
QZV8CKDp7NVM6bMlYhiKFU6nfWk4yGJZgQRouq0SHv8NXZJwM8IBg/q1HmT92TyP
3zj6J+jeVPPr5vLnp+3oVJ729OFAsWbFusiwB2F57fPo3cj5xtPN+mjwe15080TD
cDWNuDqVxi/dr4Mpf+W9SD1o1RNTwyvqU5B54HfxLz4ibzKDWhWFdufVS5ssqUm2
RpA6UCnMR9CEf1DO5kmGFin6cXlVwVk1avN7c/Q5T8YtlgbDt0X1um+Jm+R94u4q
L5xnSfhN5vnTUqm3SEWIdChR99nv/vCQyHFki6hFZOnqvatNFeTx/dUoGJvX07S/
Zp2/r/ffedmjArqeBUT5b5QScKgDpaBUW96+6dwMXeaiHpyL5KDOyDbJTAji4K9y
X32ANphqS21kASYpVj6wzAvyYKv7UsXzLiBtyB5bWdb+d4C052w7M1eMfPlgWOyd
vrX+uCF5dfzmQHQNlZTk53ccL0unZxAaKYAMIkvVHmoNee1bg/5CjaDUxxOSBXJp
PKx+zVhAZF3Rqm1TFx6rP1yD8asZjOfDQ3Yi1ImONjylypQwDObI2wRwcCMw3Uhq
3BL7b0CdoDMG8evYHjt+RVL0sV4/C9ap4DWKLe8IwTLKr7RQoJCX+4Zaqp1f+eDb
eLrVdiSxx7VqVCw3/84WPEYPPgdRTj0i4uhdiDGcxvKM/qGtt5TdNBgKt9je+Www
QpiT3OqgK1jGtclfjOWfZ7QQZEKrmgTfC8KOdJv5nxVKudbP/g6RJj3Km35wpoHU
+yL0RcU66TfJvhuc7FzSNdYe7w6D8qc7893ShQYyWP/SnPMQO6HuPTYBwR8A/Yef
4rNH7HTjHrsXUdMZRo6G1DnJqQVjJmt17GZf4cXYdXsD84K24sBbtFOHJ7u0a7TR
ExwxLTDkrIXLJrWOcQsXBHY8X8d1yPVWa3SyvcAYCo+peqJWv7CUAd1u2TJtWHNi
LHQZeM22r+LIoLNSILnEyU2vajPV2sdbw41Cv1r6I93yNrFduCH+JzcJfJ1QFANp
QXhNIJPhdTTGk5pGAWa0qh01I3JhAIZZ963mpU9jwbjRlriA1FRYbUwCOmYxlAky
CqraOLbzso0L1lbFGQqqfTJxxf2cih43rgmNNMA1lcmTEk6GafHN8Bhc3JRme7c5
wzIaYHp9F2jcpujJrcbgKTNDmoeH3gWy3BnwdiUZhGFozfYItXAuq39/XCjY1dt5
kJpK9S8s2di4MRuJWVMgyhKprHcxYUnwikTFOMA+voOwvSP8thttjvzLcxYLAu44
mzIIBFrbUy2phWjyg9bZphCkTQY2bDlnNZ9LaHxfn9nw9viYvvBX0pT8Hr2A/jsN
HbH1+H3o6tXUYXHpfyZCqYWLMXMF5ScUI/IA9RuhwqYaqGOX7JVUCpm7nbvThYYM
UzabkKvXa4bvPnuQ6F8NzCAOELcWRjBhVlGPZdKsyN04vJdq7O5LDb6ZiEr+u+2O
mA6INfcC9Ba4SrL4zBmrP1QZexGygujsbNvJf1834qmGiANmZbrUFGL7YxtWDO9g
Q0MoC9wHxoQYxNnheErfeb1ZJeF74yv81YRK/lL/h5bg1/HF6xFGx6t3QdhuD+Zr
FK4ewQNbZZXwj3RbjO46jdpdU41fTbXSc/7IKsZlOGmbLm6r30vbSUKkmgtFvlFT
vIDkcvhCsKP04TuWv8ghVZLaDHTDRsLZ06fFAENO0VEgf3Ntlu2OYSDwbWp7edzv
AAzTQsm9aLCEDZVWZwg32p+FON/lrtAX3GLqWi3WWDVx0zG5DwwMsFqhCLi6b6rN
wJl9Sy1e+GBMI20DcZFlD3hpJJp3ilBpia3rEjckDUU76b3r8seuiJnNiG9AJQGO
EChWUXEhdnLrNF0C3Cjqm8CGHL9adUzEZKicMUhYCRYDjkquBrpO8Mk3NUqfPlmV
AH3CkQxfHVpf0frGqWOVbNxQR+zRZU1Y6NtQtLYdn0Pbt3fgXhhMVQfkAPvJY75n
9V03ACvvQkCtlcdLsxlRJp8V1s8wOLkI63OAx/r/cMfv1h+ptrjl9lfMYgMsgpjC
b02Gs5Q/21argUF/mlZ5laR3GHyyNsobMD8Bfs3gBGAvNtqD9NB6se8dduNv3vpx
6yyr/f+QN8qruYOq73dXtQVQ9MtltxdnhrnmpMlUpgIhNNp4wYQvepoy0Agz5fD4
3YoWUZA7jEoOGD6QqDzHv2tYjExRZ0CIIKIEH11yrgNnNjVA+7f58IUGH6iN1u5f
eWEs6FbEUlkeIEhklB7cOxkY+zhuQ8GVP7QhdJTpkyC2G2WLSQ9IsLrI5LZPU4mC
KDCoM+N+7BAYNomF97N4OPAioQsVR0k/8gtxE3vrTrmYN5AvC6gor1NcfYqmq/0j
9aZxUMworj4RM5gKqkjGPSl0hiT5Cns4ypBBo5fFetmhgaB0c9pJHY/mwoe/S1ZM
xphNh6oMO+FGAZYx7mnu4RVWm/q6XlaeJMY4w1iFoTxzl3/l/dURZht9ufBS/xDD
zM8h9fsrhFebGyPrb2+KLvMwZgDFqqz7ztd9zwSJTBL+1tHhc89uu06UZNhZWsTG
OwMFFeNKIsVlLRHnpFjlse75PEm6ocqAOPimQ2cH54FfjTAhnPkT3dz/OjRKiBdd
qzgw6QKmdE8YZUfUZaXv4vcUosMyzniMJorC9m7L8o2G3yWKJLnt8YknUrZV6TEM
EKP9JyyGx99+ZjBUPt7wgizB2Anc8oPAxxEXaoYd/no5UfIFKEIgWI7+xMOh+k1T
pMEBygATQiwPXVrDTYQlp8Kj8kZdTy/vypbae/uElUc2F7YFixmkYhsQa/hPpO2g
gC16ukf7Xduwar0dnxpgrv5lucBBL+96C8JaHlTs/pdYo6vhAq+k3R2RaU+QbFMB
w6qdYWp/fCuUXlayD1kHwFQzXs13wYlkE+3/c8jcQoU/BpZ+LAQIeunwPKt8IGJn
PayfnGlBbkEeQGzjj7hDF7VWIpnpvIynMgl+/RmwuxEritqnu21hMRXGZ0bPk8na
L12/goF3a8YSiDl16vrtv9sousOqrXTsWtHN39TWaRnf+JX5LQfqIMGp0if9Pav8
2lkeXq9O0AEUh0+HyCdBquT1/h7lIH1oXAOyUqwnXN62kIK1spm8NZ9MWkxf0bZ2
uNrRiy6OycGdjFBEI6sJNWzFSukLF0ivQTFtn5zLzoWZJwxmECWus8XXENGhQ4Yi
Bl03XLmh8qTIiHigzrc8Pz36dgx8AwKK2w31Ke2Xrz9GMxwQF1zNC08OaIxvZF+o
qWSlwpbDKhUGRVG0omWEi71DgIrU9/B+hGqEC7MkCCrWuSnm67FL18hLaLqT3OG4
Z9JUi0Azv0JM7LMbKT5GFxg9fJUlv7rRvrDUuzLuUraRxh2PPrAY5Y0KPXvztzTQ
pkuRgS/IhnkyIuGcvwgIFealYLir6nZQq7nsBdxL+UG60tJIcsfB675W0uihGTqf
FZe0Eg+hGTp9QL8odKRU9k4RtkRRN5MYBAOyZOq4tdKYE8P831MGV8AJtSNUqf68
7jnH7zdpijOX6H3HozW6HViEOXd8aEX+lYXs3C1iyBft6Qt8HtkDONxlaR+XMj3S
BQoxkVmMni1SzLb8nNz3PmHDqMXUTK4ogxIM4ZHo3iIOX4lLwS6alaJYZVmZW7vu
hoJ8V3v5h4uJLRcb9q9ZFRzQfQPRMuOwz4jplrmPCLj+ieML2PFKETE9zLBubGPh
GjAvaTSHRE9naNGsyqRNi8vRqtStYUnH34/OUuzG6R/V6mWfG1FfNId3JsIcGJ3V
rVzaLiyT9SXHhHufReSu9akGF5VKjcqZWwDI7vGtHCr9gBpXqvrJM/+XczcpXSCY
SeVQE85eXLn/TSxS4ep8PhLeQ5WX1rKr7bGxyxoSypkjZFh1knTbYLyAKe+v0PQ3
BjvD8MxYM8IfupwaJVa/vZ0xv1WNrHmWut9HOwhRAEqAK6B83srOxtobdTVH+RSD
G2QX94Xo253tGvMCB7JrCDPJd8wN/5UfZD52vqrAVrLN3EiFRMkmNJAibqHDZrmv
onZmpMCGwD6jUN0avWrASb6dVx3IEccvYHj5kQLP4yO+vo3nSMcm0ztTqJO1NP6d
R1LbYwVfc6cG9fRmYoUi6YOmqDRHcBmKkymuNVxjGGDf+E5vH0+lv0AGTy0xEnEl
cCx6LtYUt0pR+pEanYVgqZFimdrP9FVITKYOW3F1wKZY0lTMz1/tfvI4qyCtiSSx
TP+egOE9FCMLAhzrxxvIC7AcYE8f9XyJtiy7p1x0X4ZV3B2efJpAUbiD/V6r/zum
2LD9mLLFU+FhCy1GF1RQEs1xews4sldzQ0QDWZPiUmfCXQSto2Lph8flaiSrcqwW
naQSvNkC2qtdJ2Uf00WMZ4NNF1AZSwMuFP+fU5xW1ITlLwUxUgMrfuUW7LMuLaWU
zcz6MP44EATqZKmQ5pcBZg5WBaA8HdQAbqIbLihiLbF1iFd37D8EErhlY4ra0rhw
ihQvH4rRHJSGKgaIRwG+xHjNMPuZLzNB18mcwXdvr0oXgIaHI18DynNaXX/urGZU
GDdBFJv+jY7eE6HHn4NxngJxmIx7psMtFT83a3KNM0NwZGEjQ0hUUN2brePnO7vA
kQpOxnOriNGflhCQ0NxKdExotKAFLfRL3EzAk7MBqb0ZgAeIAcZo2qawLG5LIaXs
+x1ZleDNkaYQOSYwUxRDPUTPkjKBon+FksyPvS49KAgAZMDdro6Q5i4h4Syb51sz
yZREldhI2VCzVmNdfhAztTnTy/QHkhPRDJqH/E57Rv5sSVPlEN4MtIWgJxO/pBTi
/Vh2uPb+4Ve6DWngffCbYistaCq23yd1ndX6r0ASGSs+CAnaVXnWI/2Y6+6F6kKe
GvKrG/qV+XUExD2KJ8099qzV69wyMrr5C/GFVqQR0HjOyMzulHOwodsIXrMh9OLy
vI9jP7HxYp4A0O/7L/0aCYhiRsx172U2zYjwqe6JR8wwDCkEBVDVeZsxHaG2PGfV
yabnkhIvxMbPIEKbIsLZcAaXWLtWRj00DAEwnSKl02H+d/z/JIAsRW7LblU71+2W
E4bSnEQt5xlbz1aC1wQUSDvwwTSKJQt4JD5XOEpkUsxNXdatLctdHsEC/Wtbh4t9
k3nTe9rOJB/a5EBLrvf17eDly/uKMDkLEzpBJ80fgizu0D7PLRLPIgxEJRZeDTLI
n/8rJhzAVlrcSwGZSURa5toIJYS8IiHhNRYxCapv9bHswtYyIh/BngWqORNS/Gkp
8UoWWGh/4ETjh/6UzFNNUD3Pi/5RWbp+nCfWkAdTVfe9Sz6uFJnCfV/on7pr4SHf
WmfJe2C2w1ZL+D3LLk12qF6lgJXDiBlDUI3IcLtGhUe1PvgtW2Ty3RksfnOzRFmY
UzigitJLsBKyOlGeaKRO/slgdfn9gWv6VYeEjvISdAJjXH/mcE3wvE/q/p/NiAN1
W+A1ZEfb+cq6zJazSO3ixr5BBAQ+bN2uS9S4dVN2uFfSeMhW3qRJU3kAzZbA9Lg8
q4+THwVgeIm+sBtTpOlfvvX8d58tMSwNoW44x8WMHVTulyuWMaM6sheIdocYk0MC
ahACXgL0DUn0VDkIIObdO7UXm6YJx1h/+WVD+iCTUQhlFygtgPMp6pFAW9VuGQgk
ozZiZiWTScU7FnehIMSWKUxKCXAwNpGzYuqTIea6Z+9MIxyHvUIlIPCkg27GGZ4i
PY7w0zbPEYr6W5bQDUul9EOCUr/4+XIqTqW0DkLKiLiwaeLlbo3ECdnjuN7MMuFr
w11wx8H0PzR+a9ZuGteSzVpx5qxighZ2aJrGE3YDqvL4O5R7CViNPnLS+EacPqQz
udInv33HFLQ8H/3adYoyylFSVVxOjLwFHVxp4IsUTtaLA8Fk2ln7oP19cjDmFcNp
MC2Z+lsSROMgnMaXM6PdHkOHhu0ZFRmgjnv7tJcDnLRhLM5GdblY454LGnK9srkU
sXPXR4TRXZ+bDsRgYzas/d5ZTOe8AXmLU5ePHN0tB4y6JTUGYF6ZaL0+7paM7HJk
UfEF/cjNuL5NMOXQXYNrcYByJWWyWtWMfEGfqt+rMaBX9NRbpeFU5rVpH4kEq7hd
viDLNHQr5kCaJrn27sUJQxAFu/icxXfLdjbVQlSuSVaez/B5c/7p/4japshUoemj
BTSWaVleWN32SWnzb/s3rlXmFbxaW4vxyZ2ZdI2vNMd94AWQiEuB4J9A9ptsccBP
xMOUOVfunhcPHJVbLR/ORBlaOs7dun2qFwTEgKxQCkekEFt9nggFTj61mezRjDAL
TqKmzM825yXrCBG5vlaSPpoDz/XSMpnRyXsVhWe7fGcw1CrBQDOJIVgIk0svIHI4
hYM9ou/92Nh9H5UuKHfhdqtlrYmMQUuZbCA2Xl9vL3+T/RD6AhqrWgojB/H7bT7D
UnLL6uLyWkl3DfYN2URSmkqVZrtWh7yxaGjZZQjDQbNCUna5A+gwxnpoNAHPHItT
6c3dXxTnT6JL/NkZ3MxZx0+kRaGuBybhyqTa/JJBJwnyan7hrbQ//uspmBNwUKCb
4TWKJx1UfHb7ZlnY1n8vGmSRhlPjfIXonl0/9bUERj19ghT9AQfNyWlkqTpU7V58
E3Z28nkCiwAkxDjcLIp0k944oeRDFfzQ7H+CpxAU6HWwBE74GSCcD2r9ZNJ2ZGR6
y58gRrt9kIzSGQROm2UDQpiDkZPkHcmNTcjGTB27EPIHPlT1blZSFDyS8G4iMXfM
+ka3HVGQU5aSE6pem1RirhBGqMkyMODHO5VsGeJyMEtWey+hIXvpLDw1YtgvGSSM
sphEuGOKqh4hMqXnW+AQJB0qZ7QdGwg+RC7HJu/s/vRuruEORL73aEIFNcFpNQnz
qSP5NtAirzfB/sy3SZG3QqvaJk9DNTU6+h+gCT6AmvCy+9QQXMxUOCvi4vHn2I4E
yOMcIXD0yzhvUu07svTi5oJUeOjNVSl0Bl2n3WmtK/WzRuG4miCi7/gYHoO8eicB
MayyZpB/MHc1PpJ/cjl1B1rHMeCvMKNCLIMGeZK5RfCEVX7VZKE5eKyAxXOoZFQF
WFF3ZqeG01Hl3Wxsbt2uw1dsm6yFKQ5VwxFg2ZD/oS4lFs3v32r93ZsXRhXRUjRV
bFu4bA3SytQ0/HTwWkW8s5pncV1oIEtc2gu6QiLbLxMuy96BPG9iPVSzRTEaFUZH
tmPnqkI7PDlpRVleeCr8HDx6iY7HrWLptjPdVX+KAXSATMPs79tnGnw1OABtaguP
alXyRe+xZQeP5KaLmudEtm5rVRriT+mUn+vgsNCrBfImEzO6dzN6pxve+kcwt4sL
lJjFWDZ7lIoGgXoDyQRO0025RR9+sbms0MMcnjqio9UviVeogYxGJnlj+IH8Ck50
8PM6j8XpRsv6WNg7kgBtszxA1lC/xof0NV8Q1uxVdEH5bS9+FnKa84TAZbuWkKzY
SUitk1tpSwu5I0qzpWxCIOnLbE8Csy8fgoSFPFMFi5y1gBQ3onA9ArS00sCTFMFE
IyJgnWxD3wB73ROmeI+l5BEe0xdI8nV0uByxhTB+4eaOC8NdHZ0nf4wX+PFDwMdX
JGF8cbck5Oo2mvWW7ts7QKE5OPjJOL0wBXlkkuZrgYib5mkfu1HOA/X12sKA4uDt
xSFGCPmJJcOl22xTftuyxW12FV8Z+Q8MgGF9bAf4elnvqG2Dxg1UpkUazpVd++3o
gOqs1IhnyoPyj/6z2t4RK34xSLlYGicurGiXCRHAveOS6qu+mO6Aswq4WlojojXN
KWu5sl4kaliudt7i0rix41lJYZBvYZgAFFBF3VgrUofES8hCnxPEYka2Md14So2G
fEmC1k2Rco+BmGKdOdJZV2Q4rwvPmrqOlaKUY0XjVx4sQMnqbumOxrbyqXIVvQCQ
PUJvUzJ81OxEPESg4A7plFphsrL/dK64vVijfT6MsLyVsZpDLwNbcNTPSjc1bwMd
WETa1kvLggWzP2erjrgtYuVkV7tvScSmvCyqn6TEYw/SSYzmMZ0JwvG4rNhPQIK5
z5fDXD9oUto4j1mBgF6mi/ZfDXJiJxOQiFjB11j3MmveElfw5Ysb+HKxuonS8HO5
dVDc9sUqG1Mo5QuMa8XzBydNUppOauPjMCqPlJn8KNmttm4xizmQPubgEPKUUU0Y
tbowOxjungCJZaASk6K4AkDY0F5qYhubHBi6Ic597CTTA5zNjQ654ucKqPZMXc+A
/FgAZi1S+h58xYWR0vchjkSizbzoUeIPEqhxgIE6D6XSP9bECfWFTH2WRaDPLR4L
woR/5GSEIbVQ5v9JG73IveO06b8F0bza0HN6Bl0VIUnZanzfGXim08Ql2pGP3itR
1d7AkOcvIbIv5Dp35ukDa0RHL/H9tVOT28e7ufFtx1x3QU67P3mdc+QmYtkD1B+v
HmiBni6bdVFFO3NfsYjDAGyR5nJ+ryzcTg13nB/HeksirDChVvKyHreXuo+Rnsjq
ruU90Vd3DtjTZBQZcrnEdRsW5dE2FQaJXpoNuYyZapuf4yJ8Dvu6a38th3ytAT5V
MBafyP4noLnH3s260Z4ltz5yNLBaP2GjaJCqOv88PuEZV1xMYDDwYCF2Qptk02cr
PWttV6q4ss5iHFSeFCkhdqloyPKhK1d0BjUAdWFXYG//csxnFPZSB/YvTpkLt5Qw
a2K5GZF7O0w1iG4cr3dhRLMbWI2Kzub6FazE7K7B38CZoUDcNj+3Uu7lmfN6a5n0
dDIi0lTk0k+Gf6+eg043wx0uses2MIQFiuAEc+4u6QyycexV7X8520JwqNck+jcM
P1sjIEnYfsyoSXxZ9TKdbZFM3894NnvOEKFqUKfIrKDTa325sMt69MJjPHP/ASgr
rV04/e8QYAjHTUtdKN00AjUaTzfYJ/OsFLUY/FlGfyY/i/I5bRNouzFfdUu9yroO
i6ugyAeMcc42tYZTXDtMLt9XyvxV8i+fQ4L4ffMvX/n9uzjxKgi2jBxEm+zpAxtN
rUGZc8GDgz11JoMuMFZuIrEvMKZj5AVNUjTqd31Ijft9v3HWaglvlg/HgL4ZlWkH
4MlFV6bOHNQkw/+VxU/CMTMLCDTYtESh4/GvlrTvR4Qh8ADmXvPmcp/+o/3yudzw
N01tP7ftCsecfGTnLb57x6AMGoA6nnsmF+yQ649akUHAEOaBuKfNdyyWShaY0yr7
dAovslLrt6x0IK9rFmpmTkRxk85OwmKO4bxuViYCMX+gQVsuicFJmh3IpYuaaFiX
5z2IPxI2cKLYyo7Fn1Z/tH6ke+32iaM7ylC4IHIfA1PFuRHecvNYCKSxkWZPXDNd
0f5nHZdLSpJt97yejC5U9xa7Q94fC0XaEM+dwlVgZ6maoSM7Q8yNuka7PoHwf+eY
LICEYr+yhfs3AW+tzf5oldfNEMyScs0dEb9LGz5fCmC7WinTn0bs6Eit5viL0ejy
++BMUToSPAvuU6Bo91gSASYnjqgwph7/romPw4uwVqdZ7uSwlF/bU4jvk/q9Hk83
lSwdYhlTMuzJPknsO64c9w4Lo/pwCQEGalWQH2uGwXmkuxHV7i90pWf2dvLKhV42
PbYNS9DglJNpOOG0feEierv/WbhOD0GpkjbOQ+zM/bzzJtwoT3mG2QG220eeoM+F
pc3dC5CT/ZDV8Frkj0uuaPhvs44tPxGBOZ+ab77PYREy4TcopCLJFW9dLHHBZjqA
UJj+T9XVinMSg+g5dScqgIAhY9aHYeHexmsc4A0SjNnM/WFaUUWpE2RhUshIVXnq
HwAz3/wDObgIoCLa3JbUyaG2vTCWKKY/2gtR8tfHLHvoWCLt+dXZSDif8lWsBUKi
lQroCVrPsLfHJdXp97UqcsZMOLhJwFFshEogdbCGnBbkUmzHF1sqGLixIjFXZMiv
2TN1uWzy9myRZvD1x+CZEmAb4DRLmkoAZY8Ka2YWTjn7xEZ/kyLvybTmWkcQ92Ns
QMDVEob9aEakox3VGmJMPXzDQ0aYSrGru8DCv2+o+kcI20gq+usrqEXZTZYBy1Er
qJRm6Bs31glyBCatO+8Q/FXmi4sIWTsxEMmy3TpbQgN4DVjZm3fpFPdvII7bzqRO
2EHhAsrLque6kR36EqHkHMGqbQB51OTq2HCP09g8dw3JhP5cBtCzLAr55ULDJnQt
B1m3HMGVAE7hA+beLW7C8ibu+8z9fwLgkfH5StkBW+WA+dbS3Hb0alxcs0ny6QSI
3m3rOQFIRSwwr87GfahvlI1rLA11maRx2nZnzKktVkst+eCLDFFkj4N8xAhLGmlM
pbG2nGOrSqKyjakvY1zoZle/I9ho2OxoWvVGsIdZOKX0U/Ecpnf/ottWXahda25R
aOBRw856X4Xjsj6h2a2ARjCDSpcSIg2zghLrkzm9Xbb5U6ocMhvDk+YKcBMBhr0i
6WxqsQ/jPKw+/7YeTl8Vsxw2iuGXYCYXG+KQiDv+1haJhuosnnGevpf5llvOacNu
UfXEf7OmlQhIoBQcIYAa3YxSCmqDgTIvmBFCh0xNYOy/NApyWK/eStRKGTJ64xql
UFK7Jwr2C7BXhby2fkWjwTwdBtZdKF3XpDKtoiTCC8f4vX42bWyb3YOS2D11+/nx
pWldUA2BfThoEEJRLTPiNq/lLvoutermmiuyLleFoe2KjWvDsTF41oLP7Zu155Kc
Vfhi8NxVC2eUjXT0a/wY5TJm9zvq/jirnQQ1skKjGqJtTh48pzVm4PQyay6Vpn1g
N+5TtnQoJUJIqQiTinAFXQkhp3sFRwfHbXIhCdbUQ48FuF3vICXlyP9PMYtDmajO
lKXyr0ewdD0xF34yDFxD0zCQit4Qh4eB1SBY89VIfNzrvbiYsdV+j8ARTicFuAlP
T+AcyzE7vsgikh1EZ6EqCE1IC+dF2dveFNf3W6QpuEnszTIPWmYvPZEOsInBAb1V
kIiMHbj5a2+pIhbZPTUG6rTbrFHG8FLl4C0KdnAQHWF8LUFLipT6ZiDMJc4yjPDJ
tfKRMHACfjx58BX2A878XPDmcZSHa+IgBz6WMYNWsi5Mp19d4tt6fVGmCzAazEMi
EZ7shHt/7le/x+UC7jUHdhhdGoVfZctwjVuQrP6lBcT1IjXxrpgvX9S9xzO19acr
WTFQbZ/i5SJGRrpuBQjKud1GBskaqjwZMQ/jHlt2I09kl6JBQxGGvyhY9l0byTTJ
e8MMe1BzSk50hJG36ymFndlswpLzDqV0WFVvtTuL/YxMYemgVSryM5wCh6xy6riV
6GqNe6lE2yTUxA0+TFAslOIP2KdaAxmdnMf6wIXhRczqsI3owzrpaaQ2kXP+7hZA
P2eGWlQ6bMurvzD7vApTpht+eGiPNuoIv5TtEbHJtSMVoRmF+nFGOgWW+pJk7E9d
3u0xUDisju5f8aFgSjbU8xHJwSU8jLYNldba9IefKlYwQPyMxA4yYySqByBicE+O
PDWDAIIDCvwAsLYcrMWh9dAsIw3f5AL5hU+FMzojsGbQN9kaAqwR3TVGvo4upOFk
H+qyoJiRUU89KRp43ihA85ERZIFxQtqdnIqH1BvZrFID+zrl8MsITTFSXN+d5BX6
7K5H+ZXbDtgCYnwdwEKir7khQEa9y2cRiYTI7uMnpHVJ6ETb5+oWdD9s63ubcvK4
EAb80VTcfDOOMAo/cZfeCutyKvHI+Im0Xqfaul30qT/iSnIxdBv57S1BQXRbXlD5
dpsJ9FyF/dYDJQ8IBoYjHaK+X+bTLxGE41i0KacE6HRMouwv3tUnPaCiM6YRIuHM
6av5+B5O2COIKaXU3c3QFMtKZ2S7EEyp0CQF5XrXDdSgxZBTqOVhEs149IdnSDiy
Mzd6ZSR5E2g9kpis31qGCfx6vW5be/L8HnG2h+vR72TFG1nS1lSmndYlVcanTSYz
WbMwfjfUw+mX5gFf0xHzVvXg/II2gRkjZARifXl6zuYzUDqXWk0OpoEXm5jioMlz
oBKmAd+x0fdMk9lJlEa0VCw5Meg8SF/wrazkC+WvZi5pyzQ1JkYPZ2TXI2vLCLto
cY7VceNpKSfPOGsHnOJw8VS5IVgWth0A+xFFtndKzZiPe9qqmyI2VaOZB56PzPuu
Kv6lgRiFRNrXuh/Fep4jQ3yhbeaQm/M4zLdvsLcInGisrKoP2DFNGqf/jLNF+/vH
0v34VRGTh69JLtu7zGpfwqFoZ3Yc/2EjVXz13rss3+gNdd9NITU0/wSm8wPj6EAp
5ICipSAPMit9TSgFRg8n9gpUFeHuIes7CDAa/yPO5UdJ/jkGCEUL5bnwW7aoZCrM
3eyGsELT8Q8HK9fCv36mCRyV5ApYyLL85dyda+G3I1bqkc/b6ofDLF4edDUSAz8o
tyl291a+XC3lWnHciKIzyPanFDcz9mvBYJAO+GRGJhE5HyIeHQLmhlwuiJ7z4x+J
Vv5MDwsE797gtF53GsLwqspLm5vCdgytJcWz5KtKyA5Dw9gmquSodAkMVlca0Qu9
4RcY/ygg+QUmBywBpTRc98QvZxR9uPs2PTX/Zr+LSd3Or3pabJExxny2hDUCxxf3
S6cqNRTNSjUMzYU+Iv7LMuGcUE3GR7kBr/zDEDiIcbaGLcBjsV5n1okcD+nYrKD3
iX8M5rwRfE44bVIjwBnx+Vxq16gU1addR9OUAuHym+FXrYVQj7O+fx6KVXsgn/cS
rdUbew6Y/ybYTApUfPd4JcrGeIY7/JNIaQVjn4Su30mQl67qemTfKoVG6pgYIUyJ
Ddy3xmqlRJiRuyZQsFD6X+TnFxVA/qB2KHCNNZYaMaZzRpnfH9EIlSKGObFgukeX
8OxiI1qwR5iDoht8UFW74DZXTp0YnnDr4mwzF2PuIHqEzHxd4LZPKftXhvUAe32R
jv9u6jn4TUw1yVx/E6D0ytzyv3gn+CAVJY4mO5roZCbi+2A6oJXqPtiZKd3DZO9E
CIKwW/5wbS834ctOU/94YlGZ+vWjRJYvpJd1SqKA7WU5uHOhB7AwEMdkdiRI4p/y
6UIG9bGEOvpTinRESSa+dW5LyXuazITDWrNVgW7rAQT9diGxNUSSkIGLSKrJ/hXC
DWdbK5F1ipv6izQqTaOZ/GN2ZO8Ql3yy/ElOPEt2R5BY0uOlfCgRn42l4Zv8lBKa
uA8A0Y+8RkYpV1QBN85J/2j72kgl0vZcFZdFDE5q5a2sYpOhlqQuHjiBO+R9Piiu
xbClD0nJvibF9bFKiLlNMp+NQqq5nP7wLrop2ut5b7P/i00LoxZqRgWskmfw2ctE
Jzujl7fbVHoZ5o790HV9kmcPiW/sjC03sLWgJseqdlhrdtsRCSuFwmLgmgZY09Ze
sUnUGMphVdw520SqX48QuzTXCgtvgQ914gUnt9+w4ttIJBPlH7ZQ/b4Iccq7iEhH
9wRy7bDyXnLSSf5YBF4yDAF+tfw78qGDSx/tTO3SWJggcPM/wBxL1o1tUJ1eDroH
aEBgnXJapvFYjQbfPKtaAnAqrEkKBlyFNt4yu9S04+QnEVJHT6oZY58tV01Ok0hj
CMbug4ESIydgIuztsv96EBo3AzFz7wTjjpHfPAvMaCX45GNWnu4xS/D4Zmkmu28d
7cKzpHbGKJLanl8eijZ0/L+3zqQzgQz/cpFZF/BP0gy5sTNzTVWTZLaUF7u1tCSH
UrBzaK9Npscyqvj+oA88zvAXzaqhWFxBOlg01BBP2PikYsfemI0nL3ke+GoBYuBO
2ii/pI0+3OW3wlNYjj72sosuKLm4wA7Io5caEysvi0J195/yKhdIrmHTeQaCXln4
yKAO+2Yo89zgyv57ybUK/tKKU5bmgC20zGZo/zWG9yiirrzqqg81k/GNA/bJdrh7
zQgDsGeTmKGLKelRLuPgVYVpn6dtjkxIV3AVhKOSpfGGiEUpt90tQAQ0oSdCuY0Z
8xtqvVE65TgDVZvrEVTG8CIJq3egpLwjFJTih4R0q+L4AEvSH7Z2lWuiudQxqZlE
HIzwmAudFFkAXpOGJmBvIbEDIcahKwpT3F6WM/Ho4isOOzi/atAtMjFiaMIomybT
35fJrdV3D6v/0ySj7llzlYeLwRwpapoDYeEf9n5P5Pqs978V/bW64OQDQBpifO/n
XWiiSLr6LWYWJR1OB+qjkdW7Qnnm/cqnBvNMyJf3XXb4O/VqxmKhFaHvtEtESkrR
NmZAke/ZXpRTUhtZ9mUNlL/xSNTGxOMYp5huiiCVwWUVySiAvOhaDtYLA1KpvatS
meCFzhZzmpW8MR2pSHKZRXzzvqteTxqGEmOTFcS627URg+2Y4hxkmhzxphypeo85
G66Eti0/RjcQNrP+4/fxsyx3NkNJwoWDXimgEtKM6m9Tt7D726nyAdhEtkhC1V4I
jONDj76V97TjAauQzVcHba210c4JVduc5/Sl4u//gjsVAjKVz5IJj4lONJgK1pa5
4iJDSogniKy07gxTtnvO+g91t1XdrDT0SdXoIcPCVEeEGIR/99OyVbQT5C7Sgga9
HtWDdUz+0ZaVBObq9pDBAl0SnDt02rbHJoBX2yp5eYsOOqFE6SN6yF0OIT0eN6XZ
PRhXpTj4WdfIJ1fLTGxfzh1YlD5i8pPY2Fh2/ffsjGMUXsaYGGagGbwNCuJkoViK
iraIr6CUI6oaLxDixflLJ2hpYLnMDiJqdz3GiHmnu9RnUP/o+ox20YQXW5V+4KxL
SzhZXzS6HWe9nHhP64mZJncPAaUKOO+3W6U1PPAknUH2kF4qmHkZjLnJ8pheQ1+P
c39Um35Sh4eulHmJh3lccnpmG/imDmWZRQwZHDwFwQQCFswDXK+buvxJ9oQ8ZSmM
/cl3dfh3n7N+hSRYwqDLn/6bgjQIENuWpFg/0AXaoU8AXRAp90SjIdHYDi2xkkvX
aBl6DGh70T4DGlIGxmVCWNnnOh/JHRjmg8PVse6wc/QpvulfpZ+sdUdED8sfketn
e+tFMiskDoyb/Eyu6WRdJwKdvBK1Oe9xF6G3EIG75PRbHPMg7RWR3uDd9abpuHCV
I6g4rNZ1Q1g89NKmE2Yf1cwA6qcgQ1sMEdH0aLNZQ2L0vgzdPtipn8hdeUwI0d6O
sBehGqESV5zMxj5ddaxnhb/BDXKtlVRHc3TGrpZEpz/dCaIFg87kdq34pVVAoHjb
z1P/mzkDt8VcTR8QTz8x+cqiSxlNeWAemSyVk92QjwAfvzSVhaY46dOTqmP1EwdD
Aw39iicfWsOmWCqMXObNg2H2WeKnfyKEhxlRNi/nYAxt9IQPcuNnaAk8Hmer8RpK
2XMVN0aEzgTWD8pkAu0bQMzzZ2Ykh6II5QtroFdh46s7eoJ+HSLrD42TlfhC3F2h
K8QyhtfGbbPNTIjwejDUF/yH6hP7S1gSMq8ONyAAPIOAfAU6rFSaE4/m+ePr0RdR
dg3tJVMjJE1ETe+cDshZBCiKmBpAKe7J+uwVz/U8eXAWmJ10Ezko7Bv+VHBWzyMR
85M8lMWmAgQdSkzxwXfqYu3s4G4RRKEL4YscoNJy7wiYve4SkfZChGpYRXDVa7u7
Yn+M26ELXoHAARvwyq4/WKFV1kTpA2NV2rOh2kzu4VWwfkMrpvRdtRKeOfKYsU8l
EzhQfeR5l/hVKCI3NqtCN6ouHaTV/TQNh5iL5BLq+NqR6kn4W6F9yFshj+sXkNii
sjvQO8jidnMCvN/WIWgCVRwYUuLwqabNZgW8KPEuSBBit/VVhf9h+dAlAUbxkZKH
BUpYetaQb/dLhwuiNi6yobW3KgcuURr599dV3SdPOfWFyq5iTjuwM31bON0jNEDy
vF6rjYpbaQPZxQDYa4k5y72mQ6+WnE5fATzWQTrNON1fyyT4+5cIbl6izZ8bYZmf
ca3srw+mMEdKlP5l2OruOymLY2/b9CbPOYTFZ5OU52rfP6tROvkmt/QYveoVRs/F
Q/9SmjOSsq/bT3VQTW8r0C9mCFSLS5fdI7vtB1+2Nx8yAf0/zFkbAUAFWBzbMaSG
kBTI1X8bJ2nLrmYFSIuZSRD9n1xyi90ggNxYepH66v3weYaT4DIGWMIJ1aUsYY1T
jkOPkWVBsRgseefOYaznMrJFfCPLKoQJeNhvFENGz/FFt8mBQ2orwfb+aCxEolet
IjcDd3ZmrDesO28Ls+G3qOWM/nKilGDGZhl+s/trpExXc9E9YUOfXbMrsfseSb4L
5+MS5EzGu0X8mbJCCEgRjM71kMm4JJfU59G1QCoI01W6cVRIHe9VVQox/05SAnRz
tPnTvKkUqP/VgOyqoLdbGTcyMyLKKevmqAIYhtvsTFtZFg27kxIs/ZmqBurM3eT9
lCFsskuoRbGeCR05cyE2c1mXd+utez1tqgWlwseT1BoT+8Jej6PYMBYW8wVP+fBF
buo2GtSX0WBo38cdCg04UPLwGZKAC1NX2f4sjuWGSZm+sWBMkz6WuMKJRr1b/D66
U4ibnnPC/lf/AP7uVkeQ48vupGb+dpjlz602jtf7E7i4qg5U+WMWBM0ryZ2GluVi
ML8x+hjLmNxrfur9tfrtews5bQiIq+0SL+ZhPwR+1alk9+bjuauOBBsGZJcrHqG2
+TwU8pDgOPXSl24y6fcBTztRbbG3ljoG5obahkX+0xh01CIidocSED8qu+9GxHK7
kDK+m6B4iAnTWayxIVB0ddU3xNCwBD1YyFJuaCm67IaLEx8eBH2BSuJRREoGBtXo
aqH2Abc/wsoJQMWO0GCrfXArEHWNJIXGhESOU2oM+VDjLmGlH70BMv/4LTcRCKa7
OBSh6ckt19q8QHFMj8Fbds+GX6O9/KZenyEdCY9sWTtR0VdAGR/NgZGzDwK1iXut
3oOV6GFmiozjohR9GbN7/oSprcqs/o+H0sH0DQ3w2h/J3qqzeSmthKxIedoWx0RY
LmvChxRzTGOGrZA12yRVn1y3jIFgjJb1PJFRPqYKrwZdiLrVcd60S93odqsQkmD2
YQS6EaxqBPKthy66tnRFYj6TPZwpul9/viT3KVKyQDiwncY2j2NTxaJ9fv3yGY9f
XZB8ymCMnuieodUBbIEIGJjXTioEeXFKyhPLxA8oOQVKaZatCmPLX0ilYIEA5d6q
yFIvVZJwm7CWUxvnjSojuqt/W92aMIIW/kiZFt+uCfFhhSB4O1WkhWVxI3Zm9G6q
bay/nPOvlSBz8uuhh5dL6iUp63u40wCt/QkGq6zL6e6rKy6osGrmDYCT2lucZL+a
rEcLQAZU7iP7HXquY5vqAHUgk/Sdm1IQw2S7NU+Qy15wQPoRcwQqF7JwhOitvrjW
R2+wB0vTT+ZPPgcPnQrE/MNDpNHMDBtvwitzNAer3W4nKd1sFKlWVTaNZ3RqYGty
DUdWr+LcwqBs+bO80Xz4joJHjDE6nv6PrMWIyOXAqRy8jqvTuwQSWP2E9dyjhfOb
6sE7pEiSuBqbLGpKmH5dHBl6Mk/SFIcgoP2Jt8FTsmtcplpMWStMbwOYioO4BNEy
LFP07Ec25NfuNZHbTMxE+Q1yMmsMCMKQ4wvGo8tO4vq5gmS/gU+RxFA4MIekRO3i
40HBm/OhzP3mcVMrm0G2WvueOFG6M1lQAlM5kCZg5nPyEMMTJcoKIaEZfwnAz7Eh
0i7p/hpwQJhSPchN+h6kDnO6jK0/Gun9Yi7FNIt6JydFZtzAfbyDkf1gf1SBYdOb
yL7LytLGDAwoYwZjjkaLmDDjALMzCwrOcI0zm+QlLO9zCv5XRT/gQAJ2kTrIcptI
bXcdaDuH5r5kzUgO+s5oaCT/9rFCGfgP7Kb3+uaSOJoUPvuCuJm8+NHaY5b5PKyU
3rtSOV8Gt/VIvg/H97dubK+1oi2kbAbpMumJ6MSlajj3iTv3lyfZr5nD1Gl6GnIV
M0CqbrU4ko63aT7u1qAPya+hCvph1/19GiQ1W0+fE2oiAfzi0Qlb3Q0HNX/Or3JO
U3wx4RJVRvKR2I3Mc15rMhtPnFI54sYiJqCCXdlyJV37Pd+xwu2eT5t5bcg6ipUR
xbqdRfjk2aTK/iQlPoD+DRnf/5QZECs8Fl0EPi4jtErlOEGCEF8w3Jm+N2fUi92p
TaZcbu7ivg2sUvfWAXpuoUt58gJi0xy6LzUFY/8SxpZyoMGJXOXTVtN/I2bg4axo
RSLJlLHP1+VktFV47ZVw8+Hvfk90vhi044fDEE8XgK6PXzZiskV30c+RC7YTMB6s
Bx8HKLqL//t02VJ2cC9/x3VgJ8KSYOIB2NQCs6mVoQIKSpa8gDSd7J3nrXqyuhHC
9oGN5xPo0E39JcsbP6K4cjTcWyWWPgxMF/wGU24FqBH2JVbHN5mYfOnilARfTFtz
Ik8UVLPJU6keG9ta410R3qMw3nm8EY0bUs6VfV2TXZ8gzX00ENdhcrD1rByu2f9C
E1rRlOmfGWG4XvzDHHpfUVLAsTwsil3xogII76stXCUYAPof4yVIYmSkRtHximYZ
a7Xp8XxFxG0KvcQXpEa4TrgLJpbh14igMkCsMNWWHH4Lak9MndNTIXFMyhmDpqTc
RKcwPl7Y3Ja5cGrjmCVxbxHJml/MpnJ12Gqk+L5kR0kv08BHLLUcwEg5yfGn+U5H
mgdSwsDgcSpQ+63Lq9SSc7Q3HJrRS29JhYJZZ4QE/ANfypxnk///0emfMKDrc2P6
0qF13NkjNXg4kYcvldo8R56WyY0G75U7LZzRlJz1r7YI3IKCeFnjfJJNIxPb056Y
BwkFDrOB2u78Fi5jMJclq5cIhI/PeCH8+CiJ/yq4DZuYhjCCI/4kl8HvAKNKhOJh
6qSFc/cTYFBvnnjZBMpdhpGtHWd0unAN2pFY8IcSodbeqtg8cC/M+kVUSz8OLicL
EDJbTQqNmgx4mAmp9VWmhboggwjitrAZIz62UkCHmBYqk8rocZH3y2IuoyzwPM4B
BeGNyx5+NmtNQd9zIPHNkVHeBPpTgzHndzMg0rc+9hOY5++JyCLPOO3qY84+5Uol
ZAJMgYHrteoRlvdL5mM6HXaCmV1suxiN+hq7Q5felSBBiNDt72giO9oicrcV13k5
pL0btI6s23hzSpLs5H6ThLTHJloWK2knMnI3PR1NFe3QMCFrKBK/RlKIUsu/0qCf
keNMema3R/UPCWD96bIuLeS+HWWeQVzOd1Mx/afnGuU4tzPHaw4IOGtFmv/p6X88
DY2KUQAV7OurxlOVzNch0LrkVObWuatIkSKL15dr7obhY9TSCYx+dG6dxPyyvMnu
8YMxGK0/MLltQQ+an6mcAa9mmzeN+kNFZL/deQGILteLiPsPfY4quzsXKqnWBIuI
PWpZ5yYaE9gjY5hvI0kHqEDpcIXYM/mWWHi7leq1WWgdbfEChGWStZf0OciST8QB
m/CORCXvGNs7ToREYpjczoEm72tmDJIkL0l0CHUKcZs9xSp2e/jSxoFELNsPSXZZ
hcu+QrGyO7FQrgEDAHY0w/GdcYYHU/sipmc6YwL+Lr40zyAcGdLRK0R5vN8YFFOD
QMnhi4DV4SkglNgxnflB8pw3GuoTRQugw/MySNK4P3AAA4ubUfDG/q3EtqB/MyyQ
CEjt0RvMuZymOj0oD3lUzVqMz6JXyEBWvD2vB/mlFDzN4IC+w3/7WqrkHdoALpaM
gQjTP6bSnkjjzeWqRViMAD/49K/HmRFuHFyP+A7bZrGFT6r/hp9wzTP6Oxz6lNX9
o3l5BtPgFfrAfbMQrAAo1hfmAM3C7JMO5D0TeqJcqw0IzyCxNRmfzo3iLcP6jvTw
h36S7x2U6ZITyMOwdVxQoHDasg0WHXWU0MxoB8PXbLsO181t3Yk1V0UeCB1i+nNe
B/FAYFJf46B0VfaQ74AcRZjzv/fq5XPpL7jEFND75OKYgT0kVpl0zGaSJ1kxrY+J
uWH8+tthCCiJgx7Otpftuc05yUCBJMlqNim27nGL9xjXxZ2K4BYO1SU1OidfNthc
DeVYXI8wTdAuj23/vNJuzxo98E13tNIJwXcSfje2uLa1+H9lH9zrmF9OSkjmequr
X9PbqkEKNcM/0Wsi8/jPZBn/paUlB9BjUm1Lh3BTdUJz7YgYHhglBRZMKbFYGRLV
IAVtS6YPIcP2pYXvWPggeOZ/Uyv2a/+T9eh2AikdXyt/qm+rl+QCm3Uysx/5v5xU
kfeQ/gJa++HrFtBTGCx3EPFONz5wOTy0Oyw8sdZb7rTIYgs6Ar6mnx0/hHlX9MHv
1dp/v6DFWS1GgBNHc6w0iF3RvHkBxpgMn+ricbRniI1tMZWUEW9NlLaY13Bk6s/P
xTwbTaQvlhvDxQFE+8padK0Lq8Jzlc0UheDjpyo377sfRGWwaqah/qDXSCNfkee6
LWvB+vG3VrY4dsoilsT+QkyibJy0BOqZMSxGOEcfOgfxvUqSA62A81Ok15ORrb6u
qu1/rr+czMctIC6+zPn74TSxtdM3C3OWY+ykknTFL8SLmxMwUh4a3XYh496asdq8
kDnKLeSLn9BUtnVC/Q6aJUmr3KRm2OkDIL50WPv1qw4QJvCjF5jMwkUngzpFDozO
RA5yNNuvKA4UBje5SKfZkgrWqarJO4TYx9E3szZZ968Ok+XZkMUkQ8GkY9ryt8k0
RpJvPTv+FYkpq+5zWa2sJVvK0A6EBMqH7bBguoAuI3WdeFB2HiOnvq+6d6IGYRBt
KQbzsZ3XJSfDK34UIlYSle17fmokmBT8KZRKkNHvkpPQnsZP1W7sq9sm58V9OoO2
GI1eV2JFoi6qUPdv+EnLJaDfAX7s5L4QOXnyTsRJvey9zS1nqglFsLhngmR2K1vU
Gh/1/7blS9VBZ8dRvOLCsToL2UpkOpCAgWmkc1hhcRitCB3ORct7JjHBd56jUeIe
4Z11MfxVbbDIQAP8wf2qb4Mp2VpeoG70QixXz3+D9jKyF8AEqbFhmi8WaY7ccjNd
7maFjMxXy8T0fkt7mA2C3vT7UyXBRJKUN3sLqBehL7lJDc3EOnpFZ4x/YPnhEQKk
DT1iIgnPqLUdl1VGusWXFJscKMcyzwQnRQSdOyDe4EMHVzGi/hGm0kQg42/c1Hsn
18GONR7R/SZclK/MqtgyWWT707pPX5DJ7QZOZFaUTo0x1bP8RHpr/AS7Yl23rDM2
yXLWrj2ngyrSI3oYKgwRNHqODsdatepo0LGBnrtenvJRYjfQdrD8a6dPXFtFVO4J
7Kj3/9bieMB4xnDzoyS1c/yW2xTUYeU32HnUX/BMhi9Rzvwx8HS5wRi3ut0LbAsC
Np0uUKKC6jFZxwoJax4G1w6Y4E9wgIisp/tkSLX3RQZHFdLEMOpZaq2VuLKlxR1O
nUYuJHLqbQnry0kszZq75D3j08MEVuaJ2hVhqqzCjbN8deyryspiFYVXSzhvl61I
hKldx7O9LMxON6yK24foSV7+YY7Ib5fEW+C+8b5nQ+NP5gRAZdskr0DLjcxTfBf7
Ok41gI38kvdPPMvRJicalIEp7jotsmgPzce5Bo7RHIiSyh+1bG6V2akLp4rXDs0Z
yOHwIVP4t1Y8O5G+x9QCpwZSgfXrtdRQ+m4miwQr0q8FLLN8CYMZm+mX3BH8TbNl
hMUbnIMD6DE6DZ9A89yn4b5bOB4t3HmmHhmClKMvYRh/T3j5QAtBeD2kYqRdB/lK
ZyYGHdA5texaU5nf/CVu6CqzX0ri8JexbLSE5g+gDfYDUh8Z1CjHyiBHo2lxDUa+
ntxOeQJ/zkaqOml8FLTwuKWcZhLvEGJ/b+ZHYJnBadantOmAhLmMNTqpqxx6BRuX
oHB+wWnE5CP85Y6n1u46K/BZvog2pOuEB6xajrk5dAB79x7HAaiI5CVFgqRj43w1
Lmoz91n1s86R/ZUaHO7rhsjx/LEM+Qo5PnmVIuSZE1qf0OC9wp//gAAIhAqpTqwJ
HynEiyFV7Np+pVg+j7+Dnv44LcBse5vM1TnbFwjjfTRiWqkSs3GZCfLjwhrr/OVt
7yvQEVqN9ES27iGOuN5p9opDiQf3AbWJFI7WlWY54FslbpX24Ex28IrG+rXNNCIE
c6VgUrVfoEQqgWdCM0mwgNEb5+y4j4EvI0z6pkj8VVE3YTAp3e24P5rfRZaEYGE9
7z1CJkRo7dtcKsbdytcZFEixdsdrUjku30xdPt/NlnZRsOPLyWsHLpYta9gpJjDL
UuHYHHgOZVVzoVi1JTTFr97GwsW0Coc+rKl6UuhHjc1Gz6ko+kbTyVzkblbT67gA
3I94q8wBc3In4FmGt90X4L3+DYpgLBMp4JzdTOtXRnm0c2MIaVBF7TcTIs1Rs7Yc
TDJv2bP9LRZS/QY219vEIfSuAFUbyQr4/1pbon+5oXo8xQuJUn0yG/KUAAlvVtfv
/xqqqomK/eYO8d4qSibW0ZjlihJpl1FCnDkYWO/tARxhJ2DxtYRI18Pc+0m8VimO
igHVAeCAHjzoErIsdqJzQ6sXWwYZ3QEeSyRj2ecx42+s7Pw1L0e2I7WnHsb94mXQ
n+K23ZaP+vcQDg/EHr6aMTQiTJD97wC4ZlJk/rwBqJWyGKhCNaZQoBKV8Xnt11Uu
EhpMIPUL3ZYE2GgtmtdexP5/nGi9oDCxaSUDRWwm59Iqfl7dpAlRrlyu6VQCL89G
JSeHSjFS7p9TDaZYZ2tCjlatnrSw65aIF9lQx11dA08aI1sj+SI2qAC5sF8HlCMa
qIqAV3ZnuH00Z9+5Rx52lr7HU1xJ+izoXxJxV8lhMaRM7g5X3p1xN67RyifynT0a
f5xLp2eoN2hTC6dHK1IzyjlJaAq2ud1OwSc/Ozm+9tIJ6Ys1ZoODKGF0pquj6umW
FEu5bRnV7VcaZ8z8/Gb+xvnnruTWZByOOk7zohNfkRFRlaEXyxXGC2DQi7mUH/uu
P/J7anTCaSwmkcWn0DekH1FxrnSIJhgw9Ml5yhH6EWZqP9IcsXFRNt5/XDwH39O/
QHfjekL61DEKWwbKUJCFlPYgI3Zjn/Om1jX17oUymYKI2RS5mYv8SN9lVNGEjoRS
v3EICmLAQyxO0hWUWvE49c0t2VzA6gPpIQNbPII/m8BLqFBGTWRzi/nOGFXMOj7L
oW/kOvrIxAdEnJTfBBrNOTa+oiZQCOKUV98agW1V7p3oROiGwvnxOfaEIW3ZdFyB
+R4zGXjDFqZTSg4UQBlEugTS2sBV9Dh7d3okT4jBzarBVlN6gM+8odbw4z35JTA3
lYDsHzssUC6QykHiwUyorCrpE0ZCX0e7CYMBr3XKJcqVMJUdpa73Sd9OqcbaU540
Q8/LBQ1Shio6qHYKDqi6oPm8t60zlKK4UGBvZcQs7zl9xR/orjJzkRbIcMg1yzqE
9ZfK0g/70s18AZN2eAhfR9aEjmpjazEPeraJ3YZOgF80LoquZM5lkG2PN7/7jTaY
8zgvVZIU19fTXadUYSrnbfhMyHVBaet7Y38Hv+eFh9OeKUbTu6c3dsqajaWfx1vR
WKW5BI/MCM4QpjsS917xc3jH5BeuQ4qSHfkq8yHdXy0UuhPts9Po/MnGN1CgKDZ3
apYK2Xim59dJlcyVTyEXlmsvWsvjnOAU72OdKr7fM0Ua0Bkhxg9xu4WQR6IJOf8k
3eb4xfS5LpPpDc77VNoQsb4euMdVX9uA2kfuh8Q8v5BsE1m4kZIO6pw5n9sbyjF2
IH6sGj+a/S/0tqklP3jhHF6LhbOpeQNyzwhNXomcKFi0zkH3P8fBlBHpBibQrHp9
mpsiVFGGmRt9UyfrI82PBzWs+cqXammUlMowpLphUAud4Zu2gB1TcRBIUoVDpgbD
wMITX9Tc238xKkJvMBfvdgXyZEai/A+2QengSPHSSxIx4Pjmu+AZJ4MSc8534Esl
ty/xayFzP19TjY7hymcvWKoOK7kVKKal/AHw6uCPBMXnZMZ6DtKDmEE4Gei4pW7k
kG4BSNEULaTZDogn3pqsajJi5pFDyyrIyL+e+zllQpG7SqCt/UURnmzqMd8fXn0G
RyXoiESIdIm/forCAQMpfLLkB+7DWzbLqr6VRylcYKH8u8qbSbTiB1sJmfYuK0Fj
ypcJkECBRw3gXvawV7+xtIuN652awiyMXfO9ZavTGVI7rukhKCZZ9+KzuRWPftWL
YupBDrpLCm8QcjhBR5BTEqYDlQ86IPhTM9zC2fCJXJQgCXqaF8vSPy0+S/IMEUhP
GlN50q9fDdwIUCVpIzM+wFVhQY02LFwAYzdth3CSstbNQhHMVmR5PVNOWYY+CwSl
a0UOkLZ5kDWQQaHxUkg4H5V/FFFJZ56dlpua0jSkm1MReJZtKn6nByb4uiBUBitz
5+Qdk6gVKod0k15UttwK6FVWJ3YqqhJYbnhFW5wmatP1ROY2oVIoUxUQMflz1GVN
mnC0c/sWTZYlRCBFe2vqnIY5hmb50+oKX3Te6MVni0xM0jFpA2MVewymCdFW+qyk
DCAz3IS2VOQDYViOBUqiaSQYIQTkMU1dzJy0yMte2KVkAS0XOAdfddUgW/wS+Avo
iF4vtihLRjTI/Q9uf4HtdsBgDZet1ubng9BKRil83x0shQ317b93aPYy++cRVVKl
3PByjFOtfHXY5O0ySIFX7nJeAYBURCg3HY67vZuWckQ/TdwOfaeLRD0ncnidjJov
GpM0LYRViLYuv8lFJc86IaZ15XYI7hymkhjLvN2mDSAu8m2NKbiQwfzsFb/0M01y
UMZlW6G86xeMlr3k3AJTGCjkuDjUnu9txj7dEmliiAwlIq7k20nLb4GqCO7Fyr+9
4K9Y7m4p6KjprvU+QgowJg3BDE9vMXCA+HeEptXTDas07onx5HUbmEX7ywU0CEt5
VduWYCjOBwPtiItGtrZxlSp5kguwjrPZmo/5vVuh8A7HJPvdbG8huuyZy2oSkGxo
jt2eL8cRECtz7Gl0NZ1DG4lGlAF0mnn0Z+pMW0k23UfpUyFfbNHzqbtfivOLAIU0
wQT1I47uTlQwOdJIsXb7lWZJAXKY5mlWFj2maFxgbr1Awven9xsZcI43/WXrm10i
BBsDXm68y6vRZXXaWhYwcvn8Zr8zkeqaNydgqK7JfPXi9wjOJTTGnWwhq9H4Mirw
yY1tf9BiPMziS9MSCivCzmyxC/18P4NC9uaVMl7CxNWxeB21ibqreCF7OFYp5ujU
eF6LPs7bNXkWZAqtsxlXnsejnDcqu+M+j7SSAEdaXid1rtiADTqRCkCZAxcMhN5O
RpEC6omYjgklae2HOzJ3sfiSu4L2yZ9sLZX2PzRTMV+cCfxJOALbolBc4PgndNNf
5P/C+ueunYLwijcDXXBVReFz27g7EizN90ddRZrkeBVz0k6kh8BlK/HpD56g92QC
ho+4EojuwvmYB3U4Qfw2tTh83WGp5c9+F0kaMTg0gJzfglTUlQ2KtcpGC1DPsqyN
DpcxXu9k8A2eIkEbqdeAVxyFrQ+MU5oq0S1zHToUtXqU+g69ZmPXTzB5t5qKU9nJ
lf7kwQ2/rnobaE8xgHvgRwg1dXb/xyhHylXWmylkkxKzwpCJgvlqmYBgasK1xGuS
+tF1ykHRrYz/tqj03NXv8VovFYOHfV21imZt8ZYjJ4YZLCmHw3gSSqrcD/mAxo+X
WygaY0MhUbJ0H1xwn5kflu573C7F+fnLxUTAWTRxetK1YtsCDX7l8nG/GabxxeDY
crZm5957uszT1K5bj1gbq29TuvVSuvpT+l3e29xZ+upl1lqDQsnef5z4creiy6sg
ThByUnIB6i2giZuV9C12hhg/Erj/H4pTifmVKIIpUmrj/3lw4oHyxxFK+WpBTES3
ffrW8TNq2Kb0Bp34D1gXIlBQCqCaY75HHCJvaNVphEmcNacO/+qLfLqFSH5erPtI
HORTfUit0bO11PAmZ4YTXkAB1OhXIcrNvlyB0xxU2PGo4Sp2EUfipG4vvOStYHH1
Vb/QLRgpkB/OFI53GbSRibVk4jt+Bc9q7yr/Efb/5o+FSdE9J6r5uVrkUE6d+Ni4
963aHGkpzmB/Kqw1OO8sehmKT2yYOMz/fBk0uXeV4B4Ie/sWqa7632UN4WYhUG2q
GNn3W++pgDg+FCjON4anShCiaeOKH2ky3iNb5h5q+2b6kgbYsPYhNIN6AR+CxKRT
3G7Yv03r5H+laegaCupJbW955iAV1t4+wmrMoBwvEKpPOXdysXUPv+4eIchqaY1a
IckZtJNZwfUx9EoBqE1R0bSlStoin9S0+Sj6eAVr546o9mZKzgYGmq4dBsE+ojsP
9ozFeES1ikLk+qbtcYVmZi9OUAUV6dApYyDZSLEUXnygQArlYNsYU94bhGXNJRXl
vH6M81D4lh9rlGLDMKyJcwK+R7dUx5ENUbXhdC9tRnGQ3l+VPQ9KAZf4MpmK5aSb
/5HfF6hs472p6sHLZtJ8Ow2DeQE7ec1zmUHI6Ucv+kf7NEuAgtRPpN+K+8uvUEJV
s/A7F2pnJXThihrDfJW3bs3cRzHADFfhCdKSwTPHB0EdjPenORmAUcT/rttB+IBx
IaCTLv8e71qWl8kR/7+p+SEGtgJ4pEAJdGWBQFLQObx00qsumQd3mToYl0hENJBb
TFkyhdU4g6uQwFiEV1VIEkPACXcPlEo+JyKpuS7kWm2WQtn4i6oNeBO3tbC0WTtP
231jrVXWDFvghtZjpcfRElKwir8OLUndLNBm+oJnuBHvXamTeVrlT+f5VsLb3eDg
px4/cl+8e5k52GYM/rcQyRPHheDLYbBJHIrCPNy3tOvjFAkpeBm4x925lCFNwVd+
4u/15jAFmRLxprK9/6rRWvGhbDKL7HnwNO2NaHsYc+ZRHPFqJwxGsbunjY0bDGE8
kmGL4MgEXVAESrEo935N+GsRsX9iQqvNRRxIs36FfQrzaGjwnctNeJRfjjzip0Ek
VuNFrJoAj8zK5QRdXZR8O2It89F/AKBwbLozxSDJtHzhsAkOXSPagxjgMPYt55V7
P7iNNBD8TwL0m0LG2EmuXzIclPFexmc8sYtB1A1o4ucG4p/E6FcnOy2gFEhhabqD
VguymRf362GeKDX446OYxaGO7p/ZacohnV8pgbHqQQT8ZW6wWnaR1f4s/HKWveHX
qMoDmQKggNcKXIlXw77H0nog/3eOqKm04rigXBgPF4jx4HY6sjYNpEuA/600pzws
a1BXk3y853CCAJglhf3vso48aTiTPpcoEG8RpW1T+GtnkXMKpOXu83iwiufqKyDa
kHu/v49LPsO9XJ6rCTs2IHlNTICSU+MFppwycFP+//SL1MINmwGXJXvosikMmdK3
3QsE/THvVndBjEYE1wXLlzazvOd2vrnhKWkHkUNWpHQTa3CDfNJTR5a5DJKBMjRN
ZD1+SWIKrtvnnr/pSQJrRCbxz/8G1P6bBoPpsoFdyOOrmRRNqk+D4PS+d4teC89M
eXP7PZL9RgKtulXp4g2FR2S8E32nKihP1SXGoLnnLfil5eGEA+GLlFlWSprnyCns
FnN7MK34nfTeZMHunEaFfREE4oOWTjJyc9Eou20nX5Jwt7LYrO9sGCaYrE7cFWpK
gjTUM00MB2jRRjhvF2ttlvqIU/bTO/vXMmGPHVLzzE7gIgP80HGaP5bwonaP8PH7
dmsVZTo2t1FEwWItto6oWjzI1iXyjzSsO1V2xrlx4Hx0ckReWuOCxqSpXFe3/NHc
fc0SkShx1wVLUjG2iIYY30dW8xoeRQ/tZtmgH7apKYl9MAVaDCXsgNVRgD4A0Uzs
SWIt+Die/aMFFnwB+lIctjbsyBQS7CsBI52QiTnjsKVTDkyO369cBJwkSo6X6J2Z
DeVa+qDpHbgyPk4qxBTJcapaJKlqw70XjEiMsfdVPwUn4jaP7ClNXGi3/riUzeVw
35H6Ovc5jGd6LHDQ3Av3dNYECWNE1qrng6xg/ixavfD6im/zKegu/s3VFv31JCIM
DK0qNRp3wlCvGxQX1uzSR8MQ5zrviaho4l1gA1zslEMB+9zEEtfJ5+hh1qxyQJkE
NUs+nfYynS53Yp61CHLbJuJmAiUhfFzxAw5rqN56ejE7i18SsIqBD3qtbKtvAaE1
pXJBGI7PLcwrVdC0x01sUo9UvdOqx9c+G0cCnKJMmU8WrKe13wkp7MkEGSdF4dAT
OS++2Vn4V+rj5Kl8hiakeYKbIaHffkww8c9o/FNK7sG0o39Nx6sseq8oTHKR2dtd
J+6gzLXfzIqkmhqU1loVg+9e+xHXj3GNf17JxW0GGQtP9kUS3HoKnkNmcXI9Fwmx
F4zecT/F9/P5+1kU7Nby/h/i1qkQ4HCx3kLr3n4D03rNM9hVzAFJFeFTjg4t/J8A
uMEKwWJygOI/RwHZwNTQ4M/cuvMS1/fMbeDD+6stlwYKvsXwD+r+/yKwsJPinU+s
oIxOfX2S5v4dvNCPfWVflcXSyPPoskijA5WySG8SUHdfnlSef6djQSwaHpbIyrHO
dxv2lBIm7pEzeUiTnVAJXLMJ+1hZmF/IGpi9i+fg7u8yq3AAV2ZG3wXWpNKx8XoO
rdq2Xd8W75uCs3Lyfn9Jjw8VZXc4Ltz4x2msMjlhUWMMugQZmwQha0to/jVUtJXC
elhU+vT/CAyPPE/UEOrLxS+/QNLwv9wNTC9O3hbMJeRfC1oNcErepfkMNX44S4b6
53Mx/UoXzjSiIyycXtG+24uuq+xev+O4u/irFFsrPV/IhkuK+A7RUzqnfvBT1VmW
7zpdK/GDBzsmf8pFD8RsURgHogR8l8yV4cVWePSLEvpp3qZmO7lwnRi9qQyPJQ0E
E69QyQUcgzv9TFv2Chz3JpCMHhQE2xhIxbdXs3E+yG0rsuiXgFASaJ6XYa+UcCs3
IH+2U9q3zSRP33IgJFCSwwvPE+EjM6RhUUCZN66TMgJCWDJt9ahIed7XZLgujTnH
0exE4t55X+KAB5pwYSe3O/94ACkaQZDpfjff0mc9ND1h0DHIGczrCGSwnlOV1Ojz
wHWm+daFOfJuBeeN6FxlVStACK52qZ8AJ/c5TA1GludmnEMPQY/tG+IR7HDomboc
NwaXPft+nR62qi+CYuU3DYrb4UAA4NOWTHUq+f0/Avw3WL9lQLG/Jd+i8mxyDTXT
whk3IS4Fn2khmNk1CTGsd8aQakpTAsyj/6DrAOVKXEE9y/skPvn8yJGUv5j8aaiB
QJLX8hoQkyW12gLtiJmyH488mSwATA1ddGf+SQR58lYs0YfpNiDCySj6IEt6s9JE
2FQ415EQhRdW8Q0Q9AwKVjtyQhV72APvt2eppytdDTSNS/8laqH9lo9zS4dULCV8
OH5JbsX5wafJpE9kC5sszu8TvrBeF6QrzG6IVWkhESja6MJApzKI8j7LqOCU1jgS
7ToNGzbWl8lGiviSjYetNolz7DLYa33B94eNGPSRtWP8YxQ/xJCgrjMock2AUFSU
IhPXcWXKhHuRtgdkQAl72unur4pW+CsXwbGY0xhSf6NMKtMpnSbxWz0hKIOYmdmJ
Sqd2tsge3+QUaupdta3LPh5aGKUQ623b4y/HAWIgrt0MuTFdIP0QqLlgEugZgksQ
C2TN3d1peVQh/GQeuu5LWGkKRQjy1t3PGkQE5umrM7UwUtU8r2QygWr9AUDa7phK
vmghm6oGQ1SnO0oACgE6j4Vh2DgKE3X4gFDF6GxkNY3+YVsMP0aj1e5U0DjSP5lu
/vYengz23Hiky6yiPGaiE6mUew/qMOfq19DIl1gWYHUiTYsStpppGs2sL6iNK4I0
NF+hg3Jw0uA6MtnWo6oDJYhQA7dPWPkdJT5UcvFGdEj5wkOQhfVPpNRNacVXf3sk
K020YzZvraf8BPVy9it1X+YhWGc+H9uF88HaRVDoC2ey+gxsN7ZkUW5cI847uETm
NcY/iDnTFhWwJBtJCNpCexHucTPYscLhJx9ra/C+mP77G8puLb+fIWPGSf1JQRRY
7yJWzyPcZnKCXnPB/QGiYAvuqiC3uYrctdEmk0MQKNyHmr3rqOkS6S80iD85q86j
LirBifYPe6aUXdSJa8bvUSMwjyddAo5ihE22Pqp3wAPIEi+6NKq0StM0M0PQ9CQY
dRmG//1iEG7MtCd76YO+v7MaWWcG02+AqmovGwzlzWnhIhJNuMHT2I9F3pc95C9o
ZYBWIa50ceAruMuJfO+opAFZXhLZrXGtfiXU+LTWbmhNQ5C0HyP+UoxUSwPvNwJZ
47wSVJnzUogfHO4nrRXhd2RhU6dzVvouJ7H6zWI8XFkK97fAhmuPqYwkb0XRkmkQ
bPRWygE1aOax/kTrf2yO3yrA92KU0HrDf9W5wTGZ8g0HbU0nLrlz9UeWuTH3AmrN
PJqydwIn7/mBQdJwKSNgGAoG/gGegW/29gu3Ha8fjKNzhre57pchUYCZdnFrjYXB
I8BQ378n1C6UtgrOwU52ZP36p3A3LX6EHj0k7iDiQCO0OS22Erjrp+ta6T2BQNwe
umYINVIcRTuTGCDaIQZHGUOkkSzVtYJf10Zy1IG+t9IZc5uZTx4+4p4MfJxCyUBN
d9jE4Og3A3COLM+Qe/QNcR3kApYLe4526e5XNRj4y69PP1EwjRZbO9+LMWM7fQq5
CKfkrYSPIatLwgv+O6je4yyMAmflNIUXloigaai9hVVnq6idPqQwqE4OrzQcylaM
2ihDT1ledwVoGP+xog+QuCboJVymB38OZndIkDw+IGJlh8vwMsTZ65+F/O0IuGhn
SjSkd58G5GkiY38ZXYoJfFngtECZ+OPm2oYSSkeUBK2vPKE9xj23T7sWQ9RzaYET
AxBCC9aZi1tXh9PU4gvVm4DTmbs9UvYWcvjqor9wDUVlG6dg0O+y/kkjcHHQSk/z
mb7dsZiaTJas69btSgX/iaUyQwsjhqm5vWQidOrhhK19YNO8LR9U6WllSK0POMvG
xwjGLw5c/fjYf2r8yw41h96oc7n5SazlViyIK7jOAGCNlUYuj/vvrTVDYOzJswHe
bPYk5CyCOfYRT5FwDpeiOyy4Mn7oIvpXfiEmKRlE44bNGIkNij9Ln6e9kNkaflFu
UR2dcep2YxXeEhI+WQ+PvFw6G/6ztdbSS6b33kd203yxZ8uVK0/Csb+bZqD/Fy5L
UUHOzWs7GdVZpHAgKAT9Buy4nQ70xbouBUl1UknPGw9lJk29Np9iaAoNJcyTWdpW
XOaYtqdLUl9H/rC288xlenlSQ2NqUS9TKRR2n4cjwQYYMxVg6SsoCklDgmAOTvq4
a2yTEny70RY+ZQq/YNs/OY9hIdF2SJ4y/Q3QGnH5aJU9py8tHQC3vqP3r9XJmNeo
5jcrlZZxrwkQFys2AP3nlXd7ijld2FeU6m4rhkZnAwdrCztrI6Xad/1rJ8Vt0WG8
AgNJUasXbxPjlfBBLrT1l8PVLTGA+vErzrKrIAD62BPKZFK3f5LbTJltIl0lOE1Q
0fUGKshmVW5WJ8zfY+pNMCkcd+we3vQH0VNtoN/ZbxFUppRJ5WJXZoX27S2gbo1Q
4u6Fhh7R1GxmuJo+KKro2T2Ms6Lzcg+znNvWJsX/7EKjzvBAn/rxVLpT6e+ph8zR
weUdseraqVtLUHzdMGfm9P96KNGrwna2D6RwYTasqxsKrPeFMnb5qXf2cDq9XehY
xlUxAM18bEJG6+QlxDkS+qJZQLimIb6QaCQfpZOi7ZA5Mm+LU4EpbBCX1r3M3iZV
GRKhPKcpbiQoAu6wF/DbjpKKO7o6+tGZQAe/Iwj9p6/4+KLrqkSNGeBKDyhWz+0/
NSP1X58bWdy4TBZ1AyDe6dmahpUkiWVrGMF2OmEdzFKqEHreRrIHj/XHcuiK90CF
Hzmf+imfMnQU9GFoPQfaVEhzAy5b1eOb4RhvVsJcFBpb8zRHTItvoPyD9ZFsy/Hm
g6ezRFVkQKgDWcVyMxid1tmxx9YLVxc2riYorzhTjOnYvArOERwknmYwg8QeTZLf
o9JMoRwkNzMIuAfPqTO3i8+tSiWXRNZEsKTj2ZV0YVixZWk4HwPW9OPAhGORpetV
0Yysq5L2KGjdqMNCHdHNRZIxZ8Z5uRuZrXodGNgcvu0T77/v5JGUHqqIxdQJKUeU
TDgrjvdu+EBntp9tq3tFKSP34uSxIcXeEkWQ6zJ3SWtRd7jmeGHqzUo/zrEOUNaM
7isJR8N32i7IApED3Ubvrt81Ot90rnyuEMB3pxdEpAfiIDCgqff9bL5Gsc//HAqP
wZLayeDWoSKrTpIYruz+sBgmKUJZu+3YYWiEwBtCoQu4KCKl60W2zcahnZpreIxQ
Mz3oPiNrJ0pYv1JHY+un7DTHe+7GI1/vLl+rICGXFKmHUIF3bP+6tNgvEf3dmvwi
Lz6x10YPgnAo9lBoKhu7ou8cvztOaX01LlhSSMUKQKVsK4tnoH6ftqiPIsnVJn5o
0rssALauZqfpTf53V08dnZtxVUboGGPkkjzaz0VHtKsQCK0OgVc5RBVrgdIgaZ+V
8Ct4g1n8MN1CmEnUPuMn42YYwNSiar815VguDhFmJ8A/k5SjE9NYYn2LBN7gq74L
4NU1tDlT3udHsID08Nem9vGxhhFeHh85Dcg1Y+8PZA8mk6NPx7rnEbLnQhKwY2kk
yJ4jw8Dv/Gk7jl51R0oXZ0mTByMXBd3KY284Ob0IYNhfSTNsxOmGltrsKAPmmk2C
kDLhH7iBlVtb1oxlgg9Ur+55SNX/UL+rfgirfoMwcuKr9c0GDTcB8FagudRMN2o7
9Uj55c1X6YWoaq26a/kXq5KadJHlBW7ZUiETFxOenFY/Y7B1GWA9MP0FcRXydQsM
w+Z9PeMQdwQdxWxEpwX5SQFY59nKTmtbKdPTXTdkN0pU+BtKJwigInlbAmPTPqL4
AkHCfLKcB4Tyx/kJsVtc3VhXLmE3Zx1bfo7FPtcDhZo8wovNDg8c/LraSiflEfaP
v++8eAip8NmwuQf0VPhqSTOc+2vZyPR350+QsBIh/iN8kO3V9X7/64mbFgooBWOi
SUYzAODaoOMgrETsn68mtAMGIHVOZsJKrbowiRsoMhX0RMwHewE/1p8PJr95UF0I
t7qC2z+tAChFizrgRzxUeJlNQcmq0GH6eaTlR5uQhz4POkcY8/MaPuupz5rTqOLm
qs8WVBe5IOYD6XXwTQNJAW7D1Z9Lkc/zmd4+jIRG2pv7ygYqDfl9sRHSF6BleeWN
uQiVFFOtO6V7lNArg9mKFdqW0EI/fR7NZA1ahabNK1SpBY0bI4UHZjeJVUDf0jmf
EDh4+FJngWtqTIqEKfAUyNRUccOLVruuvzgiGynXRHUaqi4fHYHsTf6Nc3LKxmZQ
bV/Su565MA/KmKBFUpcknahRc+kWwRWuWtL0pQrdtQiRoCypuJtm2It7w9DpKjSe
cIYYGGX7dW3bs5gI6ekg+QHgaJGAhTrvJ5WM9vQ727jnQRov0HKiLl70wLZQ6z+z
6dzZ66LdrGKNSELTUQdSEuiH9VQPDPJogyiZFXPZ54lTwwMtrvLK0lJFkH9ueO2+
CU02aI9jP8yQIBWu1zFkGWzU6ZfVgt4FeMojt3FM5KNwBSkNnLU+4mHc287idmcI
bhhfT1S2wxNj0XhGY3750Q1b8Snf3st5qpANJtnhPSKMHslSFr4QI83CFa/rW3OS
SXevCjaQoIWsDo2sr1t4PsPjrZ5UfLKFs2UmJ2kCNAU5kZ/rvkxQ7gByvUAN3LY6
J2GzwsgAS3EfGrxKyl0PLqzTsX+aqA+lL6ks3yexIOoLtx/4R+TOck8zrMIxDtPC
ICj9qc2Gb8ao8oD7HNWunDR3Cxkap7qQAtB/OBI6EVi5OD8YMPG+IMIBzb26wLcD
XLxa5GwgTykPolFftN3Os/7b7OA1aphdBsQlvxLYVmuuULtEUOFA9uQhjiXL+aeT
2pPgQCqklm4oZsjY6g6h1pjteVVLH/sNtL894HatjxH9iP517PiCYK0O6eLLP9OG
Fhkfr1HkXiv3cjo6Nt4Y6HvN9RDP6yOUPulzYg76CwbdOM5YHPBRWYy0uEfFX+0i
65vvYTGyA/WnUlmbkYynAdJPK2qXOLlvyxmdXqph0042CkO+cbRmiFGfTwoO0R9u
1LiKnVRIDAKR4JY8thzofhESEGrBuF4zNr9ucBFzHpa0Ir7f/GWDgGmxc3qxcnwR
vOTcR7gT8rzlZEEO82peNabDg17FoImK75f0ZLc7eyoE6DqT1L87qIFJqxYxzZ7L
Hw09urfKItUSgA3rNIiIFT89lSFLeLkkYhJgWl5vWHU7iCyMXewTsy9ov94e2SyQ
b2CX8Jr+yulb0sDzl3+Bax5q+2aVw1re4HfV2t+mqHDIoG43W3Gft7Ljo6wH+G9Q
WluAJzHXcyHEc4oDgIWmZgkPWbdVbu9ZEtn8h5EUiPCNR2+y2I0uvolLRRNQmozR
iSGIUuLeAK/V5YyGdVqZiWIU1KsUR4v6zOEQflRzDendLSsEeh2bL43BUK3ELd/o
KvJzDbk6FWnwhdMAU9aRLIVJQ/F99Fa5qhIy1CHpLn+BuiJAaKTSkHYiaV4ZSddm
foyB3UfQrdbm2lnhUoAjR7UMvuCLbyCkooU6aECYtLDkcukEXnSrIbD/s1f66FrW
sFbNtUIPb/xEkbFTJGWnExOFZhI/THqPv9VcVpp/hd0Qry5XEHc1A1tvlkIZtXgm
i8284o2p30ECEg0JfVBN56t1f6Hk28RhR3OS3FjSZ3imFmvGhiPgOY6ZD9X2ifLV
bVbP5zb2X02btmFnSr9yavg5MZOU+M9LdffAuhHhMkBqLVRKaWFt3+kne0G7vzRV
11zaI5631RHJlCNufyHX2rt6GgUUybegvC4hDy1Z/5NvBFE1i9HzFtiHwi5kegj5
BTfbcfZIQzfKU6BDzLNic6paChFejcfM+wKp1LHJaZCWeM43Kc9oZHL4FYPRd4h1
pH3wbQpZJBxMi1GsIvEqFSD7pMm/EWpbds64XWWdN5FOWEiFVG3F+W1/36MfGIH1
fMfeIwXS9BGtSQJa+c3Vg4eaT0OJh9WooExWWXJJq+THjFus5J0D8Nq5cOqi5pgX
Y9ObH44SfO19CQBRLgzvRx5dlUVxvUDe597CKqeDsaJgUZ+6qwKMllztChMczjRu
h7FNBT12kXaPOr378Ww0MRiYiXlJO7nzSv2vkAhO/53dGfItCfEcQxgtgox/CNA0
Wa6U5JOoVB35YK6XbDXzx4Hjn4pfN75HDdVy00WeRVylXnCuWE22Ckg9knXoqBGI
Kvl3Ss0XuLm3SBtqHoA6Dz6ySyPgikd7ynfRgUEkheRQvC32EXocSdGdARq4gNF3
CEvmkAgnT3U9BTmBvNOmTVFEc+juxxBfB9hVS8FlfR8wBaRAo7blQlehWeoPNCLf
9QbYNDAt9Rc3y+tDlxA6vdWENaTOid8vawQ3+KwR4rJAtSQf1YqFgrRP187u6eTk
4tx8uS/BFR3FvnAObGR3Dha2mLgqrBr0BN+ZfGeD7xDdhKLuYZKKnvlII5RjlN6N
D4Y3cNXWygTm+CBzOF4z53A6sP0nxiNqX6xxNzzNFyidciRSF84tm8r/mMT4oXEd
iUTUP4bi+RYpq6iM+NTPeKz2qjfwjcodi3gQThir75XHrRaOqaf0RQLM3DJHqBFW
cJ2E5sJ9HDBrGhPUgbF21L6FTkiEuD4kYpxGtagCdwZ3pxMsuch7sEjet7h4fBhG
BxIFFW/U2TW0ixJL2GaywWH/XrZWSzUW2O2cLEKe/vDDULirK1UFO55nhyDLm4d2
g5jwjACVI1e5K/BzlNYuI5KpH8F6aODxTttyQuwHz77dPiSxQx1qBBsMBA9CJRvk
90fHSBmnUoAYjcXnhhHdsqTVwLc2ecpYFobNFDjfOa57GDFWil86MuNvTdSjrFVp
w4N5pngyJnzW6ZDAlqocn/8OHWIDEAV/PLpm9Wy79ROBBKw57W9g+xJDReKUAwO2
0U5GvfTvNzxNfeYsAtJwDaLt10Hx+Oipgmxeocygj6JvTJ774Cx+1vRLPyrhWzOB
8bG5/86HrFnTac5Bz7MT7HBseXv8GY37zlSZW0hgYuTMAwqBk0DQp2+pzqbqkmEK
2l1VArc/mntA9VVfEaBsjt7FuHMpJpntMZjjzDsExECjC4wLcMP/Nj+jhU3yRCM9
jyky6p50oIz3Z/bKAlTeQ7bV1Rdd0a48+RSkosBuWvYGYd3cEVFZPdRynSQXKBAQ
6jaPvQ4O5Yx3Q29NVnFfEIExL52E+cSFvkCg+o7/E2VS2fzu+hqgVgzwtCT90rNc
ywVas7qh+0pFon4ZVF/ZB37TLb5rA/VkLh01oj3uxM/FjeS2X/aznGRiFKJEmYsm
WODkxzmDqmdzOdpHla7IFenffxnL6ZCXRQ8KE6W8FDi12ZydmqNVTSlxuFPDmBZi
970+soXdbcp4cDbwsUV8j6y685Gr5PmiuJC6j2vO0AXamP2OrniLuDT94lqxwVp5
BWMGe6DcHPEF/BHnVR6bBR5OKiCkPG7aryvT4ZU6gkaB7BfQW2J+tPV/syszCrY9
/UcTxhMohhoHN1OfummpqZoGxdueehCLmBM33vKfAiv1pu1wmEizgxAIC0KxgWRP
5YglRXuyT+zpwKW5FnFaNBwJFVKpzaYkHR9FBi41x+uzUDSqJ7eoe8lWM5f6B02B
AM9T2yJzYeYXmkDfl7ZLV2Q0iSEuQSMAPgYWgPvT6v4p+QQ2CRFB30abmc8gl6pv
Njid2rGMI4x+O4kDNBAIVps1Dr0Z1EgQlm0zcmj1CeeH+d4ZGLD/hiayCQ9Ah1VV
s88X204B2Yxrdxpf4MDEMXceRQ+aHN2Rgwy/MPDjcI1qpXqJlfLaEDSFgTzwuqpL
IbFufQRTQpXyUXwVybbjg1+f3hDKbzidIyrD/flxFsS90r97o1QfR6h3SdRFcbZ0
mSwjmgn6yASh11gY6KOUN8iLNvnwHEmUVpRQruIAA6Ri7dMeZYMgP2r5VlmDeiWt
5Uym9ajgVrOfg3ha8iiyOQeGRtfReXzWenYYKlUlWmVI4cmSIxELwM9Wg2Kue8ku
09zPZdumfa0M8w0hrC3RimNRJu3VafXY9gDvMbJxhP3RdhyMOqDffZQKr+jXTZ1Q
7ysIhY1swt7UFiPstFQhGOey1sMgmfPmyH6GXZKwsIAJcWah48XlPYPfRTINcBxW
gHWHIzBnnH6RWzVy5ya0/p5TaMNSlKz83LczhcNU9m2EZVhYkDJgEro7gpBAYNA5
EEAKog9bqOIsRxy+ZhjwNHqVYQmLPaAQHtPEmGdjEBP1phf2n/ysr3EZ88wf6B9p
geXyo8K5HZl97KmqV6NEH4IWCG4tVI3Yq7h9zNuzDILwl1rdFd4oEa0bS6AQdqFX
fa2huKuHcDkBzRWuXQpR4fo2eabdSCBKVngDYYXr0RiQVdiuQCFTEJI9PSYPv5lG
fPtw1uc758tKvqhsG5GaFonGMp4rpfTgiX+9tLlwBxNjuYX6UC1+w40wOpbToa6j
6/0NHNXRbP4dIckF43Krb1p2LgTC+IjGTwptTDDelxBekTAzuyaP3odhgHaZm3d9
G7A9QXHUmzfZnmDmb2rw0ZjLAItQb/JnfbTAYGvHPTKSk1pV43XdVmnk7htsGuk9
jOjJ9PHl+0fsuUGqSrQXSIWWyZMhBcJl/jMjTjmj3Q6FGfGZdocqePcG5b5bUtfv
HSL09EC2KQHz/QZ5xwq3VM4l9iP6DQcFx0FXN9y5G+vwlAaqcTX5MTwMAk3loSs1
J1j6y2ztuzZhMovx9QSMK5i+nJwqEgh9xcRGow5LUW5nFLQmf/I6K4RByPY9junK
qNffJ0JxiDqTy7zVjHPCGtq5tO2oA/etWBQICLVcKtlQ49D6wV9FjJ4oJueY7z+G
cIhnpF4VtDANfku+Pn8gCebfSKW2sVqF3ivmYggX9Q3514FOixIphxcQvpAUQR+n
nucKY0fV/Jb0jCVaEq6vane+kOPRVeq3kNprUu14GRmjjOKzR+DUic2coOt1MEYk
LgfMABRqjusC64gaUATViLQJyApfhBViyRdOdXbETlwQ/9kANLJlgRCc91S8vvXQ
wKsSGHWZ/u2wywzn05500tWnXH+ss7Buqil4uGytpS2Rzx55umS8hO6JEwt928Q1
4wHHg3Nd9zQYL7RtVcYcKFZl6XWMiEwGNlOpab2ziCrkGyM5xyzgt1ufL+GFXhfd
w/f9t2FGwzcFZHomPwplDys+uQYrg+IxwL/qEaqyHPw70aELJGmltFftQhxLLsuw
4H2sdxrIa8iWbkUcXZI6dhNpPF8WwWC1UhueOfxjsiq9JR2OUkVsrCVeQVOmiFwW
MYk4wNpcQ0nlbF9W4qMjIu25YCg7y/v1pU3IFi9PtTKzq/NVCObNUL84Xolq9tbU
gT045lSYdh7Q3Wnq4ZAns83XWbk8iB27eZlifZW543KXwCQj93AJXd+YSJVIKJh9
4l/687Ix98Xje8gzIHigv0F9usDvf4cdDKpb2pgDFLSPB1dNLzfBvNAqz0nJG4+/
Mf5Tl2J5ecEXVy8DrkTIUF5mZ7U9rQplF64kcncLJCsWFagopCPymUQrehp22YLL
f/NauGL7WjgsCgdwasXxRtNkBdmc2Eo3tSFYF39+stJjCFzQZNrG8/zHcgbX7wSq
iqLRlG+nGslSXkoEISfpSC/TKRm8X8TgHeuVE4+K8hP8EOXjounjFtxWgWZX6VQF
QIYDN2q/elSq6TEJ1VPCPM3DIqaFaeai/MIw1etur4VP32BB3mNghiqEghYjOWeY
mtxZDWPTCEu90MJtmIqgBEY6aw/FD4iuPKi3jbKGJJeNITr/Ax0hMET5EEADGP8x
ufMAg3xmCJLQj3qO4ggjZWWgkZD/2Fpbv91NCxdq0rU/qc+hmhWjgcjjQqgkC6DO
VzzaXRaI+dc4fslrrXHx431bVjlIjxkhHVnlHw6rdrDH6uU8ToBcPclod/P3Cbu5
cxgdo/EQohc2ev3iLpvNAWYByYJoEckC5NVkVXC8OBj1HkwQwryhWtnQ7hbrrGxI
phd2U1gD/Ry378UCjI3z6w8E8G2aPCGNeEyvCECdZx/3Es02oZPMoLPYTMRrbvvi
CAt8QoXTW+2eqqOU8ENIq4HcFXfoF1OwlXpePfiDwtatplFJ6Il4sToYNlkPXXE1
pJZWivIN//U95eVnXXIzDP7Naz5bCxMBdvsNb2zAIwivrYCCBm4+ct2QZiCegnoh
R1kyB1arr8mGHP3rnJVRWZ3qMZXU4rvc7f/l6d5wCnwpe4QZTzokM+qFF0/CnP4h
GCH7S8Np7sFgLV26VO82zZcHlcJlAVpg374slkP8YbRBJbhhMzMpKxHeZP91aODL
UoxNns0PecxMGkZBwqQFCexHcMhHVPwesRTaVotF4YPseAFO+78emTf2mFPnjtD+
zkxcI/GikLpFVo0ZeOx1uZZWv14B6nZKmjvk4u31ZtTToJoqoANUpJWzsmQu21Cc
3MMbMtafND+hqgtMqw56QGHlZzpL49843POI1akZNmBezVHc0k6l5cC16GZrvSLw
n2vLgT/4PV30IvTT8Zz0z4ewyJ6PpOLKvRlp81UmuJxchvegn8S7issdKl7q4ENG
5q4UoIx9VLUWwlTmmpCiZR5HKiRw/7FkeDG7KpsZ90O+j1gnllSkMOdLsyr+A1pY
uDD8YTyYNRAT+jcpBbZhoVvVu1j1V+oDRQMBbgsZmqIc9plgMmu9ufu18sWI5U5m
MOp77uK21bmBJqG6KVPCCx/S9MfsHVEB8AKSTXDNwk4PH3O0caFSIwvld1K3IM7J
wYkum2/G3LqcipZzMAZ5pclaiYih+KZZzMdr7wd5p94iKvjrq/zIuMVVZUryWkzP
8LKHLmpDZ9lY1G0tLbXAkVgrG/mex0uV83Jped6HJpHL5n59C3WabwBtGoeF0Pwt
OiQh0PmuU6xQ0yWgKPGDZNsDySb1p/ryGf4WkmCDOtC1PAn6x3LW5bMEx9tgUt/E
ZiFwNHCcgVRff9zFFGh5jrCdjNHmKpWGSlBd7AGM3XkIxPeMp+fzkhKlBe6MifJn
tM95Pfl81pXuREoS5A+3SCl2sHz2mfFLj605gZmZ3co7jM6Tvvye7ivvj6ihIpbL
PXFcoOh/PSLw76D+DMjmrY5E4YD3tVnq3asFUd+DjMb2C9VtsM61pz/92x4YuMEu
EWq7pUFlTNFGQaQiQqTGv+FLQaTi0GSXy2qTmwW2cF2Xg2Rc3qKJXQQnGQKRwnPA
gugixqRxoMGAAhvC+mjLBTlm7mumjwjEcovf51NFvsBbHabEAaTPLSk8GDvbeQFN
B2PzcRaSnJaLOWDzzjh9TbmWr/GJlpxthVIFe9bspsgZXLzJurkD2XUpTFdOEYWL
noBA3dufbis+oFkcpQijEDJpXYC3mcJAeq/1oCyRweoiEyh1jJbwqJLUnqGSXV7u
XXG6vPFKFw80yxzP+LLXeqzYNWOP4p70HWJ+e3VZw41jt+EHwlsRHzzD4VW6DzXg
9YR9sBc5efkEJEESoHUeD0EjOU/YCp+B6wYF36WlNFj/erhfv24TdjZkfJZC/mNK
w4tHzt980WCDIvyi6dJl2F30V8IV/EZ7PSw1Bncilg6STQrGlB20EuBIK769CGCe
T9zGQV2OOpwlS34v78JW+4KXmC4wmW+YM2BpVJ27/ZfY0meAZlyqrk2iNT9Dtf4X
+u/+IANkw307oCM7VwxogIwZTKVQgPMrzNjq+vbY2I/BTX8aJUzVe9uL/M3RAueK
rCGBKRycbtuw2LMONnys4tSLji/XcxcpRnT1ieyjOemnu19/KboWqvakRVEg3pWQ
/tWTQmHMApZSG0hRiT/JC0Cc3U8VhSXc3NJD5lnFrx9+tGPUqlhzd5bA8wCEQ+yq
E7WDUrHSGNOOoiY/VSV8z3aXPf3boVQ+HQeFn8qbQ6PlMctOcL1Ofr3wbnqpQcU2
DH8jYi5ACvQOI66QX+U9QvY8vd3cO+vcvB1upX12r1Nd2bWBKy3K5+G0+nLFDiES
ogCUO2JlbnzlwaKJW8WT//OGykp4Vn5fC8go2gADJNkG9uS6VlNtjWeqgTEqnvYK
Y27qt4aG3AJrKAhNy0u7bmC4kws6bMKWNgs4lZMnF6GhDVA5jNX/cF2EVNMVKfdZ
O1Y1P85HBiGFZDdm/vPz8bsSEVYz/rCaUyeQsgVX9nxHeRZhgUHZGRWaxmplbMVU
sWc69PHc1oxOcs+e25IN97O00onD5hNdvZWXVcokmiUJgslpsOKnvlmqnIErM+S+
2Psdhi1Pi2Y1ZXiQEv3K5r2VFQ3Nb2YZAb781mS1fNKSyDkGdyPNxedwirsq9//f
mmDmaiKl1MweFQL+5ctkYESW0f+MXwxqQSmktn/SnGBREvvAox3ygdSidxKgmleh
wc5FyuwhGHjT7Pj1AR0xxi+fiwNUdVCfiGN28xaUpbfwOXfySo9BYUrip49xOorB
paX6wGihzwjIG7wu4fVDGC7qbAiLkLJ53Wq8QO13dxH0e2LN1n9IFcgTpYO9otgb
RQlG69OySmev7srMAn6dHuEDSDmOB5ommpmzS/iMpO5k47gp1ODqeBoVGKlVDydV
bXQsr9B+RGp07HWReOxfbB99Daz1pWtLQlXYl4HsL+G6eHyZ+W85XG/9vzw7puQE
SC3H8/WvpuqgzuW+nptkg3gdoDD6ZGSgmmANyyWSM34rUTF5Ubw9sQxsfX8kKDS0
Ovyxh63jRCzX1/Ettfcbm7n0wyP1gY35BK+CIM73TsUXib7ZmP+0l4yBXMo6rOsP
1655TlW8l96iVDbBQz+yJgRrnodcoyI7Kxm+kUfTxqN6xCF6gKPTdRJfIv+HY1Aj
m8EeclsaI2QUXHLn0VM+8IoPbEr56qH+gTiySqzcmdUC1vv7yKIx7VDQsvqiXpr8
cwiLm2QcvIqbHCvwKScwK8AtRmX8AnWN1xGLXsmQ7AMR+SZBMBI38QEQQgjayUUv
6NCfUNjvhKe7kXs6WO87TzSWy6l3usWrya4U+tXJSiqV/TnyKqnm3fbItw+eHSma
/MdsWni+pWkZ8kDAlA04ZtnvQDibv84YJqfR35h/atD2eVuGzmbkl5kJDVdVGuyQ
rLoRRpd6rLA87I7MLxg84IK9LsivO7m22IiIZUt9w74zrsDoTM/MpC6RBnbuRUPb
CUJjQ9PWN+/HBfMa/+c5tj3tPWcvJmhM+kRO7skZ0oO3moX4qA7HODQjM4zRvFIq
3w7aC+cmz+wBGp3rACWWDcvQnjy7UNgpZzcu5LmQYfDKMIJfHCi2/vwkrCm5aZ0n
8fw01KJlRBx3HltJGA1uvq1klM15vHKypCuOc8KZ51Toqz8jSTZrhFc8y1NsUSvd
kuZnarwQgnPHKkd3QMFM6ZN1q42sl9lzbSVJ4pDQt3ZXn8hsuaCkEX3DIopUh3Dv
GgevFSMcXDW1UMAKX+RVaRAVX0/acHfuDos5BdDo5RIpAjhjMLtKv8jV/zjUW05c
5bzz1OfZn4dmqoS2mowsxPR7Onf2HW1YuzxNjMvvxnPXeb9aXm2lO4ShNlWuqPYx
CAjBYxi9BCd6nt5/vZ5+okb5IgPBRzQOecP6qafSm52by0QiEfYfQRTmhdXI4B3x
CNZPqCQ8h8Va4Q81T1kcv6/cGhhcc7G2Mz0LRFA2mL84w7E2B3ti+6izrhwCdByk
5f5Dsa3u1YowrEEV8xWyKSHwZfYGRyRSccEOaC6xMjQ1Qf5YcKz+5vBIkOd15Czs
jbk8UAsGjEltKWDTorePbplo6L7K5vuADe45sr5MmcEE0VrayJ7sh6qiJySsQeS3
k7akNOi2qtZ97/zonF+xWJ2JDwHBJSNmX79UqEK+wo2S6eWIGpm05wRLqQkSlgAf
3woEh3ZsWIa6c+nY6zK94r+n5kM0/ycx4rNIrET3sZwpwOWvzXLgUeFTeHmnm+1C
aMi5TfB09RTd1hkI6EOLzZFhFxBBWaPmkv6+RO62rzMgKMv8s5NcB2eMrHu9DhAd
V5gxCxqqL0fMuI4Md4rgfSAskqOMIL2UBt+7mS2GdoSDqddVUc4mAGvA1Mq7LuSZ
lwZEbi6ZeW4xVzapv0ImkFFJ74T0G8QlRUvY07xXszqEaUTznwZHv+akk6Rv4u76
+v+teT3VkiEKMqFL/Oxz7lFSWfBx6c5q0WEbcvmrS8VLe7KJe5sLn79Uhi/zIaXa
d7YCd3CAjzA7JocHkhWuNlyKzgzwMgfezsZiL9EGcohBHrh+FQQBAmf3npdzg3Kg
U5RKvjF30i6/1Yxv425PhIcIcNV5pIGsGmdW+55hGvwEHoKt0qbD3c1+1y+IS8an
ma8zc7JTQ8dvc0mLbHa2NOS3wRootnUbh0BjT4ShzrZKf7d56cyXGDsJ5/74amKa
2ePEUF6a9IbkrmgOOr4Dohtyvt3wbUFeyZBKHB+xctUdnppHdI7Hx49mU/VLGIRO
CLs9OwYJ6VDdDYFnKRQP5/a25ZtQL3k50cILw2ItL8an7flzHNjpzO3vOQy8Vqyo
ae60tHkHcczN3iU3s8TVCO2kC8qW4EQ+RigENPunIVQ/onO3Kp66LkgyXcytHZv+
Sy35dViGAYBIK+2AsFEMqa+niBNIwIsEvrlNThMYgeLbW9e3FagJjAf1lmTNxePw
/Px5Af1nT/+eIfluRj6srAt5qHoBpQ7QN6rXq9RSqUk9dsCKZUv83+J9c1YjOTPL
LiWyVxkgHB3bWf+Sg1y2RX6S8UfXROGfRJ1wdtbZ9oRFYW1U650aSqDym/0TYE0I
c6ZQySPDjDMlvGhwlRB3c6p4UW8nBgNB/Zxm+ZyTflkC7ykYE72Rntss4kP3Cxf5
80M3ITzIhDguvW14KFnsHUL7FlG7ryFJ4bo385yrEfXzEGI5dm0cDCtggl8KaHVF
X47oKOefMqNHCFhzKIJxnQ3RhmvNBpzc2Gel+qhZm9kVrWKIuRIq7jAO3vg1IUUA
PjuDa7ICXZDi7rWvOorHNjCgdJnBhlkCZ6paf/MiaO7oTGhPeiYVLGhogbamtBi/
BGok80uBxijHTt4yD4yosh7KGvzXc5QzJt+rGCLPVl4B0tl8iDJdpTdGYm1QyxLc
Z39ZLFIQTOY4twWTaeREgLV4TcfsODL6dZVTRSPiL7tf6TGrkH36jJoieKsAnf8C
ZsR2OIpFrK7QiEfrpL6FZpzaGhthmEYk5kfE0+jpjIOIK7R1y2Ov5ndlnVqnZ3QE
wkFSQ189wNYp6MUmx1i/ZKaNsVmniByclnh+kCC6G2DeHaujmFjYMHFzcLaGsPZW
dLCKuKH4xYZxaELXGcE9flrCFZVDQmNkSO658u7WlQZMnkm4On+1WyUp89yynkji
Ax7aTfgn3+fFWBLAvGcVXFVdj2VXGRkdYdVNlAks4vO5f+2LAg4kv5hpg4rIxH/l
OcttNCY6QNsVOVaUdg2H/uFLiJSoH2OqgdAvJexwzWhbEHvg/DWrzMPlNxVC0J1R
6qvIg/0ETN8t/U0IGA/WKX+rwSfyZTj6WMUZSiXovw7k0iv9AN7H5mUZWN9MV+UE
sEhBE6neyKknDQZozz6gG0em8CoHc0zWnzPgZfVPzfuERiQ9lV00XVk/eYeftcrE
7e/o35nBbrpLPIzDeLoaSDXjrAd4BhP4NSlGKN2FnLhc7jeAwQuwP/Jw9sMF3Zmn
f80wt/zH4tswTh+bSXxXk4RzPiwfGAnQgLc2B7kVGskPNTnEmJnd7X3y20yaGs2J
QaEqVR7yySCdVN7IMUxJKIOc/awGR55TKOJGWP4qoZyQLUINFHtzObklKZsbMGMh
Zv1JPMPIOsJLlANl3LKykjEOBxBW2f+zeCnmiqGTY5uEc7TTziJfmHrLD9dwqEcL
aiHWBgF65Zcwjz8mWD1H0XwS2EZvl2rs4HerachcE7rkU8RnhNZQAD5KjCqyhdPF
+dUal0NNJuCxqou8kSPIgSSbje+3qvRwCbsvi8f3RvI0BIfy7BqtMIfQfigEU3G2
sKGOFv7ZH3tToObLVqf6WjycOmbxKoEu6LBpbr3KifNhGhIyvFQch1G+b4dnmNTk
4ieF7A3x9QZg2CUbTlxiiW6efU7iNa79Y6dv/pZClQfgta/iLWCm6hA7TpkYgP9w
NXwA5NVC+sbqL06XqvM7TvvApHinjaGREPEdkHbhMyQpGENe2g5QbavokdjI/vBz
f8tP6vtRlpZUh1z/vJNE/DWZfpyzXSMap8bb327tZNvPz+BaIahrZyfag1FyPcxs
MfuplJvLR089wkE6Yui40fxz2fUGuKRNrhGFXLT1s3g1Um2JoZvIs3y7OfWOVNpe
IN7hjJc/sEp7Hgz/s9nlU4VaFGSz9MYtILddBiteLpH6gdqtnvmf/q1dVswiOdQj
jqo5Q2V9FOLFXXcrYU9WMH8PF5otdd3stwsRwXkFPr8qzV9E/Fl/KcJJvvKkh+fL
Cp+XxouOrck+n1MvVrxZZyMKBEzB3zC+EKTFuP8qeikezg1rihHOpC51+4E/vG2J
VEkoVFv8op7+MEyJNtCxLzIDRXJkeXgTM/uQ/QvOm3H1HNyYpl7/XkX+TOfXQGUd
HE+G4qh7+RFQon2gtWXX7uiL8SaCb0gmH7pLxxjnNGzfePr44gT/NeKrrHQZK/nW
tYcrnWfdlc/554zeVgabDZxtH9mXFyCDnIC9e/X5UImaus7blEB8tv3q7HpLmZLA
qdwhZhE6e6QnxGnctQbljdpy9yU2OGJ9I8XsOkYSwQuHFGBqa4e5NLhXdXkAt3vM
YYnWujJFkwdDBbw78hsT3ybJYyGzwelPSSeZQNz6aTbA6B7DR2fFTPON6WrIHSM7
QO/zBqNXunv2LpGaJJZOK5WQxi/4SRarqyIvTo/gjgiFMB8l1+kPU7qma3QnSB/G
Ok9SCWfLaQ3hMaYggy72AAfnaORzjzlcLFX1W/7+RbA709Hu5dE/Fh+cmHxanJG8
eUPYQHKTKVMjp5yL/MKKTZ2dUY2KduVYPo6HTb1PaUaIlvmiPSO47/3IqDLiOW26
ruV7Od65R3vd7xX1A1ZX2Ybfqa4t2Ed91G5dfCcvmOVAZkZ5PY7uiyPszciD9UVr
mp0LHHZhQCdhYYn0gC1YVZMhYgwCXJcQihp3ddDCjy2O6JZbH4kTJxA6BQrSqSfS
itzeFjbCogxyU4b8qSXD2hhOE/vYhda/QFelJi/xPYI0uxgeP2hta+CkYSsODj3b
dMNkhpK1RJ8A5utlCZ8qGfc4504LRUgotSkoaeXiJDUxrLIGn82Nybh9UMDdqnY+
26IKL6o4YvqlbwwdcQ+TubGG5drM2WmHm861M6oFZYO2BeDLyks3OnyRTwcNKYI/
UcJZU/jqqO6dF+X06E/y/ozAMALi0xZuDqJ9cVp0gVsX5KjDxPyCRetjWwaBkDNz
HAaWV2WG4XL0MTBr8tEBlou14/WZo2IWaEf2I2URLU8+1gEo7B2geo05LUzYFClm
iyEpOOfkhh/xlcTrUgAdMi2lJNqpe6Wvp52rK/fYcC0EYvrqSieD2CwW/i1xkaB5
gdfofF14/5pOgWGy5zbS8IbYgTb0vG1z8FVNATmMFiigyoEcibYEhNiKDyOt0tHl
JR9RayZ6IE24TF9v/2pF5ukCz9XjoKA5mDuiFs4X+BvG4ZfL8kgmZQf784WSLJCW
tqMDbF68QVBp4WXh4U0NMLYJ4zi6MoVEXw26Zil9FBNYU2h09ti67ybg0ArJILq4
JLxf3aFsxjJjYhWu/vrGovdZxhA4x3SQHmTGvP941tBJyhKFoTQspyb4ePbZb35J
4JaYwG98XpgFuIrB4rbTwuBsItUfJC+s10/WUFBz8GER4HWruAZ1BpFGoVt1+I2n
uXDO/o1vuwVBgIHqMZoMtT7NocV0wRBjyTvx9vOFNJPFB86+qRKshzGqGFaTyDwR
8Fp85VkciJJgti8PuWLb4pxWGVfErmCNKdvKBBMqWyudBOJNJ9AQIOLBWVTYWnvI
yp2+R4Uo4CJon+AQ0cINESiD3t99jHQpNqeB5qiUEdmC+FuAoW5UG4qXquV5kVpp
rwM/4sOjwCPY3B4fUmDpfwcZI8cbKZpygKuFuMcj4XxYvV6L8BfpC0caZUJnjMp4
Skb79ZqKSKNeSG5jaReAQ+Gua3KyJClDJwSadP2iPrISlVQP9eIrYme/eB/MYc95
yQgLPl/0PV+A1fQK/bENnbUwD5fcQXd3/fh3fMu+uyDs92OjWP+MvlO5QXr7qXBi
df26ihzuqKIwQ0/tKy7ANrxTmu82SQDuKr3iCsT3GN5ii3DvctCMmigKV8I+UoKA
s4ZC5NDhdFECb3KcpVelsp3fCs5AUtvcJJ0P/Imql1Win/rhUbqFSGSiE9rl9HVz
hfpRFFkZ4/6FQwsOCHtwshO63Fab9PvH8qcywkyLjZPM4Y9ci1nfNFLwauOJxIFK
vdyJW5c/nCg0RoogA6Dw5F6WAD9OhThRZAGjLdz1OMvVz1VJyWwfkiaHbgQ0RWz+
rn+nkbbEkmqhHv+8WAnODF22D4UX69Ebto1IVfKRiVbGVe0f5vrXHjYRtOaAySkX
CNVtGCGvAu0HRUOx0Jneimi1kVFNRa7I8JyGz6UpjQQCG0sPuIaLnFOzLConv9cA
esCdNaMeDOU3BAC3095DBAc1cqyeJ4dyK7fqs97Iv/4nBPtLjKnKOOzBtBTYo+Nj
fYsNqkj8WPqUnvswjZgCNuwQJZs7tPgHls/bFBJnEZF8rgaTn/M3ZwwZ2/2B+E4V
RFOaQe46EqXn0PB3nc+wFkx4ndv/TYczBXjOF9Kf/wguqa4sYdL4KS1RRmAS5xW0
ZltJk7qZT6B7AScKVS32EhLJJXLeSprKK7anMxE3gjUUgsS4Q5rvEjTQAMl89gti
gPgezpWeUJ0DUPUe6eecPRsUE4qi3zBCe8/52Gtbrxhnev1syuZQaiOwiaSETOzA
7nZ0RhH9L6z/vlRpdl46iE85RBRGKuai5eQrGsj6w5ooWwz1cohJVjv/jTJTLbMr
wSDJjctzLKEle19mO9bN0+6KmxHcQsREvkHSdzBkozjYozM5VCeK6QY9PizAj8VM
2EDDnY/mq05NPMreOaQaxon4up8QbjAXpjDepGIanV/mdm3tA6/mzp4SyV1iyj7O
ieznBqIBzr5r82y3OeD7v67U3DPSaRaTcb0YCthSAfIFrB4bb1BQppX1yCuXLVmh
AubMbQgOwnbCfjXWLcdu0hzvKkUV9z04MWSm6L9bbcMCmbT7ecOeqSGNFVIINxFT
a/JPHqH55S+a+gmUn/h2BGhzagl8CJ8He7/WohtxufKyl00UB1qazRinTH/bnzV+
Ws0nUFLwQMv5t971pXvct3zfb2IUg16iQlG+rBQa8DFruAXUDOSQ8KMAao9Wd08a
TXeDY1ecCNmX5v1RQ9c8KErqWAlS05NCtlzUgRAVjuIF/OWqNGkZAzsMTL20VaMX
hOysZCwKq8rvd/XUH7sb6lvpV2wrqQBSAPdkHuxz5YMrUSMDvhDUQktAHZDGN423
6+AgjHw7ZLe3Tn3X260ZIu2JJh2madUtJiL+PaipiVqrKil6sQEosgct9Bh/GBqa
ghQDsSF5po6oJGZtcK5wlzVatxBlznkwOpS6NL1QYBvLtQSGcwgSWZSVLV3JmRw/
P1In4vw3AKuUVCNdQxYKFmOwKsOwZRI/dNWyRDDS12mqHaZ3VeP+o6bdOj+EMyzV
KVgTN1gpX9RVN/Q8/eKUH49uBroPW3iga1G6ir6cT80LZ08TkOMNrync2nFN2zpj
nnI8HJpdk0UF0aJMySnoEjXzqjRhBK3JTIB8MCekgRENCKrDdZRqrEo4Iv9T1JPW
SCK3dIsGfTcp7CSUpMH+q/doyUQlR5C+2Gg44Gu3qozmJ3DvRH1FE4axNgW2ZAMU
IHGzDSalc4DpmK05pNt3+qIFCCpQatxO1QFE4Rfh9fDeHuMGoGn88PKanZdsi5NY
OUnzJjRT+5DaJuLIz86RrNW5GmkotjHGhxlSd9DXYRQAMUmzTGltJUd9yNfaFfXO
cKcgVV11DFP5tEm2v2GoMQqdFQu7LYh8j8TBczA48JzVCHvmVTc9GlAMDIs0qCLb
Xt94nXZDhrNhw76DQ7LnXncfFP0RmdAU5s1hkA74pvWbizG1lCvUWSlVZwluEOTc
z9p01UNPIHHrGsFE5IVP/+bZpX9hQiUSeDz8TJhlro4mBOGoDU03lXJ4KYXhiAms
ThnUGHsKoUFxZcaodq34RHn8/vytq/JAmQM0vrgGprB1pciODgQYnyoBjihr4Ec/
xymE8yxDioVP38+mrkBCqo18oWpy/aQNke/JNd08V8voCAQUGLClONRiWXIrUnb9
tH6ozjSjJw1lwYDYqn6MUctOCMLk3ZWbdHOLOq3zXLnSsU8cT8KK1NS6TRo/HJJ8
oQEGoR7Y6OARqIjOhOHdfRy62gtf2d6ePIAuR1wdZXMUtBRxKbjR8NXmOXMlA38b
/uZ5MNr3VUKyp4RNSiZSovdYNRjRtbQfNRg/PrmslfhE/HNBewFnHq+j9J1ylpMT
YVbX2gHjKr8uiIRRJOYET+V0NJr2mh43jR0wfnnj1mRCo0XHiwmMkYnxciEUSG19
PMIXf+MX/T0yRyFkViU7Pz/yyWW4ngh4joT3Q89bXdPb2VhP/j4RrV1LjNuZdj0t
BE3bRCMox1tZ3MNv2oYWNFU68JzmT9GguUyD+4hF17lXTxqJUrnjGY6II2kAYcMp
giVpMAljAPo23IJk1rEgU6Dk8ptXrOWVaIBDYAhX+UYiYvOrFFnYeOibwJmY6nj2
/Rn35i1472wmdMJ6ANoQFvwlFQ97WYCVLmZ/H0y/T1KdeM7kxx5+577YWYS0O5Ba
v0Tg/VffKmN0yMW097xE4EKy41vAd4WZmPYxzJax49dQL0q1+yDfficioBA3xvnX
TTDEV6e7aD5D7Y74JobVLkRp0lpFszMoqZflRwyYs9eeMmSQ2CACXC+axBisA53v
GXqQ5HHAXgPq/SY0HmwTSkrrrVlPU+GAIu3SlRgFcx/E+yQOX+TVke4VOS0RmsE3
BZ3ao6YWHdPnDUJR7HIXDaWVA1KhhBtTkVkaEzhruQJ9ItMZolh4ECGFGMtPQDkl
xq3cCpPuuaRBHxPqBoP5x3ryCIWhs+wUY0ryjWx6HhjLakoBD8rPJqGYfM2DFw0H
5WqhkmZWrcngs4+7aIMLit+Rr0+7opZnFDltK5b66P0Mr1GGD0E4kj6f33RQaUq9
LLE3eNEduoVF50dxfZA6eYRMrGpfjfVfVk5cn/wvI9WOHNAik8VyjFoMxa/ttstC
/Q/KRiWZU+EiE3E77zKnr3OBngs0mNz3xz96/xW1c58X8GJ3Hw16m80gRzF3CYjo
JAuFXFJaigWFtZh+RokNROBVPmbMQxgdYXnsR4NKPQnOvohYarf85N8+9G5amvSy
Snw224InUP2K+/lDXTA4h/f0LMaQd0po8wsYuJ5z5sTvHs7/n6mZuTrIODWEtaXB
7NsQtoWlBej4wfvX+bzGDrHq8hkZNgyU/lsIY2zS0Pan868uP2XZYfpJMvZuLaR+
NH2hRm3QWcLrovum7M+TjPlhrDjrqRgzErrW50s1Wtxkwi/ycb1dxTG7DRWcdu3r
Jw17oOwgwO9r8D9ccBfYNSXVbXxaJbCssj0iEMSmVjb17aLqQLvyAwTIMxP+YwKi
72rF7EiM2nNdiSzLPzX5aYVNW62Kj+1BHAbVoQvrsSEqWgQ7o2IPEi18swXhXKwg
7NHzcVnYPuCCL7APR+w1AZMcpeiyBI5oMpeO8Lb+HaW4ujQwNwNAsVt3OvPmy2rY
z5RXA7fo4sUuyAOLIHIqFnHx5MctX34Kg1l3SPF3mHvxpMntd1OnoceSh9Gl8fAP
F7d1UaUuFwFArspF7kVClCKT4o1CWLDrt9p0PTpYsKQWE3SBHz1zAZdPvjOmod0r
TCA7a58e5eU8qNA+zsxfBJWZzFyq7SjoXrOc44LZKNQ7BJFtKQ4uIOjS5EeSs2so
qGqsZp+fOO58gnrDHdBklqQBCIOVw870EawhbMPPT7EDciVGnlQjQyXf/JiGBHHz
I2Zno1Qtp8T39w/qQ16H/RuNoRu9EPvKP8WRQ9PJQrqrMSlJ0IyAUz2y63clEZ/H
Fhchi3XXb2MCPLqs+XkudTZbxUewzzLQ3pbobkFfu/878+gyXrhN/HHpgp0AkXUf
4vX3hyGI4PuDsZtwEZORRFhJzST+SaaKjR2aadpQTIcewwa/12lefzFAsfCNjkG5
ztspiYL2NmVAkRfjDXbHfadURAb1jY7NxTnvY3gT5QE5e42yICEJ5A5WH1TI75Ea
5ipsMokqVeWAh9bfAWpwPe44jdnOeN9GM+pT8GvIxnKWGIpAl7IdEgJ6LHH81tht
E1XIjzDmzR103V2UpboBRDZweNwi8MLB6l+HBf28z5Q5db4yffYd4fdCiEPHOEL6
3o4AfHLJIK7FAvcjzTK0F6sybiwMijoQVe9NBpcvOY0PEA9FqzQD4Os+n5hHBrOe
3ECmXK2/nbbFaO9V6Lju2+TaGgq6/j/HDS/SHR1GATRx7jdi/NoOlhdsnFt5D/10
fcxho23dwXkTYnLwcv+7A6NROEGeJCylG7cHX08urUMe0OiRwQsd3gcpUGqfGLwC
dcI2FtXMR06GwGdjmZ5mg9NJaAWdt2QDelvtUp/nCldihkAx22e6mZca75G8MX5Y
ZvXfszINYHwBLQRFBUv+oHEx3864yDHSrosmpa/WCubWi8GkBlmMNzln9fhuyx0I
M+Tu/nL+fJvxsQ9filnWCN6I+Py9d+jzuB+3+XaOx0XKnOch7NrnSKDRg9ZTpIkS
qpBZh0ysfrfmB4ZHcJ076td4AHB6b8eKOVTmamraqjf+aIV8vuhl1jIFNXGeaefq
dzWLOJaN/rOg+apyjtoECgQw35WCzwYESiB0rMWLUx68KoijRbED85v9Wr7uHIfJ
Nn7CEpafUPqZqUny1GaZd2gV5d15/oM/1bPcdiZFpuomgptv0vWv3p9+JhUHKr7G
/vWC3JA4ESmD+KE0FTrMjqXBtsPwpbkr3+Z/xjr04ZQUO/UBlFzrNM6AlWubUe9f
0eHyo+LGvYVN3kj/nEcztM6ykhQBpwutQzaMd/+VJgPQTvAnX2E5+WRYodyL1uvu
8pMlqhakhXej5sQO8RlhfDoH/DQovCJIb5N5duaF8PaZnXv4YXZGUoSt3n/4U61z
XeeiFJXjj7rM7ay/kEOC1tUHkcMRKi9VMoCJASoTyI6NtVKlr8mmN1suflS09GIF
/7zy8iqXQ1Wq5YtKr/skox9beYySKOMUYA0aoO4fdIR/1Ey0SkpUIZCwTjJQIz0+
GeeKe664t5pfstnyTZZSLz8B5IupOmnyO0krpEM6Re4QhBVJBpYRtJ7AvVPOE713
Sn6zbF8u5aD25cKTmFneyPCoA7QUyhQV9GZptf4qGDsmTllHtbzisY7Brckesrop
vO9/bgdjt4zkVQhQy8S3nOBqilKxDp+8dihYDeFc5HbIX+XkrYFW96VrukXP73j+
r11OlGWGdaHzDfSE3IWaIaFiqGhzixRbe2F0JMhCYLgZKoDsgz+eKPbPk2Dce8dJ
eMMNH2QjlkxzYPNcG83wNBG/yC/dZVbyQ1BNouGhyBKcv9p8kWbtdn2MBPTBpmXM
C8PXUxeXe5qVMnWEMcV0jljW3t8FnbNkN5DwNAT2PqE+hiYOhTw0FX4jRpUpAHK9
HP4y1rkCDnIHAfCIwHzaoDk3dSh+USnJZk5iBuD6iMrK6eqvJM8QgPP48kdtWIx1
BEyDvtOXevXN8C3pwsoo58o0kTxyxUwjHAEsFeixub2fS6rv/vVQLY5hatiBm5F0
cwsDjL/zi0CeitHT/2DXl2alhvyjOWfts4u5AGf7wxvNBdiGFaJffdnKcoAuflyS
aSi4H2mdYpdHTSW05A8jZVd9R9rqSKxJ8dxamGRUbbWNiDFgoWuWakuQqg16mG98
kNFg1ItNC7BYg2QHxLRd/mzd6VrqMeQh7jUbMGjCiAGnwzBP5Q1zuh2o3G80IG2e
BIRMmd3I9pb2hD26ZGb50LTV7CKF/UT07fWZbdFfbsSehSrPcW3zkK2eTASiB7Hv
tOMuwwNoK4PU6yAXYbxk/d+rYEfmtGadetGqUGY4UMsuEJfwBRvpIqqU+nurxr5S
4mUMK/SwovbbwlFsAssl1Unx1IskB33H01dEoGKWoYLoZ0mZP9wSOlYg4pWobWPz
KkgfeWyuo2dBvHO0RoTZByW0y5OG1rkaOUREwntc096ZZk2EJPmYM4pLv/oRX4p3
uHVDVi+j6jFsFC5GOgaenDC83p00248hXhuRUp5g95pWQr5+wC3s9Vq7GtX6vcH3
6731RQextPy0f2kziFmOCvy/r9b0IHhVbPMSW8tGibpZyj3v98i8qNuB8PAvBMub
MwDDwb9j2H5TP1h3Am19QsOEL1B6tZ3wd/P5SOtuOYxxTvSoijPRUSY54sEOCPmc
qY37bsfwk818yn0DFEHbudEu7saKV9Kze7jOcjtsOABj/fbKT1Z6ryrJdkwPSn+m
BqK4DE06l6djRjc67nRFz4vl3xzjQGPHE2caVWUrLD+TsIQ69WdmEm1Dmv2MhbJW
VOpgDA6EprQk3SpoiDQQE300AMi37Rg/qIfSrkehtJVEbWM11jlMEyJwKIBxBDKr
TNgy22o5FUb9izxkMyU7RAKKzDcvvFcPWqet9uath0LO18YYVxCjcbx3BmZOZOSw
f6QJdYLWILVxHKF95UMWKgu/V9xKRiEW0ZUr73/wjSkxSXIe03k0kWl1Q5we3c+g
1NW0L/P8zCsZbNP9rzk+d1QLg1JW01c7q1b22JQpFGeMyMUbR7xWA+jwa+81hS9d
aVdpFKJzjDZn2BXX6zz5+ah61PccKvn9Kjwk+6lyUdH+5HlEJiju+wKbU76Ow393
syrx41VvrYlCteai/6SAR/VsqCvNQMgxj1LKEzYSGIw8w14g1yJmnVu8mpZoSRiY
CIUimSRyO9h8Z4Dwd4ygVwK0jRUzigzmgexzitr9r5K3w7OgRDtGUJbHIwkVb3Sy
+1fGufH7PzfIzK07VHrsd/FoP8JQ5WZvLpKMNVYCrjQ/wev+RoS/o2pxSMSMQQEj
hoifOQqgQ/ePhV2w+APqh991oY9zyGiDlccpzM6krdtw6vBhKmgXcMTVzpt2FdQQ
sdTKLSiZHSYj+v6NemNfXezVrdCZhr/jcumDVdzFglW0spzzEOCV+Ghhlcft9ZUl
krMGGSTK/qXYLF1AeNL03dbIyjoS84VFqNq8XzvHbMVKnO9/e2QdVSDWaOV7J+Lm
naM6zz/i861YSSAohdatzJdRDaWTijLxU/mzsNJjz+jCvwdOge+bPj+v9LqPNb9A
kKppavR9/3cR+9mgWsLMHTbN3X++CDgqSmGUzb5vB4fMGLYZuhil5Rn70JSmu1ez
txcvkzjC9QLB/qOmCsrGD1E6sy4tIFx56tk8DRDK8+VF/ecxZbX14reIULwxKN6R
JfTjgjD00P77J40q3etn8FXp6xGKoWmQGolaHb7GVUVnx7KJ4oC2gZJPAQDOVxBB
tmmzN2rHRbTzifno9JdVbrllDxASQDlmffUOv0R+MA93V5Y71Pqi3yrxRDtw6OXo
uUqnBXy2PbvUxNGcKSGNR3+PcxYmuE+X/34mTzkFgSmoEu5USyNGdzkbSY1no3sj
noUNTZ8WUkfS877qCPS/PANn/MVKSVP8sPGiD+/iWJtnMe9m+ZoFytWk+tyIwYqy
4hTl4IiDQvS3Ox2+cU1twKYlLo8/MzrKt79qqK0nZ6Rk6dCwkjeqY4dKBGVrOoQD
a1VtUgGjmiVsyeF0KWUib7VtqZfQ9iaQh8KXj9153Xf6Bv1pLUYdJ66kVzlI8f+I
O3l1i1NT7yjZt0iPN1sn2lnXUdTqsHgR3cPPVImXRyX5DP0YV7bHO/aYQzTjukl5
cmCfH3hDrVLVKy47OTbtgqTXRd9WwnP/CoKw8xEsoUHuIRLyrGC5fjgwEzLKCpq6
pga7h2G4ebnmFnCSNfpA4akMNFgk6/ethPMiZUbzysnXhDSFdk9LYyq2wXgRb6/5
xhEJwCsfHycxWY4snRWSdIcG+LJ3i2FbngzCw+Fnx9svGHWuNbTRwFK5uyoLQwsV
Cwqc6VEOSSUeWOonrGMhw+9GhdInMJ1CShJBFFk47cpy7rGyqKe9gLEL2KvNVCu5
wdF5mp+q2LFuYsYVGzkQh3Z18rg9nBCw/515V+4FMn1yPmSKnsIc3mSPX3isbUZu
MZzoNKLqIT6CkWGIqusBD6kwXJjStZbc0RhWTztgQAzo7VbDOYZNEawZv18f9Hi1
6g0L8DwCg9QFYkXWAMg7IOFKwu8Ow9SA8V88IYZG/cD3yAa4QeYtjSd+5HtT+HqP
Z5o+6cr1qyIWefDALphb/7G4hOpm3FsM2LWtVhlpAEknjNou6fER+gUIOlS0PjHl
K0Nav0jxVKf/Z8rbnvDixqEMViUMytdMQs/y0Cjzq6CWkyBZoW4OKnyMdXlVHeS2
lPDL1he7b5annH85ct5RXqFtEY91zzYaxx5hILxhO8VfNVZJ3OyJwPTiRDAt4ZqB
TC8J5qbXNFHusx4xNtiHf2TJDD0Hkm5ojtd6gfc76FCWjVufcwtnaDw3uvhJ/eVX
CR3oSs5VMlOkjcXFCnIoqDDLpwfci2xOTlO+zEREwTDcD0oZ4PZYV+6C1Euczuhz
ufaw0bl7HGNj+qHmIFpkZwkcxjRFKNLC0C+H5AruKF7SLCIvxrTPPoyF81MPslUr
6okVCcRDYxL3qlLUV8EvEsW+BXh2U4UuxnGRBrHLOQPrndDg/VelyKbfSYzDwKh6
bqlhtMzBlyfag4brry8hoBDVeWpMjceXWeR2UGoHv5VqWBd8sm8b6eEolhWVMe4R
lh3dqxCBA2NeYatS+/Qi8Gx6q2EpORAIBXWr7HyWKJ00NbmcVGvxTEexyIgrXZfU
x5in8NVDZrm9mA3IH5yFk7efLnRgyjSC8QxyNanifN9xt0PU6wX8COeofNS9azbx
6yHEs1H3W11brEOkMAp/lhIRvmTkS50k5X0bXNmUiU5r2D0CaLcfZql44l2Yd26Q
t8h/lhwtmY0vmqs8ry4Nox+IvSzO+xwzYcEjuusbvF5tXmatSWkgbGKdzM2MCvdR
X9Ou62luQALOmIO4jFheYbtQilonXpWnfhL50HrBwkPUOf/RVn3chGyaWDSUprwC
Bw+IK6gfUoYfFv6prXTjUK2Y11s0NHbzvTgQSM8RlfrxYYUXDQUGkBZrXi4IpJLL
P7ndTF54qqt3miVT4CbwY1+CDQpIQrcfqRiTjm7ec1mObC+1rGBFJTctb3Ut8U4y
OOeu/dHCy18dGyauuoMoUxKjfk5UTH8JgTeV+u7OKZPCoSwrrBf4oFytp6d5R6Xw
7QiNliy5Lbvjc6vaiMvCVtR8t3rpQmhBDbkCrwwoh0zQ0J6rRdxmeXsSK/5KymIA
Q1i0qWmoG7DUMpmaxUe65tGRyf0TYrlydVcC8fM8iYv/hciTZy8lOIlx+6bSM/o2
vOjnZb5szZEedu8PMaXWUVAssOKg66fV773o0p1ScrJ/MMETuO3yrN3D69uC4bAz
gnZ9WUg+3KtV6PNytodJA3fGTBb9NO5xdnwAdvDeyFu9ruPYHgqlYz+KDSXT3Owa
+/gnYz/ETFzhjeOENGomO4E4ALbYpVAzGnDQ1tcqJ8RAHWQAlsg4LP+As/7jtMKS
1nDELAf0PL8dETnALmagKAegr/fqWuJKMXyUKQbEf3IJV/PSWVBn2m24O6L/5Mnk
k6KusAZNEw9PMjUq7iq00KiJnqemA8pEsSpqbG8fW56WVIydODxQQMUdm48RFfLD
eZx85Z2p+axghNS/0iplLsWdQ6DDJ7UAUKWc26BU+iX3kmD0T4SgumsENEYxHigv
kWfIMcw8ASKWnT1rJQ1NSF14zCndL6fMtxF52Z/6jCb8yK6FsSWNY6xRIoHhIRy/
WByV6a4mgKtU58cXcWwDM5/OFSeGpUrvrsOHZY3EUr+orpDXlJmJT7KEdWPWKEqf
NmczOv8QdvZTYgsbfaecox+jpAH01Gwb8aLKe+zpV3bpnhHSQ9xOBBNd4kQR8EZi
o4FT07WemblxmvVdVc1kPqN5NPktQz4QRHU6F69BWBnQGK/rs/f1bkxIXbS4n35N
7kKCcqvPnTfRR5a3JDE1744E5xSDw6wueMah4PkGQtCpD+hTa5usvBvghlkOZjyN
x+bIHFgXpRxjBffDRVJk+xIkGkDsz1STXV3tz+Xa+mYLcUfv+5f8e4/ZjMDLBMHr
iSHUlWuw19iUlzvo+5r0wSsJWBIF3DuxhJhsi6oksdV89aKnifOjqZu4PmxkPERv
YuLmq7LYjJ5V7S4c9JKr4nsDUEUgzqjt1c6MqpU1ev4n8VfbGnjQ8RhfIYDNmSXc
OE6mbu3BFzc7ajfuBzy9iiIaeGqTGyLZV4XCMA/+uXbWmadjHiaych6eGRLRyXTA
OyfTpQqGiv25HmIJjdJUMy4KVsqE2QvEdM3guSaJRm7f21gefAL77Utbf8n7L3fZ
KAKtat1erUYU5NrWYqNYdzts0PkdcCKlmditu+4mUN4kZwMi2kauvkWi59G3i2a7
2Sqr8BkBqxSttfoBOsupRVthhRdxHyxw8nM0H4HWR06tzX3uxIiNtCjyVUL2PW/3
oJf4+As3IR5HhBmsvFGgogLeMan4ngEIz91lHYXQGMWSWantajbPjkvB5TKM0dww
MGfZMzcmDrqJDUjXhcZMVyK90F5kKCQdokxl3ZZIrpmCUiZl8jnkY7sbKKaiA+iF
ECNi/sj7iX5YnJe7eFbCN/8W8cV0T5K/6skJbKKmTTXsh2yddu81gTVXWtuYQI2U
s48bATpKf4ttZlW52/W9Z/Kk8ZsX8vz2lMaQunNmIDvfYleKGJQBDrnGovu1Fc+s
IZQzJM1CIkp4JN62ALKPdOoQ6DEYYjsaTSeNZWibDqNjamRRdgs3VraWtJJ/DBmq
tnUQ2KiT4POGl68SIJlpwk8zaVJErzfNdJNHMOQdd6A7OKMeiUUMiOGI54UiR+S2
Ap2k3kEledGtiiSsXjbe1OBeKruu80GKmEByjnV971wF13Qz3xzX20FahSXzrkBR
9cHKriYZlROE0RONp7TpSbO48XPXQPFwaSTaw0vm1SnJM8VdLZ4yn5VetKUjVsSb
gNXAJaa2Qwq1wu/gBndKYB7GwOl48/q3cT0knR+FgPN80LkzPIFdIPqEutSKyIzB
tK4g+T/sJH4UmhstcY4IK/WRBsVd/unIXn5JB7phE/Ms2EEpGX8De+4cYacOyL9s
P95SO0DHxOZPuqFnTp6qj+O3uWXu2KFzsXfSzuLUhdyspqQ+KoPvewmdyY/2EM92
ZoSmI3ir4CiBMU0gubIWEu17qvlmdP/5XZdK5Lq3bwfXjzj80vmTZ46fGtkN411U
Fl441wm0JG9PzTXfS9hu8wFDmARRpcit/kGyKud/j27JMJEVviDRZ1AxO8iRBKOY
Hj+iXKPp6BWTBxt1gtD926TueH+/wKKYq2Mq2nrWomD51t0+bU2bCbJIvOlaMUTZ
hLEZVI3YvSweZ/zFOIAN3xlBo+a/zyOkECb/UgUfrrgEw1rFHbFXu6CRc7q8Fm7b
3WjEEFx+Go+SqxAkM3DIsTVYoynctZEI0FVjfsOQuFrv3WtWiW5C6IS2DJPfw9Mz
N3/QIGxCV4E3QckSp9nUsXfYZSjpQfyZyLPb41v3OeYZSXRU31T1o/Au08sH1tF4
377OTGx+JsSM/pZ3jHcGfXLf3n7S/4m0lhNWkd7HbroBMync7BZ6Aw/Eah6FE9WG
zueWdTVqgYjW3z9HaVSLxUgRT0kw0+GzG3aotI642Zsel2tRkdIR4LovoOCkPmTM
qhynprD1p9yaI5tnj3E/+r8TbAH8BzP/R9l9mjepwXbJM9B7LFTYrH1b8O9x94+N
ajwK3WnfBKd1YjYTqzmI3LzjzATc8VpO5thGCuYLDpeRcJtHffzqvn934HuZuiM4
7xgiYXD+L5DepqO59PIdbDdCwTK9nm/S2wcKiuIkOfTZpI9GTSvCr/mO1HwNvMDg
QLFeQ9acBdkYOwhnLPoEl51sIPkKukil4enX2rOLepQvGOYnA9KS/3ELWx4Ppd6x
87yAbpQnRXu3fnTZdmUL+ycwZfm0WaS0SVP/9D+oiRjT6r3IEvKFOCXwLW8rg3yu
WiEw6M32gQyIzfq0Y7DlVZnc85Q3fGqhnwlM57iugf7eIBMrxcn5kgPukbSjJ6hO
C/C83gie0Mp0FxVywm7f7i0/iV8cDfuQMautBTBXMQVmtDCQp6f+PuPOnIZ2wNLr
KjJ4KKNs4MU87Zir8FH60gcYn4M6lEvbuIVZPdQ7BFL1C+1fZEC1Q1wyWxHMdlQd
e9ZNpHC8ohWNkO0umw4N+Eg25A6xIYJY3ODfZnaUInmNeptnqHVd2iRYoDjtW32R
2BurZJVXxs3wUr2TgtwBvrOy8nrb+XCEZxcfNkOS53PXafKMCKGzfXyJgkiheR1o
lomA8TA5HJcv5qOYK6rRCXnVD9i5erxsDDbHhbwl4UeEZp+3n3ag3o3iNRablPuL
ltN/eV01JEBcFlp525Up+gi63zwfV6HZGMlytfbK+5iAx/G0IqhTG4EQzhXB6vi7
qR5+Z4/+fqFEVYn8GjItnW/GqYxs1aos5qfdEaWS492tZOxFmCUjWrtwTD51CC//
1H5xr4YKfhxvwhIT/5mBjSE/easPVv6L5ROmF+tGKk46XFgjj1grtktg8fW9uoYt
QEbBXVFmZIyr2kY5wTwRHKDjOEyxMzhWeAtUeIA/3lMtWpYfAd60efhuMeAt3cC/
flfGVoZVlbsCxycXnDyIcCd2UjeEJxsHnGI1F6ShjsJS5OrNZiFNte50Pu3pCFHp
ibajUpGTuUO5Ovjjhzm+1/1AyFS58dJtZzMCyrdDIgxeZiEUdJUtZVr4tx20+zBR
W1mYgz3zVxWvKVU9m/LRNVY8eCFwLCU7QKmoh5ZYGorfBDFIygkEeHOQRk+Ze4+S
bBCmOn/sShpy3Jd4HkR2qqi/bZ2fWt1SjYQMmvnPW8RZMuA3XqU2YyRniU4VpWnQ
uT9hc83aJ8pCGuuAMV4KUXH1/q+j1lnofCbEvjJ1TvR1OgnBqLDaaVNF4SGnHe1a
Dy1dNXUF/CFRouNADEpegDOqCXdCN01SZh1lmHCcLC5V0oL8Qst+NYBa141wRRUk
6q2Q05wRM9jcDuCRO8I4Vg82cDBKE/WFs1teWOGgBDy/DgER5Rgf6iUNFT8h3vNG
ZwyKoCJpas6iE9s7MT3Fn0yk9qEkHCBpdbUSBLp5u9HwKMenGVU7XZO+4Y6uVj5V
XeTIMI3ECQxmjNJlRpcwzhQCzyES1CuCXat6t1Mue29Rk7mr5Q1HoanVkvGIfb3Q
n4+XwxoU5Xt3cLj3qIwonxXNMpemHviZxnXOOoPAL5vBUOe9QxEWawpJCdssIdvr
vN7ctbMR2bo6cz5oxRBRR/n/BerOZZaINWNXdQk9pdMe2V5v5uFgwV6z6pfc9T78
X/IHqHF2LFiGF+ykwaalFeSanzroyjF+gLIY6nK3Wt1e64MxsP6VEvnglUoJdDaN
EnG6oLN4efFWemyCUPIzf9HFvfJGO2LxJ1kJ+8qTLTCAFLonwQl6D46VrgPni8y6
CLIecdzTBcJgsnnSw5D56RkQC0BndJZXJ5cYeT2XJZp63mZ8YdR0aHHiM3czj+Zv
X9Nnq7Fsl0XCW8nyWDe6nxP++P/D2nVMQrsKTLKcRC/E4sWL50fXMznDMMxwf0eX
P0hMrzInnwGC7xE3mT8pccQH2VawEMn2dRLwBN02ytHbXeUTQGfBYaLWRGs+C9+z
SkijFREaoDt/ac1DVxogH2SegjOFJVmQ/lBnrj+mSIS9PztBUyRrlObDPQGJn7XX
DA0ItANoDoEoA+w607EAx44SLZA7EK3kYlnEkSfanJ7eol85cx7GIrpu+tJF/6ZU
EFwpHm1oRwIjGK0doy+QlvVD0N3tuLDyRRgYfaa9XnEQY3yvEb/Y2RfO/Ew6u/RU
OF9Vra7yXaGemX2mDSRYpuEAFRi1+XOiD2DkYa9W06xBl0bnzcEkm8Cel8t/IEHX
Ks5ZlYRrQ7uRIYSTzF9KjgUXWqouDQ3G5j1Rz96GtoQhXQTAfgo40urD5rufhqSO
Rch1vu5TebtRimf4eLUGXv3aDaMsbcwaORhJ6TanLIW69FHJIlKl0oZjJlnFSW+/
nguwN7Yi0Knd6WH4fqZPhxpxzxhyQzfsgEv/h+ypH/vF+c6slYW6w8Ou0fL+WQh8
jfsCgWl02BeMHRs/oGU+R+ewKZjScwdduXonnC0LMQX+LjY2stzIueKZnq/xeb/n
Z9Lc9qlrhRUZJAepa3fPrXNdyNlMFKlLp4tLy/RlQUBMiKGXbYQs+AmjNAe9oOea
V5PKlHlG2F1YqQrsDtkoAUkxxCIz4l0O5qDpkLbO/K2Twe6IKZaPSDCc9APEPfVH
UybOPNLEC2Je9VcxCNWNEBiZV9fDFF+9E0k03CszrX4WMUuQzzsnyM7CTWUwCJOJ
35bsuJheMSvQWYkyY5ojTzVndaRGKpzOYi9ejA/FPeTEEuVXAhQiYCpoq2FPzDRX
M3JWr4qH2B9CisGnh0EEj0tSamBz6mKRmwe0OdZXM+SKxw4PGcQP1f+G91AeVyaT
3gOivu2p0z16X4GXt9kDuGVyUr9VQgCBlwXKmt4ffhBItpwx1/jEJaSvxxr1M6Ao
1L6b2AqMeRj5O7WHnTdOa016QaFTbgFhIm1MVRQ0PX22F7tLp7DGGkswd9Iyn86t
BoqOZ0p9L969ntCDRhY6tjxZcWDZSXzQ9ArWAKRHqAtEo4Ubapg/O+EU+MX3/RI/
7aIRk+EkwvXMtSbFbfjbyISL6jOsarEti3lvfSkkQIVeMxAqY7L1CL0nWvVs6+kf
84/G9MRbvffxd6DSTKkiroB3XaUNJKAviUCHQFp+pqcAN8Bff5hcS/rwf9ISgiSK
DtujSyeLYGyaqKznmBODA1NsPJ6czRb3Ibn7HdwwMhjBhWTFTV9T3tYuzFc7vhJo
Wsls+kStyHR4pHMqaJs/xQLn/BpiFb6x6sjx6MOIdBqX6VIvokCYsY48cOnhJODt
gvl3gZ7AcqRJRrgc+C3JiM9INsxbVomjVw4OMRc4rWxsgQ6zZcfrufvT1i/LQn0P
llMiN77YAEht8ncf6ehcFf5wOuWh28SoiNyREwLYOtR5W5NKQXUHi3LAevpwyj+U
GN8jpW3fWlLAMBZ6PfTpSWA49TEZZQM2/9j2d8qROy/1PhzNeHDmK+oKWzksrLCh
baARfJRGaCGp4bE5hrK8EBdh84Qp21kn9qMkSF88M9rjCu2DmsXRh3yOlkWpe4HR
D6sf6vChAQR1Mw6jNP6Gaj1N+4Qj6ALsp8SqgxRc+AeEmOGQlHxRU9dbWUaxQbdw
H7mFgrDdziAIM1pEDWlyXTFy3hDwKhpMcMRa6Y4O3+bNqs1hJJEEytov4saBRnNv
im/X5YXlPKzzNGU7+EufxnvCFgCuqtcJBkqY7kkcu1FNArF4fmMrpRAIywD4e5Mu
t6te3ZfE4T9AR7MWTE51hFRymruwqbbxJgf2NPME+/ZVzxq03nyN1WkGCWIkGpwy
4DBuWQjhlkBiCwVA1VYAyPAlCBPj2qZcfYqYV6IJE/JghhVL9Ct6v72Jit2eYyeL
/yZ3lOXmVpw81D6XuVW8M7iT22ZyH9JuerXOvPpj+8VJRCClYCpFKuQX31iBU9NF
VBYRxr+uDH22zzS9UvDTBan5AiBQ5zmIXMiVGLEkCvSZ7Pzc/TlK4oAIbLu6z9i2
DBUQEfDnSL8Z7wHsW/KeIJ8eSAM/bf5G6JD4Aa/TyHmb3rcAKgS6j6JUfYJI/Jru
XUpWzZND+hY9gnLF7HAhOK4DjmwI71ku8/rAqDzh2NlyZQoYwCpW62K69XhAOFlq
epmiiChQWBfwYPdrfv9Y9BlkGH1M8hB7CWK03k5Unq9T2BcxnPYS+vKkCMLB/v4T
Y8vRQZwECb0x7DH5EQ5r9W+4Tpjecvv3KN8LCxZF3G/Rb3AdP/u8ezFbvgYz4sBn
F+2qaf/7uuJlgoXH70fkHBD0XXP54w8mo4JQJeTmHVIBrwvUVx5F+6XKXC7G0iN7
K9gLehltpMZOhZ+BVamEa0DyANL/Oui0A9uNETIUf8fUJa+6PrBWao3cgrzmj3vu
YR8cHUNrcUmIDWKcR//BUU2wjqt8RN5iyxZyoepqvyHaSo8ezsNdDHn1OaSYVs8X
dbrVJ2m3UyyyPWjZDdzLxfjtWT8YRqPdYLNfYo13AUtlM20nWP0XCLyvGve3g1V6
CGZn2/w/gi5NoLDmfIbJEXu2VIba/LzyW+mCj73MXsrJSejejbozIm74NDXfrnbq
725rTYI7keLR+h5ars6EZ/hSDVyJPgOXB6tpiLHJAq1SwHHN4zFHnd4CJMiGfJem
k2m5otV7rBnKx98Ofga0c3T/6/vE7TvHyKEPjBj/q8GMAsIbhBuyq/7W2kpyl8SK
+m1XfxiLU4ku1ETQWhhWsKVcLQddnZOV+eg5nBkLSpD43e2ezKnO2iOvwxkvA13V
jiZrFo4RKP7n/CbLZEh4ALmfdjjCTUEtegFl0F4m+o9MeyDjofDp2v/52atf/WOC
gxLQJ8Lbv6hwHizwvvW2kzFdhoX7aUbUwxu+zqShA91G7mbk3V+YxHpwQSVZG1a/
tXmdGdN/DLXYT0Mz4xSPYPfoYTYU5p+CkECHAE+cdHqKldRzHvJethWEJFBgj/W3
J/gSgTOzhIytv91Hn27m5mLxgVsx54J4itjSzZN3G+ZjVAjg2IS3dEJ8DFK5Jumm
8s7vLy1f75IpnTkVQAg4avNnxYH1lnK5jZdr1QdZQcD9JJ28Ds7Fr1Voha5197Ac
qxMooXqCzt0PYOYBZO8iAZ8tcIfYGc2CdpNajfmtxIfjO2J5w4hOxMe2IowKoLct
O96V39AM3iGIv1hSXcJ5sHRh4NM4pydEUJv57DP+YCzKUWXnGmT21SHd4rhVaKqc
hD5ezPywnApU/mEUTVN7Du9qG4ewS7rGUBitG5aGfiPcV3sKmz97o1fhMxtjZtdN
3Ap3l/O/5wWCFuEQ9OH3FMNh3gRuigR70HvLrlTe5xwuuznbcilkKVJLiPCuY5nF
Fp/wa5EAPdNUzb7O+VzJ1lAVEDWhExlGVe5MlDdjCac0CEg0pD76EPsBfbWrH1WZ
gtX3sJnMwjehXRfZ+kZ0vYMx8EhQWwlYFf/W4xI0BhYT7ja1BxGXZbv7VrCk260S
dtfSZVXNlhtdnjjqFtQAqrZUfNdl6wQ1s5Xd0FvsKcQoMWNjQGtbeVzNHaS2B/FF
OCP8jOU7JvTC0TcsFfCiramKsiRpDCE8mqPBLZSX6RZgZm4aBCyMaqyax3WKttNB
ztHmPtvZBJf3v36RmGICh4JuPGmdB79t6lcP2mPRiclAfUNkrLEONToBcqTZM8nk
tOAqQKpi1djzBd8P59S4f9X8cFG/tdOaSGmm1ahN0lx7lPD5zMi07SvQSGXs0K6X
K1+LEK7AJtjPSUcjB4FqOehPDPK0sgRjwt8dx6Z+FDi3FAULnRMHrHnr2V0b/hJP
1KIXXtVKaRPlUdAtw9wjr2YUeLqma5ngJJO0dSqMNqgP30W5VZ99BS1z05Kb06yb
gsa+uCb3lzX//hl3aKE0Y5Z1ilvqOFFdY49pQ/IWRY+rbtyBdoQY8YgoGiFPOqZw
SHXnvB3iRedvUzyWb2MLmvcoMXofqtX6F/x5nSGSPoiOoBh83nv8Nkjz72DbFUxO
6jdR0iib3ZNF7Or9uaVx42suN8PUgPyQ3xumNE9o12aySzq70Zm6+hoyJT5r/1a7
oLev2FLgVTlrRXA3PfVGVnD2AupBO9sdW5/43kd4PxMNoSwpMkKWJkB9rjHktTop
lrFpbbhrhY2AnAbpFnpjzlyVKt3wgdScbHc4yMUaprOW40BGxTjMhEEtVhca7/eq
qXsW52DP/bUuYlnlj+2p3tVCrkrPHLZ0HZWeCXh1eQgaE/sX3/7IgPujyQRtQRDc
AqujydSv2gxdGoCFBoZBymPOYAgvcHzGbomQDxzht7c5VkVHqy3Nsilx709or3Rp
E+gafrYUt0FekYDlOyKccO0NLBQclNUWqUIvyzCi9Rw59YXcbe5CM37WgorgreV3
89ejo2PbubnZ8FYOBPxNenweYnkURm/JJVOoQWJOZyPQgIVHhktknKreE12SKetu
Eg8ueGZCRdKG1jjVG9vx3P9fW2ccFC1IiFwMvsKt+xEptJ1kKdqNU2KivBDcxibO
7tPIB7tSQ8ChSH+CJCGwoZ0a3PlDFXvz9N8cSayB9gguTW9DYrtc5z1m2yUJTvzG
BuobYnbs9ZuHiVLQe3jR2nP7JjT5QJ6d6IFRk/ZqFxYXgZaZSGge8OXDC/Of0HCT
dEBVjk0qB2/JCnMq2hevpewq7i2UiOEIKypru2U1KqhfhhR3OPFaeZ5a+p4iLGo9
G1Qlxi95ILHj3oHPG1rcmXVNikLHQTIIfRZ9aGBbDLljAZ7MzSPvp8LzM5UDeLhc
oZ0Is8+NikgD7s0t76TMyekUcc3XW+9gH4kf1Ie80CLkS8uvmc2PHwZpItGxPKGU
vIleG3f1a8oaedAuOvHtRTKn5aLlwdczAMQ+yv4oxPvK1XZxp8wZt9PvZMZJwEa0
RqEbcaJmqiAgkd0JEDAk4XqZbS5kug7im1WuZKURKd0lAv1Nx3VpA+om4bKRZiiG
GXcT8ZdxI76JUlxH4NoNPD6a8Xa6NSarZWQxEKFlGHrzgEfQKPcjox5oXvK2ARHl
hdI7oLCxPVtUKPKkBdPz2y1jwAl/irF/QvFWAGrD2dI4KgQvoH81X14GgV5bW57G
kJT935x6i2TjMXyO/ZrjBSNaCtjSiFSFSzype3aREDyoWM6eWniEH8iXJcU/rXoH
RDHFramFIZzy+0qQzpS9Kx9M0aIvJQzU/kuYSfLu1NwqUH/aN5IO8QmqxbvtkFuZ
8wA1cMTeh1539DPE0/4paIo10DKzWNNer9vZFZONgM5hd4ctlMdxi93L9xcQEtib
XzSAEc3Bo4Em35H8v4YOt6jmsn9GF/lxS2qD3U4McGLCEtTplzD6567skhrclQKv
K1ajgoMDIB5hRq60ijWy8/HjHPzDAeSK2n1Vm1IYTxPxHtZNR27CuajYMdEGSzM+
FxhFH1+kiAvk/S0BUPIslj1Z5ayKnh2Iaf2Dpa4yPuVEVrheYQyy1lXCGnMVUAtG
vjeOoAs4HM+mfOA9thvXfnb354toUxpv1ChkI4Ox04zlfJLzvxYbVk0HTNWw+nRm
+rjjIIRDo12bQAynJlA+hXNnmV1m2lQKssOsYKX/L/aBJ7W2ehCLJ5bU38a33HsH
l0wZx6tO0XyMFGhkYbU6cgXh4Et6yq2TJOJrVZ2PCmRvJYccg3Rsh56OBCLOAnT7
DV4K/Z18WwInh1kYQXlQyVSGn1bYzqNJVkEy6DkvRoorLBrV9CjyArFeYgzYQopH
lceWg8pulayIH9Q1noJEvHv4uscDkM6PA4M9Lgn3HuK1VV5pCVfc06OBA8HEsi5F
cGo3RmFGOZBNE5ewdHwcGTj4ftrb2poG46nhEALFb8Q0W5lHCSnZqGky7WH/JKM+
6iFfVaW8amrlVEhZDPjXrR5QqgtjpVumn/jFB7/jnbwLbQttLOq52fYghCdJO6Tg
SOuMGj2d9q+o2V3Y3sccyKLCxzkswp/V8EMAMH9J49lQfrN0dC3IhIawLdLjEGd0
TfQMBWCZRGZp03wvn3REQzAWfE6mfqJaX3i2ebj3rntYrw0PwYGZ4VJQbxMilaMu
zdF5a3d10/1+FwBxm3gHNBgaRsCH6Ed6uN5/V0j5nuyJ6rCD/cSMuGvkIgaLH6TY
CRA2dIFZMWECk8TN/8UHSLiaqu+LzD3DODaE94OiFc1FjM8oA6lktnENEaK2zAuY
smTpLFYFJ2Qyvpjg8CixTKuwsCnwEz/2hVqvRbN0rqw=

`pragma protect end_protected
