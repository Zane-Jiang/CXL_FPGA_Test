// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gaXJ6TLcF3UD3ABRaGilQMdSzHB+u2Z3qunDXEvjl2LJRVAek9PjyZlHKs5V
Un1tp0MCEPkvFKV/XbSEeJ/e3GC6GZOQj/ZJCjFKgBjCqqHuFEaQLnikEX07
p5VYVs3xAaJW3ed7gUHGTbroIjFrmtGkWOgg2cmfHAvaDBqbwC0hh3xaq0zS
ZvO0kB7L6wYjMZshW08QiWlhe6J5DRencI1zyhiy0wgZoEnI2zayGjaj6s0f
nquojzS/OL5KCTDEj4kwd+WwaLbsoClSqTK4JCF2eCLJ6oo8zd3o/cFGjSkw
RkO95R/fZ5/G4xwCLRn8oVRnj9LcU/GdYmIKsYLRiA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E+0EQF/ThvUFC4bX5z8hlGq4Z78x0zto3j8GctqxzTz+urAeurDJCc1SqL4s
EGrxek3718UvqBPH0mKXqAVGqBHdcII2Kp2mWyuykorXYg1SC+N6BLRBNPaW
hTK4MI1X3Drya+7xieLrih3Qy1wHTKgBcmLfLhTvdo7/bmErV5d0gGlQCDc/
HKYj1spANmqmQ6FNIeHKkuRyNiaozil7yCQo/9VHLaTCNm8gp4+dp0lnKjTH
IOz0jom9gJUnwIx9sHTwRI4yTbaZFuHblk7iQ/2KazcWauYnU/oS131WLHj5
r+EEb0i2EUhaJq/itcKys+xlaXB0w4+dpEo7JDVSBQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RNsWdM480cUuhdbx7sWzqeVo81tGvjmdiIlT1u/WjNVKloiD+hCT1OGXFWAq
Yv6NPNAzapCDOOi5vo5U0Lr0jRpDyJ8Qg23xtAPdXZjl7yg3X3qDknKK9rOX
wJ7p4KWDrb5clPe7EvlB8PYdHX0QIkCJ5tIUhLfSxwLGKoIC4R0P6jRKIin+
hADm4J1i5xjxrunXe9bKsBkWquKueVlSWKfL8BCW7NUTbwmAkhyTBBHseQvv
D8E2tWbsPFt3YdT50TwyR5BfmWgFFmYLjMP27+d30118mxg757e7mSqy28eh
O+tPlOwulsI3p9hMaUpQh9EkPWc9QVBTd+j9kBIfiA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XAa5m0s1eWzGDVdXDDza33yyKUMoRqW2x35I0EMuOFnj3y/ycmusaPCBMuFa
3JZqKiQ4jYcsQe/NY5taHe13sjBfAKiActGCG8zVSbYdrGC6SVzRo8V0AmWQ
4J2ppuD6pOYMCzTzvP+YJidKryDA1oWSGS+xQdIKOx2LJzAEcxk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GV8z+jW6PQisDoYfINWH/GYQdo4mTF0ybYHHIMmXaw/PVj2tZyRV6cm7a8yF
JrbajNfuCRN2Oaq/FrtW1M0hDNuD1SRpEUohwuNCqM7d594ALLZAP5hiM/vr
DsZ4YUXcsn/kayCIsSG15s7qwCyZ4DBgz+IjZPreBwPciX/wgEdBNzTEMqQF
5Tyzl7c7iQQkCi6+uLXo3p4HqV46SQ7eL+taJBhSwnLR3PscolMVMZCAMQXK
+8tv6N7k09+H8A7KFmJ26gp+cekE/e3+/7sbg5/RbYkp+4/AFSmCHA+LVJGs
cV3/x2yGN8hgUQYRDmTTHK9iFAmg0IGOHs6IT9pwtVtnAExTqPj9gwYbdW5I
djKAVH97YZKRuyhW0h7ycwFUPfmSJ6KfOuQFGJ7Z+qldNnazl8nqh0v9XQzZ
R1eYTTCaJLPxDsLaHxFqqdFrXmbRwNsh108+b+E4dTMTidQ2SNeJViDig1fN
nV7NuwmSHQXa1d+EZaUiyxyZiJn4IR31


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FWe4+7K8lU3vsMwZdXaAsovpnAdzPx7MQnqkSgtSDLEs3xtcclo0HyDa6l4h
7xNGjXY32vWixcXalDEdj85+u/IGpCssiquDy7uZLxBFD+Xhjug4AgCW6AFY
AHOBWIlA3eBYuKLCjXeUQXJSanlHRyHAHe9+QN6RFcMrgN3xplw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ASt1ce8NIMbaWcASYgJ31njKlPTDLGEdM0LyhlPvE438FSvpPKlq0Oy/Cu6Q
o3JJKuR9bI41qaJdXY/7qG/TRkuZ2yZgQzMxSgLzlxnDu99uTkEIp75lzojz
hvJlfDX6HndNwglPxxtw6pRAYCL+cLXipfs44Pa+GexLPKLPFr4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2320)
`pragma protect data_block
mIvyoRoNlJ7KFT1eofLlb2C4v9aDcK91E3vhE4DFYuC8b3TUIJWDJabR7Vzs
nF+m3FdGbGeAmUZXkygxVPpuANLlUpfLDAGKyfCfwtRhQkIguZkaxDaW6izV
v8Gb3IcQkVtPoD6cVcM9SLXPME+4w/cv5qXtAg6ZVhDD8ASPcZsKJ+U7A6f5
Ymid/1RsupuQm1OvWdI8v/N0OruruEG5bzjCtSgVYWniyquHO96Ldz2ZOYwj
8+1akVEDoU55eo+6/wTLvr6O6MeCiU17sYnn/MrMWThvANgd59hpk6ldEhp4
or9IxH40sagth2HOrTYBa5Xx/ISSqUmgF9Sc1ev1wZNCmhkAdf0VmN6hU2Da
x80OyW+4hEWt4aideF9hlUp4ejNnyxZH54D4mgQ4TFe1CNiLMHIH47cplQx+
G+mcpsms/EqaJJXyCKw08QGIkRO/rM/9Ta0jTxqDqd4ignrJiB5qcPaP//ki
ZaUAoWcKM788C2KIo7SELu/HRfdfMlgwR3ll5XajvsaL0w7VOWA/g2kjp/lK
ULNPlr6XiBmKt9ShAzIORTNKUjcYQVwdkEmGoOxGe9Bz+IQSNjlz8YJOQLGG
u8Xa0++OfCNwNLphCMUmOzMuYilZ3ZrBe9NfrzNkJcmoGVuez6llCnQ07/H2
3LqAzjCs8fjNpQUxaMzCZzgD0z7Ng8BFATxRfD80j4I4yllb12q4lUZmnjMI
rjLMaNXrRuwsKfc1QXSWuX6CMY9TKquYUHyNBYKT0k8aloDcA/aHFLOxgxTI
UPhZQjO2Sa7xnLqAkcbHpgPvUoyxu/V90WgVIknk3nJcKEBYxFw46IF/6J/4
H8raBdFqmnccKqsUlTmNBPlfhgBUB+y1m2IwCBxj1mlXmqtrOQ9bHyhIwpA2
jior6jAU9ren74fjwxAuBvQzQdqfTAOPFg+fGzxLPOc7PyIV6cPGkhLPpAW1
n4sM4TyrfP4AP2BJzgQJWEEOEptORTgRlrf+I7bKC9kaAQE3JgYfEemd89nH
xW47qXMLXRaZXkyAMzlv/WMsdA71Ox2qT6K5wmfwxeCp3Df2kvJn+H+GFb3d
R1hJbH9QSoSwtfGopMkwkAWrTQ6XDpZyk63Qj84M/VeDOJk3bA3BYdfFaRfj
mzOtc31iqJBSldw4yXYt5zx+tipEvUBhoFbzDEXgiUJqxJBHY/iutdkY21ly
OY5vMy/QdidUVeRjBd2i3ut1C/jYZaf3+uzOi1n6oiyUpsJcsFq3afh8KBDF
lLR9ALa+4Gk14440uJWxW46OyuJB1N9M/497oD/uok7+fFzwEnuPucSX2VQ5
icDqwqkQqKqRx0o1xUoc5lhrn4QaKNXHABRSkMqUerd8cqs1ODTTrJj9DkSw
kPjBVsaEwSup3jlhU7xTy4bL1WA9j+lpLVSIgSosgKFANKHns/EnD0sQ3z4a
DoI/y0IZHhWCaTIP+zHvnQI9chmbS4GKRkGphvsxZqzH7R1wsQnLTIG2ttmm
4ZYS/O+/ivQmQi7aITXADPmnVvG3ZUqTvqfPq/vk92TUq3wvz3x4SPjtRz56
bA5AOBgjg5KVw4YGNjlp86Psfz8QFUoXA/l3Du/8dglDmIOqE+lXxlCpZQdJ
Gy0Js2v965Dl8fBI92P1l6CW+wRrZNCTaFeaCfMxfEhdhg/x5UJR/DzRmpLP
FiQCaC9l4VQ0wZOL/i/sHkHuAAYfv0QDO52tbuuw1ZztERAuPTPFfc+RlNMJ
YcUz4CvoBN5rpaLg/VFefFJ4QfgTkUlOTOQIh4BfZSs7o0z6Xa8Ym4kQSO3O
Yv5jYeIhcgZxV9n+o8WqJJ6/zoQhqe6PxUQL5Pzhy1DKuorcz+J4D1sEqmrH
u5k5G+I47WuTXRaXlWiFfEnvuAoDa0LB4LLF+lu66Pq6aaTmgPjdqaey92bT
DYEzlf7bkepgeD7l4QTLrYkhc7pT1y0MtNDpLiCEDUgzWVdvS/JEXpHyQEi/
RNGDSS0jHZ/VoyxTs7urFdMKUDxEoAecaUUsgfMtPIkUxeUnuBTfIW+ehu5+
tLPWEETiVNwXjaudXTFY6V76MgJgRl7C94CJbrU+4z0xvmQY15iQDKvwrH9J
+v1mtFt+RddGpJbHH2PFmFLnqpQtTC7V+Pa4dfGGnjFa4OUWLPv2jzToSUdA
ftMJTXSYwKES1V9qGogzK/rGY/k7C8RJI0lczTk2aHlXVKHq5NuYIVDEVarj
pJE6YjP6Mv9ESG7pbv58fOaF6rmYkj8pBb1ve6cwmdo8rV1I3ZftomV9ue1d
tvjQbLm7yj0puUxs2O1Bv/kdLVJJCastmcG4EiFVZfPUK+HQVOnCfu1461xz
anvm6REPnNjg2VSdo5HdsjQYD3lFmf1CUlEUmxQ/6jkuR6pxSTUr20wHmO9k
r7yFI3FnpcDDyHGf0fxJgGNgqRdC2megVgyZi6hPYLt++zYRZVA/4AAMa/gn
78OBnieK5p12qgBYL9TwZBD1FAEq+opAfvZqoQHD3ASWIL1bEeaB5dRoJ5y0
3xxAiYl9OwVpOMhMdfh0taSvDi1/3jpqnT/hVWBQW9BVDFGz5GL0yRuBtQCT
KzjeVhjXoIhHdvp1LBVnp+TJ7ujPQja9YwryP7NCqN+S9uY1DJIwHqjnL6M4
4LjpBlvj1wwLTvfF5eotXcKHHczliw/SF9bTn/ceYS+iDKcYFV5kz2ccdW1Y
dHZz/sJ5J7jNT709HlloUR0HdlWjOr4NVvI46r1EFQDdlASuiH0EvFZB2XUU
tbcJg/XNFLOJMub+6Sxn0H3FvMDfVoWL7qN8/4cyEEBlJtGqTEyi/zzb+Rq1
/Uk37jJtGN+cyzWz11VqvNuxp/TGuZj2EO2LycEvlMz9eF+EaUCVGzsdazxc
HJg4cEtQGyemtVlfiw1EhPTEOwbObpb1/883V6Licee9swQ0j6oePUPA9K/u
lSRnomGnzfftta7VbU1D9HQaIWOoMBpZRi2ouyHPephVCvQwD+lXvmIPJ8vP
6uQBgvuTYCq7Xer3Lyxq+q1LKxGIZEZCvR4y4usuJp6V2JsQ2272GNVtXB8d
3fbcdkDEtF8Rx5Kbybud7Vce3V4XleXKmA==

`pragma protect end_protected
