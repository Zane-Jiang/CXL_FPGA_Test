// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OYVcVXzNAPQMKlV93Waz7ymkuHuuoVvazq2YE3+lAx/Jq+9hIKZv46OdqyxZ
kEZk+Cfwtfnhx46J2kSV+NsQIFnK0Y3w7c4/TGTl6a8Uj7sZ76eRtyLiU9fw
YXiV89jIi5J+zQb+7UwQGixmq5o1dou72MJAsxzGucUaSrKGPXKbrqdc/Ep6
BqRGJ2BodmeAuHdDtUsGSQ+hb9lGv9KjSDo8kKYPQpqCoX3bo78x6ktvCimr
418wX5jNqiWdKp7y/NxapyE8hsalhPv1ozWfYE7dwG+zqoyFdwCvlwim4/CE
DfOyVHwHDIAd3YHajBWVWZFMo94Y7+ZV/Xj25tD5Lw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eg8QHaVJZS6qHWx7gl4XqMUlDJKQv7MWcAp97Pyk5eqLWxGp+qgxYri10Z62
ABv9gkz+B5DYpO4n0TArNBsW9M3ITXS50I7AJz220W2/hPPSwvZbAF8x/AMG
q0PPOyLxwZEF8J8KlYzO/QNxhXfeCrFnRMECwwkF99WAGcJsFNMthrBMVHlQ
XgqefS5F6NPU6rbWMrqN4r/7KHGUnY9YDTcGW2ORjtTWFxkpshg8eIdG6cwn
0XviXWBnvXZ6yRCbN4yG5/0TY+gj0505zKexuWOAs8p2X1TNQ4bGjMHcVB+R
iOXTHYFgiXd+2lfMUgy17KsJk21PPar6YytQhrAlJw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Iaix5cW3QXzXCIot362rTYUIuhbd/THTjTBBEAhobD7IYNCc7YX88LxMmdzT
2IeAGY2EEf0fytWI33ai4e8Wmibh0ks+Mm6ojUFWpIT1NTCI+qfCRk3RAE/d
FI7krwLxKucxdsGw+fAKVU3nNy9OP1k+ZF7/hR+lT58Y86vKIyycPHIziu4k
9zgqbVbH/R2SMNtvL9YBjl1obZBCNcZsnL9+EZYYFUjtzpXtOZoJX+oLpXpU
CZzlViawwiea/oqwheU58UnJIgmFVRAoKrmYoBJYM0Pyd6n0+CIaTh/3+4iK
6cvMhAIMtbkKaTnEwHCk8aEn4N4aB8S8DLcTMduq1Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Jnnky/OoKkXV5JrkDEu+hctbo43wpndcB9DmujhoVhmw4a0C8YF4QECA4JtS
fhO9iAhqhk+uiBzxFdLTSLrbFgqSH710mUAmzFUVSyEZPy8qSPM/KIPwgANK
EArJ7k+PeWdCbm/MPmk8s8yRtncqzjWvONpgZRCDbhfGTPhd8iA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ED0X059TTyR8TM4iOtYV8lQRTJivstTmz1z4c/qcO4Y+Pnj2szx4O1oGau13
uCnTRvzfgXpSdQtcq80qYAZNmB5ZEHg7NKo0ttATkO+2TZEeVwQwc2ikIIxO
eSUKaJ+TsgwE6IMZV0XbZpoE92r88sPAP1M4rjTdF5fV7K8dZMMrCZc/5A52
5aZ5RzHxVooisX4ubX0pdFJXeFuq+lk97+We8kAGbrF2n4gGe67xBDgL3oIh
qLAKdb9wefqjr+iXBbbl6SB7Vcfh+qLZ6OYiG26xHezexYdmtVx0n39ssJ1n
DGDOkrGvfhiEg8ogQGkPLVJsblaMI4EK8SquiCpEQ7FMJq4FgUhD4rPCQPi8
tq5rTXpe7Y8wzPkwDB3bslm3RMnKe5IlYwchb22ON6zis5twwTectzGWHE72
S/YXySAnhOwYaKoL1cF5racMXcXwAXeinEY+sRErDxkz27Z1NsnziC3zpsr5
N6i9R3Vlmy6FmFMnbnl+Je9lMLv0eKrd


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KEs/1hYB0OXa0YIfDuOKk15DInk2Cl3lsHDj/9sdykgXw3zPcwAMoEbq70gK
LP82QohYr9J7ga8RD+Cl7LgaRx1n3GWFx/Nkz4Slk8KXIEmiGCR00nVwV+LA
ywkwt5ResIqZSIJ7rLFhSb4CXvWI8Gz5wC6e3vfqUQ/2pF1D2O8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aM2iCJSOgFr3q4cR5OcuKKoNUQSsqzoaq/rXNUeBDd59+i+Cj426rXiBSRfD
otucwcrl8BodaKr8gJm0NXBSuVw34vOtC37z7cUyX8oINZQps26sJLK29Z+r
VKw9yHoqBO/FTbGrTJBM3g5s++UEzRvMEIL8MNn/oo0emEhwK38=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1296)
`pragma protect data_block
XRbhHEoFPWO4Tb6BGOYExfv1oU+ZF0qVH4YaLx9PosooE5bVttuFqFaOFh+H
wXe/33hD/eI8/ibzzO/JezzNKiCMHwJuVAczj9ja2kRd1WgBubbjlf/LSQrf
mFanoZCQNLR9bY+tDvwpPgcARf2a1dxS4cnIDayP0YraH9SotUidJLDpNHtZ
//30aYiVdKzpiv7LN5LSkLzR6gjxBgX4pPUymDL3viPCknwoh+XYsomb7DLH
DS4taiedI/GWK6G8yt7R69DOUZYLkQxcd5nCuTvzh2ApePoz7HpOuEh4yj6m
ubNeeHlLBf+YGZ6pxYr3kRLRHZZImSOVogWbaktPnYqco+nkLoJ12K03UL9H
OxbhNhogvTjz7Dz1+OiDTaf5fWsnhNgYUI4OcvMOp0IonagxLKAaOAx+lM4U
M9TKE5/W5+/18YDmXMEGToYlyVT3Qf/FyearkECKoD7/iIcHC4mtOSFzyRVX
hC/5OL4q5v+rh6xjLcLsXyCepbESYSyyOqSq0nGTLI2ZoMvIu7u1u4eijh5Q
7Ndsmo8MoBxXF13g2OM5KtoBgb2CH/wt0sJ0lKc/7rbL2Pv2WEK7/0Sn9U6G
3t8qEgQE8NBe5qR2iwd/+J6hyFeoh55XXE6AL7ViGGHWQXRdI33j24ADcl/K
690+v/WdzMCbj5+8IpDpw1Y1e0yJ2LmupE7HouRa2AVt10JFVmgdP7S4bmCL
BGzQ7o6hk2G/kLAbH5qI4dA/bfEKjOq0Zxu/PFL0IfakLZVzvPjfOpYqTYsM
UhpwYHTd7GBp1eNl0QAR2IeXPEM8YHYWp6gvEBzEDDw4WKczwhZl8bHxycDC
EacWkq8uzR4y4zupv4vqyvde4rsr1latILCq+ipHmB/jbT1Cm/IhxYjKa1D9
Gjin4AGENbHT2q2lG7wA1d1Rj0C9yRUQoWrcAoTrFxVfAIjDHt0Wwu2ncRul
1IZ/nktWpjQ7vO8TvQMvohO7IE+N7kaZKCdG3wKixhtuqOAhUU6Hxg/EYwpl
F61PTBPmQWiWHgsmSWZl+h7LFM3AL4OfqoQ9izNBKIIg3SIJ+V1Y/Y2Jlh68
8+LLdPSy/PNTZibqVJx4eYBK8yC+UyqWCXjI5wRsnhLP/21vPm1eTJ9zu8+C
mHcCEdZ/Frcx+yTXOkCtH/LQ+kprJBRXt+JIaTOfP+mN9CK4XpJ4gboJydHC
CX4mJJe7y/85uDdw+thPTQkD9f+IK2Boriwmq59Dl40F8Fz/U6R++uLLkNda
7C/4N6dx8YAwEROYciQK2mbrnkJ4+b8oF0Y1TqavfOJC1sG6TsY6vfWyq/qY
nY9WpLfWnzdcvBWbkC9GZPjzlpsWkDdArgnnPI3oMGsX7Azt9SGs15t4b6M+
WdnINLg3Ltzvo4UqHfom2EWLoNfkOrNx02WnF/soj24fpV1J4SWBu/yTYtRT
gn1rl82r5ygGEuxwOOaAHISzgejAW2KQWj3EDoutpgPYZJtiMYVMnfWvz/A+
rNckNDa0THPf8A62/giY6XaiQhKjxr6ohO4+bfcsQuDPs4Wwncs3ekiMXx8q
TecDjC9wJBf2lgWSgcl8lJJkP361Mi2rYHZHtySDtqe+lV6bX3sbKDS2CCtH
/8JmubUf1TK+cXk6FTlQUEE4Im86gLHFnAkVxxLX1YXOXNsLX+2znevt/+Gc
UMQdI6rznFmCaO8XCaa6uH+4CflKFzdEpqRPp/k2XKxV8UMQ

`pragma protect end_protected
