`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
q9Y/yqrJJVx0YxqBtzQ+ByFImaOYlWkPmH04Re6uJ+YxqkOF/j53kNGgpN503YYU
UAHUO90tXstKOBLx9fw1OgN8yyeXezXo17EndGfH4NTJt9cKnrr9m4SpkOL/Bnpt
QCUMh/FYglG4yW5vZ5Ms52h3oSMxLJV1NggHWJv8CPw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 22256), data_block
yXebmLLNngmngLchO2BC3hOGIbtHdiB0NUD/x7I3W/buZE7a8ndTiXjq9LgyCzbO
+LhXZSiLRnL3rL0EL7jwdGC8NEuar2rHx4208y5ed1rK8weZCg++1hiI94vKwulz
qVadDrF5CrD8hkfDs2yj/X/DI2rBzryhIxw/Yjg9dl5l4mrFfjPdV2ZCQoPNBBr1
IX4x6+jdknOlKhZdnPSah6fShl9Mp9rBOkEh2diHy0TDzsUQ0mbjOOUS2+udD4rs
E7xv+0WekmSaNWMKomkLqin7qRozXodLe/YWlAW60R65GgdZyKWoVhFselkDpj5l
PWPkYf9p7J7wuOEOdkppgzg0SCQs/5vpzNk8JAW//8m8PV8qdV6Dwf76yzdIAwGg
srDplxOlANCnmrQ4+8OHvOPoUcWtj0XVJ+PHG+U5YJIQ7QGQcApWwAWcZMOwzHgs
fmxaM9rx2k8qQsGxBU4dP19anGnQ0WcUFSmBcy+WKXujAK8YwnFoND2rB+OirdEW
lXq6IJksg5BdUhRRrbcdisau7ViBqOL6HVZO2jPtQ5vd5BNz1b2l7+ccrapzi9OC
LxH75dGrqKgwCRC9EiYkymJWMseZX3FKNA8tKOkJWbhMNMgiEDqgmEAQCB8IM5OA
xaHUSpLtp6+sXP2Kweeq7bdgrr0pv9NOXWWv/j4bfPdREmYyFEP9iaOI9WQZo1Q7
kIwUqbunahIPoJ5C4rrR9wcnQAzhFbmfjssfyj4Idd0+AFBthDMYvr1HNugDlRKC
PD33MjJuB4ls31VG16i6RPH089WZyOXootuEnQTaELZG5GrPacn5ZH7T6oWP4/u/
VfDniWiwq2Xh1hr7kyXaRr1aBEGyuOni81p6EEykZBrb2DZXZ7e003cPerv9teAJ
ehgyuz58wDVZBXUmjMchZTX0SHWJp/RYZgOSx0Yas9+VTo8H2LgeWjua1e59KJzu
PW6VjSDPiPmHbeC0cT0meUS0VzoVd7FWF6curlWqtPOLLELvmW46GBL/dUCZpBZx
Yf5O7IR7nRMXllsiF/HnkMlQNJr6cnw0PX3/zO0idIDBkwCSQxRj2uyoEVUSXbkE
/qq5tTiQYmCWRrQO7j0MHqPZC7imwNF61AmbRfQ0ajJgIIldiO7B9sstp5TV1gWl
bDEN+wEpeFbbqIgcwDspELzfOhrUjVIPGLVASEtXXSmN3/NIEJeGy6Q70y7Kdbhn
dbAYBMmLnO90IVuMHuMkxcYp65QLixgapztLbULhShyZySxbjJ9LKVkwP49J9dfD
u9uw74zVL10elxZhZY9jad7/x+LRxxxQCn4vqyVa+xExMmikOlJOUhPvGTJwFuC1
XBOcOkSWULHCGFMvuIHoATn/rXtJQdhZCpGdsieacXRNPA2uOYwUq1fqf5Gn95YO
9PB21licBdd36l8NdjJlM93+pFAyo3A6zoQYebnBaZXdyPtHSPyPxc7ogknhtUgx
mMAhlQC1VfiZSjO+Iz8rhTF5BbHTI4GkjiwP8+1/7KyifulygIumIkqvgw4I6ncj
MRM1cTHhhbahXsVaBAgW58tiUMHrawHXjTp1P97+6h3Bekwu3LhFUtJkxFX8wkpT
7uPX+Y7ozx/lAwADxfaTrmiHIdFVid4z+8lCaEhf0zG8k0stPuP3OSMoL/ot/4a2
rqQ7i0jriYx2F+w0IeiGYJqbhcGoHlIbkf3o3hQWWB03hr+MLzDJ3lc+2uqQijaX
EWu+3FeKHC3WS50tlbrocjaQAG7FCzc/3c+Dlu55z2xTLP0KkhrEvzCIzZGaD47e
T46wzBGxEpW4e8UebJ0gZWMmTsG+yEohT9L9ydz7Kox41hjujuCovDqPUKYGDevS
rsWl39liQFC4K8Fnx/9MmNRIzcB3MAdQZ3Yln1faFN+zeIJ3MQIEehfVInX2+CuY
jxwZvaMImdOfu1ChDF4ZtawzoO0IwwcFIDxBs0qxmLHuQGAHbMRKCDldIOHzpmXB
36hQn3zXfJ8SRLD9h9Sh0wSkrp3ENPbg0XawqkycL+YSq/sNGHN6zEUTTFLVgAfn
bkgUE15ylMv6WWdu7TJSTGvrefNhFhdppgGI88+Ppscckk9jqsEH4JRbgcvGw3At
nAIhZnL3Q9XBzc5kvX5F4xA8iDL/C5zIemp7/3FcaiGCSWzPGloda/YorVkBkMj0
6Pz0d0O8ad3sAqnzDpKm1X1507+PybyObtKYLQAi9akdnu/E6JOigIW7odsS+seZ
Fak6r5NJ8NIzFDLr27htnYGvmjPeGRo4tzHZxvg+CjYIrca1M7744ZV4uwc+9/LG
QVuTvEug0V/E93Olrl5lwU051w4IgIbux8V3Ac6zBtTltJD22d9EEGfapb5QZ5ui
bw7A5isn5xxY4y1nnWxZ/YVJLYayAwQHxogtCeuHmVBmRBTc0fJJSzmyUQiAXydy
WlmpqR/cywEXSb25TZ5bnzSfdu3e7VSxWZ94rD9i1SXQrvP5yP8BDVVCSLgLpmHg
THN3nXjjT/Re0npFXbzJq3YpbDeFkQe2eZa1+1IThg738E6qeBby2pYI/c+b2U0B
NDzcivN6RpcwoEeKM0PtPWo57bgN6yNCok72RRchGTkG/7xfVQrYwpS1BKcFeo/a
e9YiWtJQSrpQPPkWhpCDH1HenvthYJALqD5pQL9K9fxsh3zNnQkw7ox/kBXZbLYf
Ov/ZbabxLLIAiUaDpx78Tcj6wEVEGFqPDl0OiNrsvvcI000ht7MtuYSORGF4DVjt
VukcfZOgvpVTac8nR1jP/fgyxoG5GeKAfJqwuRkOvPeVqKnr9FmvEcaM3LoBOuye
Enxf8Y4FEfhWhxbXIbjJMosZYF3KWOHdqqar3yAV7aeu9ilzOsvf1ugRZ2Xl+R/4
E6g8yNrjJiNP59yKPOG8berjM+T3bwifO4njBx6+4HRXrYdCXo9qrd9DJIZSPYGX
M/RfXXDGWqjEPWx8B6RYGFCaG4+gJao2w8uuF8YMlnGTOxW4cPB4jdABNCcE/iFw
lxoi7/RDdilxLAk08lWTR/g5TWiSIFC4KpxCX/h91dY5f9Nrc//l7D+FK9ONpGis
9Hp+w96CvGFwlGodqUkDXYAvikxFNpXvFMbi7f/mNf+mXVOCdOtI5giXuJgpc0Wf
q5s7uoKAdQaGZ9uaxxKFgIUYchtT9zZu58ObmgtD8KrAISXsDRBPEgMpuftcrUYq
QY3nzWU/HdaS0A6Ru43eyovq3EJxUZPbWVTmj7PLMOQUo0JdaiK90GYpzT1eh01Q
IAqd/T/k0+nCfxVscJhM9JCrSkWwq3bpVGTMoB1qjBwf7+Na4njTX45qcFRI29jz
wHN6kOGPdtV1r9joHc6z/vbO+Bb3OLFiYznkcRoUfdtLHOnahVLZpSa6VCrVf1pw
N1/5ck/xobVBz7VRia5mvcYyTZL6qa2dOwZyE8uqnXZceEEkgFJfc7DXtcKhEVcB
zeVw3UmJXGJg0NlocX8uE5aO4vszeMtyOy2vJ8/BW7tufQ1JOzXcQrDPTam/8mb6
Vo+Ud6Bk1/5VYqzi+3cVqYaFt6nzXRenss9pa5ELNrIqXBO9q2D/Jc4pirsnaXfz
THy7etf6Jkj+ZJ/auvEzo+jVVTJbltL+iOrC4LcZfnzPv/i5NAnSX6gJfBj0P8bw
3zqcNgMCNlvIhxv/WPmKXSH5aXEBphUqOx4yff4yA/EUle9qReNxXFdTBIsV+BKo
5L/hfrMU+wWEEHkG2VPQswhi8S1DeiBB9sNI8+/pUFXH4rVGBcAm7ZWZEp5+SpuP
r+1fWNNqUlSacSlN0h8wMWQo7+cgTixMWnRpSYSb6sbJcPSmFoNIQt083a0m1wnA
vDVZGsXtik8+Qdp2ysn8Io5zra4FL4sMvNBs/IxtWL+4HXqVM2EBS9CJeCxciTKy
Tr9xlViQnhk+HuO0jsN25UPqLWYSdp8qKv+fOmTYcH1sW3X8BiNTXq8JhOG2JxzV
E2dcF3TD6/tFr4he0YV0uiLOIDR1VzsssT3PxY0HLYKKAkDHd7r01v/DBedBTCpf
okhdo4P1ke/te0YEp56PuvQKAgaiIWtPrsbQPQM1LCLdTohRddJDv+boyOyTc46j
1DspEFmDHZj3MJHxQVJFc5PFC5JDWzfio+XZBmc7LNEuLarNMo1oMCVEDkNQDH8A
7D+cOJdQCG3muTbUKchKLKUD9Hlg0E/18coplhSKCP1Td61n0I00QPDiIBxA6vD4
mp9x8ioiw9gHFq3hDtf9OkvpxKhZKJvKHnFXKbNMvkj5MCxs/qH+GNTGXvOlR0+G
R+3KxVdnk2Vso8yMBO/TLnReowW24dyJ7wG7NFoJgLBgqoLKMEXiyFM+uGUMOVo+
UxMlrjG9rEYjyUgw5PyMDBB8uFyYiOo+dLY5jWB/lt+eG6/2ls7C6dCHKaiowhqs
58or5TeGptDDl1zYlkqeBjZyGZMLPgvwsP749EugA369D6/0cQXUDFJtl4gjciC7
Hy6PQUb+IAi9M2gGGict7YCHzLDeCobJoCAzJBINJvBdW+0ajcRR4g6dgWpdIVeD
uSu25J6V6EyoWVQ4dCBfp18G5FW/q/6Qg05xLNceoUI5k+wyxPQkM7LjGw+56FDi
/UBEAts+pZgZe5Q1Q4dtowAo1CYx5eeANeprMz3JZUFfCJkRxTMmgbeHPZDGv5Vc
0nUMjNDKRuvgOgWeTahgVSU4Z3QkHRNjKzTXUpDpLp7sOVJKAWbqTdY862s6Ag88
ogkZhQJ6EzDfJJbnEwu4qEOak0DNCBW7nOOjAwWpRMoOllp+9LTfz4Edt70TDOxg
stc94KcRGndrON4RoFXkzXNy77Unpi1BTWosJSzmS0BAnT/oOLF/0oWvz/yYJe05
zQj9BaStGvWPr5En3MB2gNnXPqmM9k+wmzQU4TxUp1qeIgoxyJmPQTup2U2lyICO
mPSVUS/48/s8hwbhx+r2/AAT9DF+iOMq9FoRg2K5wWbMUL9cYFgKNUNQBRXGRElF
/Faa4XVN/yOWJmKCaBVHL5E0XGa/8k2PXDXh4DQ6/O6ekLI1uyK6qIMyG+MvxYkh
+iuvCaA7lgmeuUFwXEvdoEHoQAzpyGobi4spNqvAVupc1fXlkjArwUUaYH/ne3wj
3Lf68kCOmsA6Ivk/droTlfQJrkeutsgaiSHKf5QEFBn7mOLq5eoFkWkidumyCUZh
PlEDLrNB27wCOJyOL8LaoVbfl+xcVqz3vxDdgStSby/qtGjrPKpiQT9BzepcyVM9
n/qwjptOYGA2SpHm/lRj/fHk5O+Xp5Iy4IMSxXhhrFmUw4c3R/HE3RgMTsmRum34
aS8aGFojzHax12DmpUf6034IQvPCi17v5Nx4rWwV/JpyIKotRZu3chw0w2fLLK8r
mwJaMlC1xPDU7v6oLZyPTj4G/UM0utz9pfq02iSrbSBAqHr+RjgXNgn/U+F9mgPl
dwTMHHrwiGGp7a+voYoo+fTSFq2FBAx396QR4Ugy2xO2Y+YXMXlKB0woBZ0WoXli
4W0sIQyjxET5Hel7j9atv0l69XNSvJ1Fj3w56GlCNEOIohUGhRQzb2AuzlS+nUUO
fQcqXGsDupsqMmglPuQeZQ8Su0AtmuzFTk1XKozGvVhuOAAUozL9ZASt9hZItqox
yiXHfxsjAuAVnfGx7DBQqCQsDJqDQNa3tjt2E4GJpHvOnuxgr8IEZOk2C1D3p64I
FzMUql9bBNSy2NVCcu7cwonb/asOI/e7A6DI4AkFVhNHLgYma0pdazA8cnIopTQJ
Ov+UJHesb6MaaDajrhLsvhTcMouAD9yNVAsxPkktnHEGxccNzQDg1f5A8f2XbUlC
gtgLTbIVROt3wYXymAG/FC1m2mubQVRjh41TIwPMnQDFpTe6xNUuIWrzPdpQ42eg
lYdfs3+XcQIC2c1eICJTda0YgzX/yj0QzanudUr312WLPB+yU9Y7jfVOBH8BpL+O
8VnTt2npNBabk+ew73N9O53Ek2CsOQ78i6NOA9owVK/9q8AU+nnh323OIisSy7Dc
Jv2FkDdo3C5mGm1hPvOJ6kzYt8BWWaW0qx73I6ULs5pmdUv/4Z5IUR8LHjbdfx1u
d3jFb8diJzdkvxhfULsVnENlhB0F5JesZ1MdG5gMNSZXZU0kpxbY5nhGltSK3aDM
kmKcOKL8tQmRUrQAoASZlmVCwZXTzhiZmpjSnKFfuk8C/ac2cRHseTJL/xvUldog
ZxZfgXL3F9vRpGuWdRWP1oLNr6LqbyxOfjAehzca/coJOmRJJwjDyVlQT10IB7Vo
/kO6QXFQ/PBahL/hdwnPdTS2ZHoIL0ED/ODRT2Sgqrtrmk8SRvgFr+kCue0XeSta
zlCSmDxkfRZkaAf1IbY7bC3CJ8QQSCXtEjhBjPJoRUqkOFHvCSAFFwCnT1Uh8VyX
yTL4d2C+X/mq8WyLUNaceN9ALV5htftAzUEOIadZfS6JzlRePu+9OyPvZw0l8+o9
tFZdwG3qJFCUXBwPw6QO/uo2sOjTOULH6JytEG41+AMXX9/cfMR0BReOQ+hdJ36y
McvXSa+noTIK3prm2qudot7Deza1mH4u2CTqf07dPlk8vPY/0iInQXQnDH7y6hwx
TeBzl7YRqkojJq0/Ev9sPGnFpXWmmSg06w4v5jYmuvATLvY5q5Cs2gM4eN2d9eTX
fZ8PCJVtI/3QnYeV+JHDwWz6oxHJRCEGItfGRb/UUWHqP+ssT72TA2zyzvvOYt3s
J1sy32Hp4rD3Pq18o97A1dP3vR0/9Tld7s02LsaNLij/sx22kb3K843gqmu6W+oF
11f3sSa8OYvsh8NmLiwasbYNxUbvN8dgL8pvPSa95k95RBm37z6j9T93ewU/9cwd
38M2yVqP7nEPn/EkIqTWwLfZWHyVwUs+P4/fas9idTqAXtl/cSqIFYCSZcojlh0T
dpGJGJ3Wvruic3TxkJE0qfCQQdJTEfUZHJMO77PrC5bGLYYWR/FC5YAW5U5XMG3/
QsblzJG3HE19bkOvZ+7YvRChBJ2E4gqleHT3RA8NXZ75oZX70UlitZ9HJkr7Iisp
BZsAlSzuQrysERRf8zJBCwjcP4xFTCPJi7ihKxOxz/RnD/kFTBzfG1BGD2KfDdyT
xgjbGlLFFkK6AeI/+8bg9OPCXII5ZWZYIYScbs0ezwZXZDnAiDIBOuOORUuw1Ble
6Qeaycik06vCZXXV9EuxzQMS8p/G1cTMsa5tD5C0T0ZubTVPsAmR0uIDFgBBWvsd
L5OemcPZJ8FSkQunICjlTVAbsq/WBhSfcUM4l4H/fMvK9c2MVz2lu76sNrX1CzFH
3wHt3j6Bt2T/TrFY2Dmk2Nmt71eR2Z595plqm9mWXQlyPM12MSXFHUABWmSzyG18
VUQT+3TbiXMq0Gk0ibQlPuN5NVPv5qr4vR1gxoqQGefNpbdxQfcyV6MB+Lu7XSia
jBZSTz/UxkwKYnt6PPQbFTieY6NnWV8micEX7pSoHczm3RzfxGW9OLUYVf0TmdUr
xz35QTuZaUJtOT8og28S7RhqFsGtVsalGJI2faoam2MBFSw/WThd2r9mGvDElVF5
Gf9nUtLO0sbcKm0nbp+jlTMPHHhA07+LT0FKsrlAT/PHPQGJ1rhkeYcfPORJiGyD
ZA0wIsqmdOBTMBhQ+KjhmZ5UVdUFsueT8VH/DDwtW/nRNTxKOjDAXCCAUGPxBvRI
z2iz1xRGbM23P/fi3PH9P+wVUsxirX8Zs9HALE2bCUTnHYFfPZqAZSeGzddIyR+b
l/MmGtQPEObVfBURDfncDFN0KeHT7X4lUIOmSW6eNj2zudSfBTeV3pQnWRvbzZ1w
LXJ9PyuWbRV8kXKxGV068W+vXJ9gn+XQhJwkNgaJRAspS3Ei7GQvu6QIR9FMFLSI
2Bh37Mqn0v8uITlWUA9YJ6EqMZ9QxlyrbeMXi52WJ20a7ZYXwKoWMoIz0fn+CXQw
VxDSFQys6ABduolS5Pvd00w1UzyW4bikTVPyK7M9scroIajObgcuRvayg9hloone
IPzCRhE1XnIGGqJhxtJwAO5P7tt3sc1oC7zsMF4SI97XcHbTWbhBC6sDBO0+KEpy
Q0rpJArTpjoSdbksWWIGM/paWzsTU+BQbzm9Y6/u16DuKJjlJwA6NswzN1OnN6Lu
elMs4SUUXgq2S3R2IyuB0NBdh9ex97PGag8sDO145wG5w+uKrXo1WYmul4KUiOi1
yVFt4vU8/j4EcWH23DLQZybShhrp5ogj4ppVS6CD/25v96Aa+VHOBjSfAIGASz7N
VrINF531yr4+qfy8BG5IfSWYDabR9pOQXFlQ55OYMa7u46HbSZQCkCwqUtN6wSn4
tmRLh0leRbQHgwSk2hP6T1OGAq/NAlsxujyqT9QSj7T7imKSsyZ9MNZTAi8Xt/If
OICE9ybph4YGl2c2MB2XRO0zMTUplsaWhiursf3JqF7tOO+NOc/B181NSZHC0lJq
yCUNw01FjmkTG30TjdbTb90/yF0KJYE+GPkx96Ksz5J09qBcREoV1JvSCuCKFgfr
F6TOMdwvB6SnU9JAwimxB7EDqozjV9iDxY2ygU1pg2mm/rhIUbAPfKMmtreg2P2n
oIClXnUI5vQiKBrbfvdnybeLmqLYW4gMDYzsTO6dPdfdh/U9IQmq1io1odu+5rUK
uoa4disWcAe0/tUdG10iqGsR7hY39X+SoXFj9DLvug6fHNJNTrPyHO5JFDXsLHqJ
jhvvRd3id4j1VbbhBa85/juQmmYS7kU/ozcrclTa0cjbtuWnaRJqO8NxbYv/pu6w
BpZtj9B58dxXYDkyNzUdVMVnpes852A23ceJ8mOmgDFir+e3JK8udS1s5zjaHVGP
7X8DaQEiu36ypQAfL8FYL9EB7iGRAQYbX6B8YfA00iQ82JFIocUAibJCVVf/6mcF
5PoBD6cpBachm9igLS7Qo00/y1fj7zowgsq0cXFDxO7j2CR3WtCXCu8823sn9eMV
cERTopIm+P50ZwgmvwpG5h6aGJR80Sl9rZXP9bh9COlJqo3K2o08/2Fb7/Z4+Zb5
UNQoq6/VGglMtzB16A0T+8Raw18BZxhZQw9zdGsuv1nzy8eBUzLx0MegyDbFDGaK
oV0QUXVhmmm5mhDAWba5OKjKYOGgXAYJ70LbwESSeQxDrxdJig45bxeTruqWdUnf
LkEBLDbhRZQlMYhW0gj9PhzrsmvvDn/wB+LP/FOBBk8/5OkmIRZ5r1MXTsXvybCk
GpWTQ5kwaQ05l354ApvY8tcM+aD6my7hnUWZ90wNkdvSLgzoE+SepQmQKVtXic9X
o+QQrmRrSy8/V/NZ13F+3QTpHpIiaUD3Nj9xqRZux1nmP5jUtcd+voU0/U7Sty+Y
JGMSW9t7mt4y3HhKm2BHvewGH5qHEoSmDLSctsLzSRDRpba2WpJYxlD9veAPOhF1
hV84lRRrG3WNt/7UEzvuIUNX5uF7PRirmFZdiuq7qZaf1wxFE+dfYJCKsOSWeHIs
UfwzmaJ5XFq0wwNKyGg5DcBtnkSUatvCOxGOJQ5D4NqSw60hPYSgSx3sUpNVrPmZ
CBIapbFMT2tafTjUcI2byQKOxaj+JZuEOqTkEf8u22KMBXFCxvWLvYLTEd1JxBJa
/+i3XV2Uzsnx0N9kW+4n5OozMZI1g8gglP3fEgSRvHLDIVklJ0ALItQto5KYuHIA
OutMCDWJbNkq1Z2Bp5/GjxhZgELJtY81qXCMbMyFMCVIm3aXoZvocAgsVQVQTKLP
EPcbhJkkQRc0XyIymEcdBDOKedQT2fPreHg9N1PapNSBd20yM8y0ycD344EhtXCR
AkEu8a806VH0INzn4F3as8JE1pl4y+4QUfixccXvVkwo2dDqJS7zeG7Xvvjs4prL
Y0/qJAz8Dn1EjPBDd4QhFdlU9GKtcPyWq26ShSEdZNY9Vc+dhnhQ2Rhvwe8Com3B
rz0jmxT/iizpMNzSocmgyVkDAn2oSOdSsomgPl7xF4jfzxVhzoB+zgT4Re0KlIoe
m+6JmhYN1vsw0GZeNluJjL1XVTwKcoMsG72gxJs29RAKk+mSeDGyMZfep8yiS775
a/tsgpWoA2XwbMziCEHJ01cGIvkxrbe/CvJFBZLhkDEj5f70DH3gS+PKafg8fIfT
SyVEjOM6CCH1SfhTdgrJOPDcIIfoGXQYqdIyVLo+DOIm+6IKqqsZYG7aFTcqgNBI
7edt9QiE3nODY0j0bm0OzvkcvhwMoVcCbF9RXHqb2XXB6cGSilg9O00WQcrD+emY
O46YikvMsKvlUpRm0ufPyC+YKLgHv0Evf/plzab0wPQaqRRa2fB1M4wi4+DiJmBI
DnL1nBRDNqZd+0Qt9bhDl8jQgIZOI3OrzqKbTQHfxeTpz6Rola7vXb3o+6QSAn1m
iXWDE4NPH1QiIp0E99rr0MW8tln1fnPagSAYVntQp9s51YUyExLI9ZFo93Kt0vR9
PnDxpnPr42aQWZolV5S54dO+QXqEcU9c7edOt8kG/xd2exWq81dIvLMMf3/DlDUT
h1Zk53iLwOJtOSD4ZPtE1lek+JcWoWlQeatq8fXEdu1QXyBoAmMY50otlEkDABKX
g7niXRjQYEJQ7heZD0jGY+z3o2aofgj+1GTU6YAbpnvIoc7PClPhEPBYLqFKkz1T
fSq0U4uJWi4iVvJhN5vQZCw6/HAW3P6DQ8nWukn0ymjYqjebAaTFAe38cPeqpVYZ
26DCC0ER2dviAQoluw4LZnH7/FTJAhr20LQEHSGsFPG9BdJOd9jX1+dkwWcCuSmW
HV9QCFK+FcKO+XwNLA0S4GqfnWSJClIm+qV78x1cnozzCp6cEGo6kFCUpTjm40tK
VtQlYFmDq59VtAIWyDPzITZv7XoswLoB7HQ7a6iBh4fTQDq/G31npVjnzSk1SOZ0
C5+9gJYIE9zxWQ9GSqTGgY0eBl15GXK8WcRU7xx3XWVMNAFolo+xeJ5MnILlnajn
U66MnE3Pl25fUQu+jquJV6ZVfOdJWd/ls1+cHksWOG6KkDxiKI3GU8d9S+y7kvif
zCc40MFoQdZY36pL3G9i4RPnd+dzwYfFCaWXYbBGjga0EApORJ21xKSDGKfBD/tX
JXPMBDp7FofHmqJDWCF1jaEIqeD2JXm0QV+qYb7wOwPdbGvngPHJuruJZ3DA650F
DhafxPoHTvXFb1c8UenyH3z2wIqKCasixEs9/CgfYSILsniYXCtUZe7ldoi7PmI5
7a04k6n0xcOwzU3Ffe71UHyARfcmVRfQD1DHIs8n+EMQ3ED5iADOXi0R9RVZoo8x
A+M8e6M5mkomB0JN3K464OJ0kdndT+W1dkhauCcKko0EdzrybNS9N1qUeMKndOLc
qzomXs3BMjT6mOjlthGl4sP7qq1WPgLWOjTO+FSm+Hmv29T960iQdLejEFw0HOsx
8qfi3UbuwBN9TIH+qcjSWaGieTGjo3W8a5pGi+WvDJ5hrL1XzovrpqDbRo6Ytc8z
2TY4JqqQRxMu1oG7D/Ok4Ue7qhm8PlhXt/ZfteV8zD4zq6HAGre2NUp3vkN9LJYj
FtkPD0CwsBicVoN96VRy0OyxdqHVhUxPlYPnRAEb/K8J3CJjuPJgRqwWmI20soGw
t6gO4unpiBX5w7kq80J3ZFVNTBUq0VBDZStvyRSu9DgUbGD0VGsSoU8vwtd9JLpR
sm1PbqlGKLhdAyRHUp0ZKpYMEY4ohyKPxjU32G22RFFqVKseX+NOlK+TUgE/r071
4YHej501fq5AI4Z9whnkwNbU3OF6TNHgoBoMkkQR6AdL+1uhTOIrNYNcSs2UY1Z3
7HxJW6AEr49KLzxx6/CSiziBM7s8o+J7b4jxMmPlyy4HW5UbqqxfVajW1trlrDyE
oWpRYqawhrV0OqJXxoSSG9wWSfZ83yJaBFanCsS+UbCh3b8XrLb+VxY/mjI1iOsl
x7Jf6kFSiW8b6Z7cbAgr6JjhW7rKnNK1mduKlH+6+DuYbZjfR323Rlhw/iMjDqg4
2PWICgFXD9CWrpmxRUXtzmVl2MaOEXH7MeHF8xxbODuEqhYXoEDbf3n7TLRILaSV
0T6+UQMGoUAC9R97CItj3asuDX1diynSgc8NevRgUBqekcL5OsgdgJ361TIDnJFK
UPsl33JQo3Kvr6z6k3XdV8tIPODEbHTrwez42bbrtDombIWAAt7nRmQzT1TwRSZW
hspLFCzH+SvVGaptiVIsvZZTeywrQjXxuXebp6NA/sbpbFdm5EGeS5B2uLYB27/G
QMPouthMSwLkSVH7UU98oE1mSSnu1XngD01/TfRTOAIdXoIMU248tSFkEUPvODEj
lHFv64BuPp3yPwBIHniD9RaJfKBPrUj9mk+GGy0DteMEU8PNIbyV8vHZzTEzryFU
l5xx+uwEVgBhFsPfbn9XUvIfnWTwRXa88hY7qQ5O7FD3mgHihuTm7Q+uv1zDSE7U
l55K0GNs1DxivnpEZP1TwghdiCEUz5dgRgd+IHBLJZpAPEeeFqeJF887q/wURlUY
KikihW9A3rWKxLXsfWpNg6c5WSJ2XCtOI7LlbodWWzbNOWISJVbRlTc5YhXupv7b
93wNXrJqZDnohhpGmRigf0zhXUi3W3fZpv8E4T0zsX2twtc9AQP2+slE5MHTj8GB
AjVOG0Sb6X9OEZzm2l3i+CEqr2hicxpb3i/LZ2iezyiu78CJJMfVKv3rBRtAaVMe
bGfp1Nj1Xf3fVXvLnYRWoP8UrUjhmsJrHFf/OWtaE5l9yxu4Uf6FT20beT9ZxWHR
pcfvvpt8DCFiiL0SU23VR1wJx4xzSeBhf2kh7HR7ejxO+7qhY39wOByvAbK9gxcO
IIEdDeMs3N45nzkZ9R05Y24w11iPJbU//DexZn15S+xL7lSdiCLaWmrqX9hdERoB
hGe0GrTnE/e9Mbxxk1WY2oZ5E9vU26Wzwyuc6U5Es5S29nwSji9svaju/dQFPn5z
w51EarEC3yBSAoQpDbURL/qchmWDpqHwl3mgewtXBnRAo7MAakAffzwJK2YnSZkO
flL9LpQNwy/t+vobCKg/ib2yPcERKUk8EDXAlDPOE+5PTOqyey/mGVkDBTvZfuWu
J85BGPAyYSCLPQvUMIVuzatVp8yboQTjf3RqA4QlMgTABlzmFv9YXXUmjcaKt2yJ
UN1ULed0Mz3d3tGwsXFns4YZVR1nc7zjN8tn7aTfcuVAClw9ebt9nHYm3zg4vnEL
cs0sA+m2456T2dVrv04N5gpHYbvLGgfoHcd0DqoIAw8Ieu4lOBWhkmNDNCMcatrk
88a2Hgi4195lzLw4RyPTQ0d4uzWz0LSeFnsQsWrlXudLjuKM4AdB4UWBiNiehVI0
L4om0B7C1N2fPlH3yA9Uan4AvBqjTemrL3MVZxeOjAD4/GX2P7RAYlj/eERzAdD5
hYpQ/ovF9GtYVwwmfbYBES/tft5mFoFyiWA0DiIIVbdjQklAkWjUURam6UAH6V95
+XlsH+m89DNdMLlyS56n90PxOLNJwGmcUU4098mX79ky6OrMHTTq/ZTppF3IEjob
rSi4pxDDwqbw+0+/joB3h04Dk3Ti7sLIbVKHgYbPAf//ROjDFFvochijJ5nyhVqP
pIx6cob/ofZ7xxPkZDQyaMEhFfeIPOo8TO4w9cUAwY3SJNFMBhmxF+MgYdfb28fi
ZVBZ6apobV04mlnFobsdBouwpPn18XXeeCHvVYW8l6tH/sjjUPlyv5td+hu26jDj
9ChlNuv+qOgoONq/YQ/LGUmgm93LDqAjEmAsCuoPueGX6cDgFPvm5+ht+zqvUSyh
FidLpo0zOT9vdKcporlxYpNfLPi6SMx2UEn5k/MbYywNQb2xF0tx0aFogdUxjCxa
KrlceXkVhs+3/okntq9vM9l5F2Xg51SDF2FFRXzhRJnvqOkRHllIz5KTouM7Mzot
diFTsYtZmwiFv+k1uyFQtpkx3adfUrSB2zN90PIK8tws09y9UPSmpCqXrot9kUK7
UD9JmoUBWuoaLjE6Ikb34PaTPWx1BF918q9TZi+e3DfYkNGZTon17TVHA+gmtcyo
1qTOAYVIzdzOGwIhKWAeDIRad/8GKlokr7AxHZYTWuT3hW7FmxxjWgaLy8dnuxGe
xirUuLN1h5CPWmzVJDw6et6rn2iSLb8nItx4ELsqwuVJC8nk1sLBLMt6WvdBmaLV
TcJbsmZ3+0sAucWB+adfwHnsNVFCIqpXvU4iP1nUx6b0sXViRxNgrirL9M30ZcJk
AVW7McubN2ZQBeSwb43Nm3n5CR6Sw5q1k/zg/AOcO/voxVq6mghPDcf/y5DmS5hb
/4n0zbGDSgl1xDvNDNdBK5UWx7eORoXPVF1B3rUB8O6rEj6LZCNK/0LXO1yUH3MV
L18aygjHGJpdpBFEjucIHYsZaeGzhG/TvpNwjJ/nMTFP4CBqPd/EHMMVP2OuVsZO
Kf+iFo78d7wU3AInlOGTN5PTWaQ1MWoW1+k+qC2BG4zyq0N+TsFGeKjW+GzK30hk
v8nwZhP0P50FN+L8/+kChC2i4WZxrMh79LrpCdYERYbs2qkJl88K1kzBDJ0E9mfF
absyLih/GUiGSXw3DjVNArEAtCJ0BSXeyZV0QsOTJToswdQU7rG/zcS6Gdfk1/hL
i9WS87h0UuH+p4ggfN8OWpUQj59ctkZKUH7zyECqeQp57Y07fF3LXiR2cXuCN6Kz
QRf3T+u81r8wIcub+rIFXJhB4FUyYFZJA3G4NMFOO5b2aT1vwDWA3AOtkATCulvJ
5U8VkvEEVCmm15xVl7SvrDyWkyn7J39InVUIXuyu7xlGIfomOcdvvd81P9X24fC9
bOCN2raTG4eVLioSIY11Rjn2k4vXGQjKBhblX1iylm8BviWersCW11JwM2RUnZE5
SG7Si+qryOhJhNTbT+ZpRFizR0lbbB0KdoL79IEhD7MdSxCf7b7sOPGaZSFrixfs
LcPKZRsqed867gmTH757CUxlb9PjDGoaBFi3iFTH6mUMyqOYxqKNCoWGpB5W8WI6
yV9hR0msXeYiK06ExDMokTs8YZu21ksTmr6kbRWXuKv6I80YbBaCAbd7Pocnhc8V
3IzVDOWdY/Evsk+k2ww1rD7YYnjbGqPvGo2TeeuewSfkFH5Zd6k4SKSpC7sl2oqD
edgkPbJ7GOkyHzT4mvfW23IMWA6pfKB89H0O2h39tMQFTeugQy3QA3WgUfAcZDXD
/QHihcIr6wBj0/ToDueLL0f7PmABwDDUpH2Jq1TSOvJuDT+f2N5my4Y/QW0F/Om+
3tdE/zAuuPnmnijT+T2YLKx9r8hSOMykrBHTDYe2YTEMPo9dHXA8BjeNYz4BQvHy
i1VnwggzEvrSF0Xd25eT885mpViolnFPmQxlHLDysRMoWAQnRmW2NF0g56oH59Rk
VgRUQKyuDrjaWPEodxyOFcs0ah1mtyI3ULmq0MwtRCyF0/NKW6RpvM+Imcz6wwMV
1/xT+FtK1WIhy+JLNThur7vy9hSYHTqxC83usfp7V7BGo7a96d/kP52KcU3bfW9A
rsI3HvoXA/ZNOFjR/NXwiXCayMOeFQN/Wdp8YeVewfCg02ZA5JMZT/eIeQ0uD2Um
bsPvvzj601mzYbC7q95U7j6i5MQD6rFQyz3X+BMBEWj6WLBhPZ+e17QuKxiHn4VN
wPvbTkXiSgu1HR5eryxWj1ZMoxfdaTns73b7HTm4E1h03B8JF9fvhF48y6kXlyMk
8UFLEB9OJR/KAT+EEh5IdyxrMC8cwULimrPM3AnCVKjllLMvRzjpCj8vydKMolk3
yP6UH/qhmYAYY2lqGiy+aqf0SkFkGCR+usZvaAAfWBl1jV6u7iq8coJggBFeXBrc
aeEk1lXkJaPLpMBrc+0RDgcZQsL8zauBSJj2fkI4GpHf4G1jG/LBTDPmiiDc7Dpi
mzPvd5UB1vDpONf2Z8M5x8c7L1UTxSqeq8JwnRVVahw7/7FjnqigEruXgAcMI759
1lEtAosJGrAEMv0R0ko4LkmAyjR1lo99uh7TWmPwPUrzPfCUtiPTfNsN3dCEc6XP
SAbW5YM84Bdwzdksv5BTj7eNgBO+4i+qgaLuZ2TNoVd9WHGqgoHQpl5uB0x15Q34
xDf3/tRPPw7GnnZTgUFl2srGYLAbl1Ny/N037vRdIcFD9T+o2wyYC9DFro1umQlj
FNXuMWhcIlmlkqXl7zUqLh8DJW/WUvKGGnISz0d+b5F7/kufTTudwJnSxu0iJY7E
VPZh5v/GlOwlSyrdZ/iu/6VtZxI2wqiY6aqhTa3RMCb4ZAF1DSzssQ0ndFggXHJm
VbyRaoABKw7QLA2jONKk28dxan8S2tUWzWfI1tg647Qb0q4PlaOQpGsQohJmqyWy
aawD0VHvnmdmGGfRzkE5uqYQcxmPyW6lJ1AUzx+lQ28X2tu+EnZxh2DRSdlMdaXO
RSe5JoDbk6Gt5Ix0wzgxUr/nbCg8bNvejc9uqYHIszZ1GoW61qLNgMyrL64ohoap
XSCQrziGLCyFxvPLTmHfrA+p0uZRnXwkv/DYHl+J2kGnS1uUM0fFaBlgkNZenjZG
0XnNYQ+4D1a6qFQ3hgO3ggTvc6bPE/0UmFJPSpEXS0oLpEs3WTfF3WmeHGX0Ss+M
8PPawPr3T+k46dzljyQgN2Go19lY96YqTGQkDGo8Ib7UbYCy8pdBPsCez1RQCgnz
ruSI6KDdaV3OQh79Hl9byTTsF4KFhoTIYXDlH8Fp5Ie25iMPbR6KT8+wY4n6Q0z/
ygo+EK/ke7zrkNbUTP3SzU3y1ZAEx31j+LN5P0woG9YB7Vdf3wZA2OOHIb+9JUHe
AWqIRovC6ooaUZZDu02DIusqrjhoLpj1EMkot8qeYgcxJP7GH2s30WKgo/MNnExv
D96r4qPmgbgeZJIiCfDVrWDEco9xg5h34Al7oNtlpa4dRu2YkflGdIKwEGqTdj21
zepXcHGBmhdyC9k8KaJw1IxjKqw2qly4UFnhXt2k7Q849wlT67mFjXiKVxxePpof
UngJqJneE2Npsz6YwUov4IfsNnBTGpYlkCM1MYk+O2dxbKFx1w5cXYwMbjAABBTz
ObO+C0nBG9pkZ6sk7rcMgTw0Jg1Ri4SgXxbs6VVm4W4Dzw2z4w9kCwoDxItrU9oY
gRip/jfTaqA8b3L31Fs9ESBKZ2CmbnZDZRzj7c4fF+8oBde9qZM8FbGHriQboVAV
Vdj1N1IJc2MLE/nsS/Y3RxBzkEVfYbEsspJy9i9FURUixl8ZIQVAd5ryBNLWfvz2
xDQF8aoKy29KBBAEdPzQMt5MsPXkUhZmi34IRu4aWUnCyZ+LxoclwKMRvO6MthwL
0Bqxh1HsIwzL/gzhnJZH/WXzjU1Av7fpfoTouSqgbN54LcZG3siAxxjuur7FLQUk
Cuyd8il/UmUBoIp5O5i0U0QnD9AF+cowXdzrGxUZuXyPzJvHR7Vh49J5gc6u/ieP
FfJrQN7xMsjdd8CE6x7j6+wnHg/nQ3Db0dtPAMxqnfSDIo16kc2XE5bcgFRNnPzR
sqZ2kBweu7OnI8tdQsFsXKdtaOD/PcOEoyZzw5Ly55RJ67AVYq7Rpoh4XVJTl3LV
NYDJbVTEdn0BhXbbs1kGs5IGDqVBST3sviJv4QyC9eypZkTqVfbIQqXquzhDYzuu
06c4hunHCfMOtJ2Lez8a2mam5JIxY30b2GlpLJR25vrs7CLFKHY+KEt8iSHPuam5
nCCf+qjUzB2gFSn7os2mmEYleXVG9YICB83Ip811Y44qDwhKnN4maJaiwnXR/CLo
NSJzGuhorrurXj/o5xo4xsRY9IMN3unrU0iW0XWCSEE2hiKKIZjmYyrBIGMI1Mwe
8jq4rq4f2TR9PXPCAvphwdtYDwLl34kxatZhccwH0GwNaraeAvSHCQmP5Zl7Fjbj
antWVdeQUEN17O8YfyAvB9/ZPSNHY6NdPdhI6bkSuhiTr0Gq7igemKUtb/0E6CG9
jU5ut3XDTB2RzBH6tuj3VZ3zaykqhOIGTkMpzHM1Rn90tehr9aVssJXP2vDraenp
d9GNXmFSehKdQdfpheOardgdlV9YXf+mhsVovg8Sb7BCz9WdpzxXjs4EEMNaVzCy
zTOQG2kfPHSP33k4ewJwU0zRUsMsGUlh3jETpTghGWmbbXSQW6pm56DgHPgLoO8x
Ty2vmf3slvYNYsRYchJ9VPLERqHNsABaIubF8v963tydZWtKPvOq7iNKbVw0/8/s
Vp8BVme2l9IW9d7I2pnChk4ntNLGt8KUHbsVgSPYiKY/h2dsg3jQ3RK2ROnq5Wg1
okwgbbrTTTGtOGsZsucozEt/fWavSPz/ivdyN8lpQi2mTkCgnIz2hpGoSuh1NuNL
LON9afP4xVzQN8cr1bNOVEJDo0sCvKbG1cSJcxNycmeaCS/wdevGG6c1leJxAQ4d
EVGtzlYHux20Do1mz/JaN9aKkDu7b1JLQcQ4l2sWCNheB+xRuZ8KtqND1E6mnrx0
sJ2Wuqcu1ROVIOB1BFYlZOtHe+1cQzWodcAnbUzIhbfHapuFlLr262oqxbWNmdxF
kR6XrEyiaCrroLBlEzmtxC3oR0K4tORqt3KhLLLEGk+XsheTzqAqJxSkcqWd1Eon
+olfWLG+pHAFQEmD+fVGvlau2Inq+0KWKfOwQNIgLv2OXB/1SmD7vW4mIOdKYvQg
g8LPGfptduAagfq00wQ0q5tIpUmYc7zcfB+XFgj3Xn2T/+gx9Ma2ZkvKfNe/3Fzz
fQNTT80FoCYOly3ZgkNu/mO4usN9aD0yx7bQUJ2Oz+Jbe4O0MSz030CRpcURG84R
qxYKhWFOeeea1cnwelVKSGzFulNbeDgpKDFEVxe9P6r7KvjXYV5wYJYZBQdZa9Rq
BPdG8Yxi9hw8VYocacqwlbqTWx6WCpM0bnW6Vw6bKtc2qIv60djgXGOiWEJ5hdrN
4A3V1UuMNTdjAdxYPaF1+F5rqOpciMvB47g4NTXcbsCQJ3HkTq7xgXnrI77/9brk
cyhHza8x7QJvjbG+9ipvuUSNM7YvOxMh4IPz8rZZCuxk4TkV1sMvRxUWtDV+PX0B
/P7RQAtG+ygKdlTFqiI79xI2c5cbIju7dUMvfvZJpFtyjL7xDDR8EGVG+Xh/XDnd
uBe1rJR284Z2Lmj9MyL73c/6XxthffaFBGoWqrWctOODtoOq+cuA6ioYWRrpabhM
fDm36T9YeSYXILRDoY/8jmWGICBoWvPGPMN9NoekJ1ykwWkwq7B7x/EqNLrFjaXs
eesA2Kg4Rm11Cw1iHdvSnrYiWM/pT+D6+C9US2EwOOTtJ8eexoLwYRiII1JG+qS8
y9fEev8m6xIcrJU7Je4VeuYI7ht3CjJPM4705bszuxMCZPXhzYM8eDtU6ClCJk6Q
Q3KVpWVHE1wy3vnZFsTmkGcOnbGgzpyQyz3YVv43UDBIA3rDSR2zHsDUomvYV6mz
e3MnvvFMcE/SMbfZfDR1YxRxK25z64CaaqbA/U+sSiv56FUi7fC2X/uaEH3hGVw2
fBSmbc0QwEN9IkrA6VQIKCI4zbzyxqyBa/wM5GR1J/DMhxS3BHLVLMamqCDfpAPm
oIltC3jJTXK2hHXQQjyAa/PBhdVTjJxLAsExa+B3oU4bxSz40jiYEIlss7YCm7OK
3Pg7EizrQiFZ8uJOWCrYOSH8EQWd2Zx8Dla3N/B47x50oCTJDlEjrMfm1g+IBbv6
l6HY3F2iTk7PxD1S7sNpILwM7swDEgPZOxVAKwpBULIq3rZolF7AfemnMYpVAfa4
YzTe7Dyz8VfhrxEB29ZS1MLcmAhz9358SXO2c97zAMF6bleYZRPUYlTEUVKh9iIn
FP+cMAIBH5S9ONLPPEzAn/Yi4+u72ibb1VuC7M3yrPWaMb8IXmkv1DT+QWbudKcZ
S/Ip6yMR+0m3Ldy5QizBHkH335SFw838Q/LQ7ASlQ7WeVx/27dGZTWR7GL7VTHcG
+oDK3OSRe5q9CNSC8jH0nwG3rdT6yUkqKLeZdoe9HPf5u2LnhyYRKdbelltfPXnF
EIZtcjnZrH2wyfczW3XA+MPsivlFHZ7Exy6IzhkdHSRac/1VZWM8WbQr77ogco3a
/HKRAbZ9dpqmzQCh97iCGN/yhOButGMVDa0WRxxFYP//Dv43OC0iSQFCvaP+IHde
4UiwbqE6hjyzCE541lQKlpDm08lC+UEaHpkjk82zj75c5cxViYPLDS8T+wvVR7ZT
gRViSNQbQm+xfgoqSN6UPdhymP/9NT6ITPpehvU+xTTI0/baE9mZPsk0hMgo8CCO
IEXiso47+vIBUxIUjGoWNrwi2VgkqYdfnUfcAEwRwi2ufT9vWCSbfE09PSUD46qB
u3bkmmfM8scisWT+jvJna1k3aJ2szBMcFqBVD18AO+a+GVi8GPwnM6x4bETMTug2
D52fjrCW6UTLXTykWp84ic3K4mZPu9xBaW+UaFBz0TA9ASZNPsno4jxDVwGzw1T8
tSFKRd9GuwNaoc+uBjqbOL6B0ma8s6aid/0O99wk1gMFg5Kjr+96Lg/KrvLa7vEr
E3ZwwJvOJEeSZ/fFl9tQ/phCa9LxgC9S8BIuZMmq4oR8XXkT4XxUWp2polg/3DL1
pIGApoXYOexzfDKR33cqry+1n5C+6CaKvqEMotMo9ZSPpcF2ToAQQSsCj+TAPyqc
I9GewMluRlmyJeh9YP0qbdESVtoTkSLnpPZRD/4Xg6vM2a5kGXJUeS+CXUSJfPge
vQuazzC2HRR/UQ4mLgspNGLPgpoPkBSmncXwImHppYT/GrIPLHXj3n5FVYXeKXg7
hLIjjudlKQviY2AMeZCyBh6tfy/ECIsH4lmw7G5xR25p39tvMkx7fpYV33X5OZdW
u7KwUYbJvUb1TFXSW3IUXLPX6vYhXcKgJE9aT772qX30Xxr+ft//uyjXOxtFv0S7
FLZM/X2KXYRosdHO7XdsqLxsYypCY3K04P6ULxQUpJU0h3LKO5YDpSPIXvkyd481
7j8bcFuws6E2clDBO86tka9iXRPu4XVdm4yDuNEFT9QZZmkE31Wob68SSsvFzHtA
th2RfGYg65uBTWLrh45oBGCc/oVyJtycEoGwbBTwgECBs9fatX5GqIhkxBeVbsWy
NYcsa5zOVxBl40CQ2VgZ0sIvfv+usqUVtmyn+2L6HKVjq8Jtw+SVGgMMyIGZqRnL
+rXWNxsvPXQhE1d2Xne68ZL7nAOxRAhWzbkQKlVegHiuvIxaRiVe/jzpSomxwz40
K9i/jOKZgCwx0y/5Up4d+l3a+8be3GjZjN4kqyUd3fudwNCm7DMleNglUoHkRdB4
Bk4J3IGIHkQq+suzOwufy+peHSfrbmzPBrwmEArL0pmrt9N2Ctl/hZSzY4edWJod
+5CJRfk5mMKe2KnZSiUfQR7iw9CV6FsFISk9aimeNqVxKsRSpe4X/A9ve4YbIkgX
p1ccrt7qpYnR6LXGRHiDnsdcPjsE5vM3VTaxngrKoM52Lzt4L3qoX1jf5l/9yqie
FOt4rYYfpD1sXfW0B2vcHljU3KcRqSQu7ru8rizJEe9ChYngXgKGwMNaTHlTts7Y
Rep0XZXG1My5auqTG0U7Pj/gxQ8FTWcb4hIdy8SAFwCI2xldOwfqgiOLAcMmqpo2
U/itQ8ldclKnbmsjLZYVLeXLF4RYJlZPWNfEbR5DdhGdIQ+pO3TWo4crUebCpIEF
b7ZpfB8TLK2GBJtdlBVAkpQGFUnsCUBIehyZJRjanKsrUZuBnkGvEVtptrCtvHTK
0AsEZdD2QgOfGeVHtAK3FamWSPd80yepjc+5nhFNXZqNNXbs2NExZF5CN8aJYrKE
occsva4oj+Pn7BXC1BMVUzCaYBE4ANHYDyNTAWKntLDKdlRvFn25HOmV9xOqZ8kn
/tXH7iuwRD4TM0QhJ9qO1NgCNDfouJNWyn+GZ/FG6A6Vd8G4MzXaTX7X41brciAt
REuyDjrgC3A4Oma3A0R8sZqH8DmoFcWEYqvRKYqLBVNVSOHXtAZro/xKJVhDxdpj
KGbKOUZPQ5V6yRVfCJ2jS2O848Lcr6G2QrNMK75Pr7xkaHMaRmsXaLFxVi3oXNpp
cf0TkzYibDA4Ux7TcFnH8Cp3gyGd34uA4f2jadar9vVFN5XhIpZ/6PX7Qx9s7PWa
u0e3YHNzptcqiMFmwIgNhB9y+xRKK18KhmPXtRrYajCPlxxS2j+MS7NbRX5VDS8M
WQaSTUh4fQuJJdVyPeMlWjh5w1mpc8YsJPBFMs3kbrh/zqQF3KN8ffC554js6dkx
bLPEzW0gfd+iUkY1HOUPrGL/sNBUEuL0n3Pc+sj4fH5vrNnWg5bq2cbtHo1Y7Q6A
OjVtJqgbv/4cPDILfojbESTs6Iw8rYHHXJ6IV44Am/jDcR+Kj8MOFpx4nyXpa/yn
LVgiBhtKLt1DM2LH96/lN08UPyVJBM84va7UAVojqGb/OK4NZsYMEKZoMS8Dsg0t
3o95rT9uZEeCsv7JqYmskZofl/JPOMxR6riD+n9jlpOH6JmwpkdfB8zvQMGpqes+
V3N/xjGoiGdVYWoeUnO2wqAls7u92kp1OtfwvSiRZQcCu72xVsAmTNSmMYvk9Xqm
wYBtx5dM67sJCNXMdL7cxh0HILP4fnHtHwFfDQs3aHFNPaTgKCpy0aYRBj1HNbyV
IBlE5NE34K2iIPxc1qhWOcS27Kk2SqYtyLQ6kF2GadpcLgPdXFEZPKa/Tymk8Yys
a0mN7KQTLr9cu0Mvel1lBJrP3OyEIwNHi9/jWcMAEcLYQgGsUglSjiauUrdXWrXq
U3QGyU93U2GPMEbaJKGh6Haa4g1TVK6EbvoUN5Kzt0r9QLbTlVe8wDiMnGHflNUm
1p4b6mjSweaao9wTNfzXoQTtJs3CRUifMekU8sjYTrNusRvt+xAWBR+Pnvekfbl0
10+5uQ5lmH7m4TebzZ2KOPhMwk9Mjav4CNLD5SafKFH46x91fQT0o2wUcR0IQBAi
77CKW7uOP3waU5kGAD+CkUAKWxalIhB4kN7b9abL/Db+mZsYJHdDMJjxiZzmBv3r
m2YCfyVIH+ddEVurCWEsPSGr2apj/1w+MitMRKhVAspeQfGVdCPLYYdCLXxSVzr5
7Bea12t+kbG4FLuJP1xY22gP4J/l+L/HL4jxd0i2h9iY+iCF68WSklzscxT5zzMF
AhG/yPcphpWm0zi+xizpBbi9hdORU3IqmIHcFGl39lrp0perFUiXrX180VDRnCqQ
t2dNtNjVDyCBZ8du7qeH6jvwNvxVBGsg1js8A5ISoY9jBIPJeQV3kbSRJOlpJCX0
dwvZo0etZWvs9uxNXpBeI2EnOUQmf/Rg4VGAKfwW+hKuVc8ciELvHK2yoxx/U6bo
AFA5bdLqgi+5LIy/UGpJjwzWAQ62ZLaDFYKJlIg4mwxtxW9oqygrQE2YEslr7PJt
J6rKUCxxHk4TKMJ43yhfbErs3NCcYwnJdbNemMRKo+rcw+7RU/e2GIgMhcieydah
dBryX3bUcwEgl3lRYRvHctn37cpPWCITlR0VMvwDHG/IpU218nltTBusj+XvWDgE
O7xJxWnwq+R2CrHoToHp1QN8xb7YwTdjUWqEfYAPZToQ4aw0eKdYLKY5yQeTMvHh
0lRz9zc1pANXQcw2peS48be8DKMb2WhE6zieoiaXkHw16BbQ6jfBWnG8KXtFKotZ
7FVvHPkWxtlXgbtJYZe9mE9NVHPEFYjziwMLjFzJLdqW/5kX0sooT+nl+OP5+wBt
MJeQvygXxDyrjtbQ9kQJbzued4RdFL2u6kRCxNIGeTOEgXKu/VFRoHYrHICOmcGQ
SLJc2QRQ9TFIszTXWurrTON7iKCHkjqryfOSHHi3xDYKCEe9EVx/2Xnqs+lRyRAz
vFmfQ5ZnXpkSAOQEQM0dCJMReKzBzZVk4SSAyWQKSitHVo4Ce7SMQ8MrJTcBJq8p
DY+gI/1UVRqwKwe+kiunZoMIc3mNpAPkee+wNtLLeC/XAdjpX7KIkjogLkvim1Pd
dlJ7sUnL85dmLIErHOt0SIg7EnXcEgqwzbBlcC+JGGxoTK5re4iA1MnBVsVfIytf
TKyth48bs3NQDsT6W5+PcSBDwv+i3pc5iVmdtWO/aOwnxe3P+3BwGoU3L5EgY/j+
Ly3beqTL0Sk9E1rrZ8wf+m+tDNBWk++TL/x47zsXXlkcH4ECBQMDTEqCBt4KY9Lv
JLmh9XfvPuIfYhr0h2H5EWYXl8xMqmAcrbEOJuRU1kDixpUyQHu32UJCKHJyCNVi
GqicyhjbBfteWFrwZnVfWcvCNHUhMkDHVOn/yW6MeSOVSprbeHMNQNOHIVZJE8nl
6dEunMLo8Btvf80ihr62CSR8CI0mMY8HwO3LrcH6bj1RMZqDov5Fnp+OZ4L+HazC
S+3mDwgagrKWAb5gGJEdT0kiJ4mVkKWJDpetJ7Qd+tR3sGnFr0WzvikYH+djSl2V
c4DoFi/vKJNfdwXV7UtHtEfHZasngK5ySKN/PVU4mTAmOaIuwzoC+67km7vEVbUI
uETWYPUELKFi7FTLE8/9ZbI/i/wHbX02mdqPIDfx1T12EOP7btLXrqVk94Y0Pqnj
9kbs/anDHuuWm0xgxPgMmhzQkrx0JGWBLS7bdcpTGC+eFpJYHU3H+r4FGmJJTX6p
EkYQ26WEeKpfVqYwhYe3bwUC3caDpcSTGTMDDTRWVKgIewwhxaNvv8dWzh1vveNO
Y8slYPAoCYlS+dC6VaxmD2oW8GKM//kLjpUmIK+SmJ6jgqxjC0hdXgQ1gwTeG16n
XvTRcwxktkjvFt4z/lYWmxtLNgPtDkbRKCNikq9/0z1jOjhRjkt8QmGnzlPAfFz2
imO0JsMy+SM7LwO4fDb+wz52mVGWGAVcUO+F+PLE5HBd35K+pWjDxV4zh127FuQu
y6bYLFDRXJvdyzDraWHoTyj1b5NI5HoyhiVzJL/3q6jHDHG8ME6Vcfj4hraF4yMW
loNbsUINCt4ojCpz3WcRqzz6pBmubxg1eI0XltU06YSyXcezNdmaWnsA0/oqSMbu
HI3ovXdO/W2/nHcNEemk7UTLjcJKqlfRsUcmYQ41NcPnOlgLq5MVro+MYBNdo6MM
5uVwRIdNyVk7FuRZNAJoDqTMoq8VU511Gc/ENWEHJ2WHSPqsnixRkIKkLWv+XKhu
aw6nuye8QMZaHXwWZAuSAFwEz43NwSwtnQtG7GCL8DmTVdC3y4yUpu/+QCKdUlhy
VKoynC0f10xVkzS/1LsGwrdIBeQrM5aZ0SXxNx47OKYj40jgZPHn51Gi/5pMQQ+y
8KjvwtnAcCyH5YKRzNKIc2LeYj/1VttibO1ZTTuN3ZXOeKtqySDR3U5Gu3w2myB2
/TNhNAZotFqH601FyVGAGdtMX5ZpFOo55y5WscY86POPIvhCNurhK4iAGLGniwrA
8RHECdl71HzSfh91AqGWWXXzDO44w8ikdi/AeS0maBiZGVOYymb7rywWlYocIxog
SVvh5jOGIggpeYi07Ia78kZyrOjZmFPNnH9kO04bb77wtp9hU2dm2uWFE4B6XHr3
yGNcfpWIzhtKHZkR/+KowXBRHdlcon6+8LC4GF/snWZyFxWLGpZ9Tn3ENEDmBgEI
RPvLljCxynfvQiaO+XMv+EFE5qFAauvN0CevD4t0rQjpQwLX2cbGeMpMejFKflOp
3Z46xr2yWpVMzDNE6HP4HGuhpwJ+1V0xtIN7t1FAg3B6u7Fjcrcw0Fhc4gNmdDiM
Wjx3cAQLNmGAGweCQofbyf+22lgsAfWa6gvrOUd7WNhG0fQ6yJfkLYfwBhVqageF
CgxD8+7a0B9CplVtgD9Z2oIkSc+8Zz7k6UcmmEBQII3WjAnXZg3HEjE9Bkex2la4
kr9WoHJW3cGLbYWvzF3tEbVilCChQnXGw3SzngdaJSpwpoIUqd0iJK06tbtO/kYJ
XNtP5VMosvg5bPW8oICE9S3hXwzRhibqGRySHrsp1I6eNDsresbMn/2q0A5VQ2Wz
8Wkm2kgCIX2XJfN8n8qCJklJwJce1BfAMQgWJFVTVKJLR10aijrN2V4CzOk2dlLt
1KnVcWHnhUH8ZOj9ya3u02qp7oBogH7sm8W9Cwi+t0Aeczjq+PkLU7/lV9r7wyUY
pCjethB0hxZgLub0bwKbdr1g+rGaNii1Fryd00P+rfZGeQRXJEfUcSp1RhIcP9tq
z6bzASHAHp6/o0F2f8vuAJxZCMvuZX6i7vtSxwcSGc1o9AMMEjnvzQoKIN9ubU1y
23Pm7C2hNbeTriJNzraDzqNaeScevigLloPs687hQPQ0wQWH2m/3r9mUfjQVAwnk
HahBXJIBcpAIqMSt+Mwq2TeATr+Hjx9bSip97eqzbPoM787noMtoPGdJOM4wzZSd
zQnxzNIzfMFDTQuYsyra/PFFgLo1BuU7OylU4vz9lVdSTigv0xmbAV1VUQyWeihr
kW0A8tjtNsTA5Qx699L0CxJPLcuZCICus28GCRNhCJYdW6vjgTRiSBefT2dd4fHT
T27ulXjat1NG1GlvJkdtXMMaK57NS7Zi7wkkFgfVkkZZj+E+xIqO5dXjmvdU8mRQ
8X1IfDVs3PQgJiWDnLFpN5tZ+VkyaMexVZAOaRG2cfGjwTZh5TjJFG5u1kckV4Fp
/aGY/hhPDg3Otdb7qiUTrT4FlT3d0XQXF7w1FfUFIlF9FPn3zPWYmGZYQyy5Thjl
0MqTteyBAXxv7IQ2hokrYPGFGCLWs69Hwf4bi6/vSTB1GLUTY1z5wezrZyYp+3gc
YNZrLtwkmt72kufsIz0TJ3qCXI7Rk4fZjYcvEkEmcBJyChpQyssDZSdAmGS91/Ot
gFw9Omudapc5FvrndOVb0dUi6C+EsSqtvICQSO858XZIY0pFJnTzuoe9c+PKN80s
o0Z07ZA8zKwtv02IHMdCA1v832QHI4j4oXOQqH1IsAPpKmIydSYGirGBwFY2+nj7
ULkidOFMeeocuKI6KF3hgFyzB2zxsIWGl7Av2XR+IBmJmhaDxOrPdkx0PDpv3AKp
V9QbK5tUdjSP8WfNpP0hCx7CTEaqSswRqI9txKdz9Wa6tv5s/0eiZIqDxT27dh6r
QV8ou7EMPwcm0FM/WkeoFTTVTJZx3nMC0Ri6QG5spCbvGw32gOWHoI6+SrpvJMRO
YBQDY0Ddf+rUGXGwECpdOTIvlPcJXw9QBWGsQMI0PioXCEb7VYhbf2n2VXkZ1ikV
s1Apl007O/Ofk7wPeZ1lAh0AtoUm7Ba57Fgei62Sd2n5PKXz0K0tRaMDncRL6UqT
6eoXj16uVlkYaKxizRF/W2+ABA1XQhxeZ442/lmcQrlzDfPHy8H5noq3AeHdCA+Q
PA6pk2CSp3uIL/zyMOP/yRy70EEwio+MMjiw/G7axn9qdpaamNu1vboekHfn2WIm
hnufSzMIBQo3ELNdkM7LcnKzB25kadJYdDpLByvj+04DInjeJG5+Zc+VitzECdHD
z9IhbOwBDGwU0Hfrzfnc4UfWWyDlBy5vQOZYuUQmrzgSLTheYwUVoUotOMUIkHh3
kT90K7z02t4Gsu/1Ls1Y/ONzueErGP8fhT5v1DLH9r56nLyOBuIm64u2QtHry7ik
8dXiZuHyavP/TH5Unj3skfHQ/rMY3pdWZIxQg+VBjHlLVuob4o0/xME9gu09y6iE
ix90qH114pnMK8aDtvvM7MJ2GggSNcTn45kIaecvwQTaqMmYGcNCEB+bTcgVQq1A
NWyP0AVRBWEYI93A1rIM6xVk6+B3XqRQu8fgJ4bYuKOr94rdHjJOFV/lYaJD95X/
BqupNgyzY3z2KxyCutxCJXlDYE62x502+CsRetRffIe4hhlqGfqPW6Gm1T5zTaKb
in47DRs+C9vYl1wXGdxkchip9gymdbjt2d/GsXsKqGX2mkRcAYt2w0m2Hw2buaZ1
wuatyUI3oXOrTJSHtakWegUeR7EQgtdSTVU73t9ej2NTYGvPzbId/qkZ7yXn7RHH
A0rTgY4BkxEA5H01PSOKQtgICqzWQRo/ikxEWelWXdVEaan9HVnPTF14sal5LuA3
3wSJ5hb/T5QEW7lWmkbja63VD32TLM5nejA6h+FziJx7Vp7gpwwc+UuJdXlSdLqh
JFbdluw6SssdFTt2Y++zZUblW4MJl+l4+NBHpV4TGpGCFN6nEmctU1dHbVfKrYnv
mwTqlRwkulZ8EcSTbtZzEuLDNvhJCWXCAZFfo6qcFYHkId+icUBs53PiUlm6GOIh
e/ft7Kz1nbHZVLHSOmGsGH6/jWrRmKJW2boYi/87EI0gFjh4+R4EWNdxQbZOTvwC
YL2y71IBp0lp/MTyJ6YIDU6/4df7/tBQYwmxqtBfHArcAcmXmE0u14G+DVtQfS08
JilW1XSmvYsgDfK8KneRNmjI1xBN0tPquANV4qQD6P3nocnR9L8tuBEJYYwg2yK6
Tbg6P9hVynLn+hNkfTouyzts1LnhkAsWkKBPIWVdpO70QJHg4Yd45RXIaTni5bLA
wlDE9WIKdcHsx8N69V7K5ZXIv2X4BQs+mE0pQjMuosWEPYODoEj03Q1edckI8yqT
gMAeHat0unn9/KNrQkn0Ne02Cj5QZgv5lGweTlWZ32ttkTwNimLgr1T/LX8PFp0M
PmPQ7lgv/lI6b/PdneXM/jz7gZbGA33PGrAh7fwb0hrwYcOVDGd6EAN0saFkPnGy
Z5JDb4ZU8xMb28vKnwjplwVjwnkG5NdPJ4Nw7hYqmzCrtqFKY+RY+5ncGKEYI52q
Pwg5ihd6+EulkwUtKCBip2/ZxEpMEKGpLQgsMhHuO/jXH2Z+rp0z4jxurGTLZbeG
ZQKvSy3ffX9CegGc73lMwVDFfrisyzf7/+/KbQ8SJNQOStCFbBeyffLsas7fvNM2
2PXu86Jo9ERewM/cjlCk2EGp0HTDOChjvgYzFclaPPVZc7Gx2sRjC2lJpA78HVgO
jAFkR4LMOjzCJ9tMHQCCW+hstZ6ZBZYQ5th9bN0UfA8ILLUF5aQuK5fWzq+OcIhM
TqVZSsaRi4f2stYdVexYBd1BIL8M3g4nrggSV77sU/3GJQT3cCGndA6ny/NMMOZT
3ZV/BR9ULt6Hj7wd8qQhKgh/+ArGkmH8of3EjYbfy4hmCUDr1WjxwMAsU2mA1w7W
7qowWF4b/FyP/W0WjGwfDEg3hsb6YvDR3hZSwGN94kI6C15RQcJtK3xZkw9VGCI4
SDg83L0K+9ShsNQHBUn7fWoIz0xo0wFKd1RdShs8AVvoFgJGMv4e1gu1hgi4YjLW
UBQ8WqPuxiwl76acFN8tCTQM1mMpi9PRGHUKLS5IXWB0zfQdwZ99XJVCT63XUzS8
i0zi0Iplg8cZfD/F2LXX5NzgolEIiKBGleEip8awnr25tu+Wtg5llNhz9xArzAu+
TL3x7/jdXPAbyfIvwLkJMIbJpxuHpzheg5Jixj/M4zLdXgHAhUC0jb1KsI521Amv
0R7iCXVBhhyNvesxCeGwWdAJsJUJT+zoBisxNcKwV8xlUf3dyoczsLbb+W+NJ5Rm
Ay9R+6Ug2Whf9yFz9OebB04iW/mDsHsdy0adOQsqAcgYEJ0XPxG/mNJ4emkK3kW0
D3IA0ojQEoekXrDtWF8DdeLVZ5dENFIvklgLCt0ZoLvd21ex+0ivyml32yGshggB
ShE0NpdeG/IcWqBYOCP0L06DblWLqv0P7gFT0Db42AeAURb+tc6/t0xeCWVf+5QV
AuGK+keJQGT0SvUEcG5jsKoj537yUmCON2vTvrIpFMs=
`pragma protect end_protected
