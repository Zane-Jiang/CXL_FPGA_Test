// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TTC0ETvsvoKKrPUfyx6KFps1TNNjqe/W/1XoC1aTYtcV73ojaAjZtqjoQXe/
iEWzey5PIS6/+wEzsd4k34JjdnIoZMsBaVgfB9vPw+GKMsSyxPuj0p8Wj0S6
ULPaiaFrKnl8WFrVZLPZZKfDOpd981NvoMcLLE2bRTY4Yk8CW4laPuvyB9IM
66IeCIMw8lL7NoG7IOwYW01ETYHwnsSXh7+xPhkVt0o5CCkoQKmuELzwJfDq
OIaUPtBc/8SoRKNYOS7tuQeIf/nyjmgBY+bKuYMO7O5199kXgdc3XO2xQCg3
6n7rUBdLyQNqDen0BWAggLlW4R9GFS+In2drRaZECA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BWBgQ5kvYVLV4bttjwdi2scutyazycY803DfHzCt25yK1ropOTFqrcNqBAA4
NQuYdUEvVDiP31FG2MBvnyDt7hOeOryJGl0ciMnIlJFgR/TNskvAGZyVwl/2
XTosDjtT3yRbny7l+jJI1FRON7FtZSqf9oVseZM6BKuno92JsPGMroEFbX9m
fpkFKI+K73bXyVFkBwXg2TDxadjemZr0WSdkAIzH69YVyAppjM4l9jIMyR04
CBcuAYv54oHyj9LSgT69fIQ/cM1qhpWBeaLXQGHXdlb/qgQl2MpkZ9beM4AP
ZuJ6Yjjo9B64l5zNjzn4B1Pf7wZGWJgtsY+BXBnJ3A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o7F4I+RckiIL/lMZZUhd+azZL9qJzYN74/U3p3tZmQjfkgFmTh0L+DotL3F5
TdYyTc2m5C3psFD7vFAp8d14VXNyByQYHawyHl/xMmVROkFxTlTP20KAahAA
K2AtsowGFfakFBnkTDmGwspZQ5t3Lc5kb79DqxkrLjLT3SFspLbm+Mx7GAGM
chYAhA1DEPZkfwPpSlu3/nvstGgxrKmclDjn3v623/f7NQV35k0WnT+WdrBP
f9yiWbqfIP9lY4cO4dpWDymz+mRfsqGTQobqecrNwa+3lwbjt6AuYTwvFNxo
hndaIJHqUUabSBDXa/WpVt1knPBGMJUP0qFs4UVuNA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FHSme80C+Uq5YIzQYPR5OZradz99PpgCeQaRJHCNTHU5c7ADcZsakKKE+rFc
CMY9sB8jmwpy3C/xaLdDlh1EOzbl2zxOrpBBnHswhQjoczZxPYofW7Jr59xl
x2kGpEHZxqKorcK/sFM04Alxji2Qha/T8LhyzO7TrAwTmmSufpI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
j8GN3mfFbTpRotgYKrfyY74XuoRbu7R02yh5Dj8GMaK6wLKJ8ThuXFyZoFgF
jePP8QrpacHPYPVNPn6sUZDjKG/hwIpHTTguS0nKf97MF5sgqHbf+43d2Myv
5EqzPRczcccHu3NKuX7P8z3AigV9jHE+xD6fA7R35colZmQot+2c7MHJsj8P
URo6DArEdV57Hib0nt1stkiOfgp1nEwnaCw0MgjQbHOCo+8wE+VOrHR/OweK
VzFFWTlxCkVecXAfMaCR1l38RFZIt6pyPliNEUwQoKmofyltVXLKRcke4+fJ
3GysrkMMDcvpAahu90ShbcAssMzV9Vph/exdwI3nQ4YXW1KAToIypeFpJAbL
0Jn+Cc1c77T72WmBlsI+mWUckr86BtJv7u8gYrxNwnavRjSbEzIcWfpSrtyg
uIZqsEw4BujSIhFsio09Q35zAsJGPX7YMFZmcA8RqlYg+owxcq5R5aoLs8Q8
IWFoSto7Bi8eJLgjf1c0VD45EROe58sY


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RCGB1pSWhT/kB3oIfDSsX6Awrvwwc5Ae5kpNesiVt4UOwoSdyshSrMhL/upI
Uh2Ww7ZEJAcDh3FGqstlbrSAhDBNuwAWV9/MD+r5q2IbRDGKaJRyOIhqGVnz
k+hWBvvyyMdadIv+vEu3jH36C5nZiSBwUztghIg5Idt8j3ubE1o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R9tB8Y1UlhZxou5qxcA7PSB6VPWp+DVik4+Dq5O5Hd0WU/aEEmMWEX+NiR6O
LR6FwfrJRy7VxHlebrKaCYi4N+HXTwKrT6Oe0oAij2bNbL4tVFdOU2hF0Xzc
xwPehlksu3OxGxAZLAZ7PWv+FfoxnDkIS/KOPiF0ePw/PvgRvxM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18432)
`pragma protect data_block
OUYNhjM/7qQ8scQ1oRo5BBIRsW04ZnD6LXUwErKZeVWZNNfNvAwLGRS3s/Du
WrghtDhh1RYu3Zqo23wRVqLYWS4reHRk3IIVfOtpCEGmIkAIt8EnZIOogVZq
Hsuo4cBLU8M2xHy5GuqnXz2PV/53lS3UYDVTY3SF2n2LX6+3jd1aeN9lD/Kq
d/6QhEckPc0DndovdNp1JKNdNzBva9gY3agJ8lUKxdTa4TkDCvt1f1s+ZIAZ
UmyzCsEITgfZQ/h+iA99iHzon1MaACBwJP3LuqQkUiV6iBkXXq8MjEUjuiXR
MCsmQMbrEtj47bvH6DVwwqpjpotJP7+EJODPY3gonCl8/JyYUiXoOKVbSTFE
qg4Q16U3LrXWrD/ZQVHn+AUEsOYTMcIj+hCxE8gu9O2auQTvRULmelpXE6VW
gSxAXfKgnPWxkoQDolaD/WQFzoU0Y9ijUakm6+rEvCAC37L+cNUlWxQxGiSN
RlWIILHdaGp3y0QMxF8mFVYCvl72Kbc4q1Ho4EDX1/3r6eB59QjdBXdzLN+X
NJbf7ablhOHfNhA1Bgq8pO2F93+hKgm0KjjZWnLEVPs+g/fd6KP4IqfJWA/O
ORltx9b62Lh1MFdrO+KaXlEP6Wh1JOiF6x6BMBRDtlesh4h4Rf8OFiyXkIiB
SJZZCroC8ntRBkKRX0anOW/cxTtam3BsNWovpgLcE8Q1K/k8nu2986mGnyWu
BbkZ7Aw5VTEsv9UvVs4mCmBqXovFmZWlD/X7n9is2wewY9df+uGSMrxJ/W2c
yFYh3ci8FGnQOwa1AS3lUCNWJ1Yrsx09kA8/5qrre1aSRvlHBc82DcZqbx86
T9RTV9Xi+bnNeFA7y8WzvQxutAOvJczIFKUTrMKBbqpV9A5RW/NTJd9mV7sg
27N9o58UN97NbDZOmvZANrVb+MjuthITzU6aCZyYYe/kxSm8Z9/zVr5d/6xg
EzRPt2zwhb/Lifz9mJUa1MiDDXe1ReCFC6C1ZVAnAlO2+Nkwg3fWLQo8wQBk
YQL8EZlyfQLXX6D7QndPavr+eqIaiBxC3dYw+GCheoKZxzADYzo8v3zrwkBN
59b0TdGe1yTypoz5QQAncuF91b1/WOWjZcuhFGk3WXuXuhojFxpi13igd2ov
wL1JKIUstu0S42Y5DHIXT0j65bW7MfSBcLCF/TnWP/Wy0RZtBYDzJCVmHDtK
oowr2JdXyGyVbnsbH1Rgk7R1SqdV6qrAvKnrGk6KB102gW79gI+8nJVvMP01
oVYD+nLkp+QfE7zz5HSa0uqYrtXlrRopjyR1ISkU+NEIlJkNZ61lApC2kC4l
xwJN0dd9/s3A5Tl/j1EXbkKb/zJY2VhmfIedKngUGOppdGxeCTQHKvckpcUr
CM9Iu8zsKfzf4nXzfFjvi1wjhTEBZhW/abKT95UpiqPFpAaBUOkQ5djRWxZt
jEPge/O83j3c/A11pJeKJEChamFT6syibKVSfMKsPY2SwUrZbZPBhGSU+J09
PMOlxhZSncOEZijXz2ScKkkJgDMrO4X8v2gDlW5WICgYoDIaqMw3pZ1jWmXy
2e/9wwRpenINFYlu5joow/QFTsQzw6RqXAEEbwduhJ5+yiFge7Hybd0GmyoC
d9AR8esOe0BkxBKSsvSVdNTPLp3UuU/JZtQVOh1e8glK2X83YJWodhDQSAxU
8L/jWcIrKXizXw7TL3DsQCDcfXh9K3wPHTQiL5XVSLtRiLTCy5fJYXe5imUM
nN2MqUblllp8PI50HTgprXa067hrjAAGIwIe/Qo++PZTowNZg8TEJQsdAdq2
6VueRYKZDGfsrcM/qlnb4lLOShJHqtbWk+Tnjtpdf/UH+4XQRJcx0qp8kvOS
xyvgJ5d5f2aLhvNxE+L3GC7yeQA/wYGpSh9zNHEO33Gz9vP+uG6Peil8ONjm
djSkQiFJwbEwbpgDMzi1zMmi/UgyRuo2GIgM8Jle8xWm1UAXuzj3dE/ek5Aa
Hhmx0gI34e7UBNP2S1xzu5tghPGr/Llkq13lxIPUhkv4mGlRcVjssKRuwEZG
zK4dnKr2K12Lizuphaf8bUDULV51yYPNhWlIwo+pDS7EXw7ljSBcLtTXV56t
xrL6WW9P+XD59+f2eyfiRosXA9MIgMAZUTGsAl7ywtrTz3+08aq+njDnJzTT
lwLufZovbtgM3tPUMyVii4xlasnd0nlEtrlGvOyiKW2iADdO5xllRvKXPBSB
tX4jKzcBF8Km7t73x+jZS5EmetGXyotPHBf05OxkzZ/F1aCaoC3jRs6ArH25
nEzIgdQRQNYf29ezsb5kZGM7EtRmvtAeoxhqzSfTLTEkOF52Ui7OeOOjxP2m
l1SKQ+oU6nYyuB6w+kk6cOeadraqIuB1uPoBljVU9qfhyWQi0M9VJ9Do7kCf
L6FqXDreocEBUH/7K+n+/N6kjp+KsfCrD779AQkOp+KwWvU8/PZ77hSN31pr
YzvHDbWaoQVrvIbkqsowPlt7gDHPmir389pcEPZWjVI7B4sY7GNhhPfvGkRV
UoLiEFlqeuJanPc86T+ZHEBlKjnU/Tuu0itxnv67XDRRbKbYm2LoQ7jK39aF
KEQzMGdgF5Be0lAUbjM1+rxT6YobRUvfbndX5itNgm/rRww3JUukiFGNj+lK
5sc8GPks3AEzPxhuaTMwWK21Rr2lJi7bmXop9figZZc7E/j6lxgAstdinxaU
RUTTSu4qhW5qmrD32Xgd5vBadNkqNPLxPDqJvF38+mKD28i0scKr/qXR+hRu
R7w17fy/OaAcQsbchJClxuFbXxDGOizzP1HLnB3jTjvrjTnonMQuvQb/eYJF
1MkO/U9l7OKc5MGRQ3K+0O+P8PSN779z+tOkAlt5mHGA0rMLQzgVCibiqJmK
iURwApFudrdYyVLG35Gtv0dd5hp85hU1VLaandM8s2zpryEGKC+WHY2cl0wg
jQUHHPY+SuEsj8ZA3+aOsvBz5xfSxdsgcn8ltt9rPvJmkDe2DUJoihaHZlq2
7nW0g8b9JI1GO1F8i5dhvp8HIMvXiC3VZIonHP2XgwJ7U0OSko5eUyMtXG41
GyH9ctc9OC/B78tk5diwGctx+hvAdJjm3qZP4T2Pa/mU1sjPyHO1DoU7vNng
EacPQ9eRJ0PRkP5JkKuztVE2khIyW0oFozVJgBY6+kl21SLIGOtBOI1Br25P
7LUvv4hoNQzSChKYJy+fNPUUVueboFd2PCXEDZUex94TBnKGPjypJPLPWhwZ
12coH13qohH2TjFQZcxqB/qOiHHoMjawkQWEMRYSsi3fsyz2X/ushSS0827I
hSiV6vOuVLCsNoZsM49Iu7VE3UDBqv74m06lR68TRe0OmeaEsth9O+awfFZ+
dtFQ484RFNi81hdNRHScM6xfr2io5Al+EXWsLS/hfYxlZxdLHBdKCxanGXrR
V8ppvUNMrEVLl66EKlXCFruVqKoOMuJLfz29gvJoRhy8OuwL9fXeXCVBDInm
zT6oZ0tOr0KMJClThyzAv30b/i1eN0RxvVGa6zKYaP8C8CIa9+IY3tGNJFQ6
tSxpQSMPYkndR4fk+AicaQn6hlwZNwq520irqOkTyWAGtgElNDzxaR98+PId
HQkaTugl5MoUBMpyh1UoVnEODgz0Cwxd2OB+SxgDmJVAsjh8RuXHylGpn+4K
P3WMkAhDTgvZX8WUY/kO3KiowXgg++WxWl8ZGk3ekmfZexewI2bGpjGFY6fp
+6OIIfQHI1PZECfk8/6Fae3y8MU+swGJjM1dk+QmpuMhqRiBGcWr08DDbkJ5
lTOatBlwoP09vjDWgTAU3HF5jcAHL1b0mIzMhuu9Mt64eUYFDzDxlLQB+qkj
2BnDd8VX517OUMTN+kc7HTy6kodGGHBWBf1f1ifQktLYpmohOkr8JZdMnfnD
F5yBtIoB06GPYItSRTLBQWh7xGpL+z12WYUbLirRPxFazFj7JKAEpWL/U2Un
r1AaTcO21YLNwtY1FjcCSYJTIRy59TRgPJ1NQsbBjE1ngkDrECUiYmr4P6HI
Hi/9DJVXcNa47nIq4Xw7FzaminPWuyvlSeWO0rEG9sRhp4uZdF3LovU5HHgz
Gdwt8zFlMxMXFuf8/tz8gfm//j9O2EKS1WpSYp0Tka/bvdUjsQ8dpsI9EDuK
BDDRhkcCa5JyBvhn2sHhsmFaNC2Vycn3CK0dwtvkW3jMGvO5jvRj2urOqSD4
qjPMhkxIkwTaoUFzQbAmWJiYkR/a/5rbBRu81XSfi0wkq5Bh6yZrP0mSfzle
QM+z4my+HtPW0e3Drk1NT/tXHS8cmxlE614aOKYoCimj6HO7bPJ7c5BmCDjx
yz7O6yWCD5tjNMPtqFkmQeq7Trt0A9f4K02/d551I+AtKTGKjLFksbd+Qfxt
2N1Uovu7nQHmlK0/IiZoD9kHnp3f4kBbiXVwIYQTosDDlyteKZYqugAoaa6f
CmNuh3JKgyAtHL4Wc3qmLRkJwuhDlWlIB8zL01nQFM08G9i/oHx5Ucv8YDxg
I/xiSlevuA/kAlDa93fCqM7YiA17MJi83EkMaHvkyNGqkku4odBqRLLEcaTZ
2J3gMKIsEs7oN/aLC19fWeavXuACUVsKYSqCSraLo/Pt5p/V5i2u7fHnIA4Y
cJXkw6WUZ+JMC7+Bh/kjLio1taXnHxqM9gkE/1WoOJG8hcLI9482U7hJm17N
rrl00LyU8DR9dHuIhc/weXPsDDAJI556MwajZ5J9MLtdp+PKFnxfZAAKP5C6
hXfwM+2Hckcmq3oNzeb4HYaDaOb9MWpBY653AIwS2uEYW/jaWV0qu1kuyShN
cZ/24T/IpKBc2hbLjq559ezzOrci41ibwX6ri9tnucQ9eAog9L2ye4f+Vjap
1GWG2ZCI/lXEeDax9XbihgEMsyncK/lw9wA35axAkEDCw2ru0FkwhEtZFqn2
tqwT6EWNJNn/mhAqvftbehEFUaSe44ACa4jgRVKKAiaJrmLHfq+C2CgLX8U6
gkDpmexX+zJfVOB8tzfk7Rv9mraOhVt5RAX4J8xVc2mCOnka5q3Tfhn5hq8Y
8afdhd6LVd8EhPPPhJzJK75YFTTZ7RFwixRUn85eFZADil41wOlXiwUJXPLm
pNW9FRN5AKZEtgUboLQpoq0VhHPnPhi2Hx0LJarGvvkrg3mQHXby25EgYBgV
lWAqtIoZDN5g6rNDBnT8SPPC2WoM1tUnFy7t2Sjgd3ozQxRqiHPkUUCRkCRW
Hr5CM77l4yBnPxjN+CrMPqwqy3TbqB/SxKtJpXkgE5AQ0onhaBw5mQM0PxMH
nRtJR4ytXqKwz3VgPenKD8zVgXvwRtXEm0CkFYgbviut3JJpsdIQOJS3sE4S
2c0p98TopWyO8jPIiFNLfhrDdoGzeEuVOnET1j0Jlu86g6tes2p75uqlPs1V
Y75y9nB1/FC69bLdXKPN82LSWrCIpIcDCzIoNqfAL72uxB8/kA+Zhob80Zkp
IXqSVZvbJvGkrCHB15oVoMdfch/rQlXsR8JAkVBBrDfCdkHrMST9tAt8vb85
8TtTE0jU5GkuCadJw1OJKhtzwsi/qsw7H9yEDlp9qqPVsMcOKti7/5Qs1eOr
a+M6YTteSEunIv0EIqejHy7rN3qVlMrrerPfOx29gzSLpH8f5zOZywqO5n0S
2exfK36zhckxIr8ynr8Nz99fmivYgY/11z3WPtlCadnvUoqEmoXUIO9Lxxx5
WxZw7UcQQx4jN5j8WCbcdwd0dy/zzdiqvyTkhwggu7Tx1fU2V4sPbVfUYSBL
Jaabi0d+UzAedBhWvRlWqDLXg6CYN6cmtL5Fbr7l96Vwox7G5tbpx6iYZu/e
5UqHt/EabUSBhtAaPsd3I9GOBO6YvzbufnjGsX3e3UELn1O+OQc8BXY7Dh1T
0STeQwBLCVyg85IBKeKfqG297pyzpKvNBKD2LtoZ+rhpcSsPcrkXzTiC6VFw
zBncyGaDPjdvFrxqktF1cw2C19S6go+McDxcag9lBl0qCrO66Dino/HbwmSJ
0moycNr9Dj/JG/hGz/aI9VrHBx2KjzuJ40364F27WFs0HPZgnFsceewegqNF
+Yhn130hVB+ZL8c3ZqHeR1w3uYTT+OBrg2rraRFauVoXCMAVRKMU8Iz5Q57E
8K3Lr0vDM+Od7gMJHLWDLDQUmDc2j+hw410TXTqa7+rLtjB5BfYPWm7/5L2T
FoxCtIoc6KkuE3vSrifMGwgU5/cvvehfQWBCevIdVIrjAYDL2RMzcJ53T5if
h71FFwGiZwnjxIpgPQSjxhY7domFtIsydldnY42V1714RPxi0Xv+lSTWwj26
lEBNJs0sBs05DHSnnJ0SzoR8/CKHoYgLZGkqT3pkbESJUTGuv6E3bMLd1h5V
MGiECs5aZHNVj7at3nx1DTrB964n8OWGAtDkDzo0b+L9zkGSLX7QeOgBjuPm
VO0oBYxC6ZGxeVW0Pz3aPSZyY76PA55Eq1d8CFtXMbD2GkEowqO0+7zgXPJq
JhCvVHQw2KdmUtVJOxIaKPqoQWvE4SZTo5p50ydQhl/c+LY/uFM47DhMK2Bq
z5TqUxU4hWLBPkqOLu8GEjFIrLzDlh2DhtGUwu6V1ovyPnnOMMZ+nPsDw0CL
RnzSCY3T3j9JNS1i2NKG9IvpkB2g/IUV677hFBkjaKJfC8JdeiN3eQF4njkR
WaXpGKgGn3WSkgum6c0SF/embduDGh65UfIpz359p86i1pEJg+CAX5YO0V0n
m243LTUK4bq0DXLiMex9yXV6ddrJExEzowOuLYljGUEBtfGd8HWdjXiWLE8u
50o0Lz/3UlYy+WuQMxN79900BkkG0nEhHbgxm8jW3ullWGSXIvOBi4L5m0Mi
z9rYJyp/oCLQlmZVdXbA3oCaGPvjYMTKMofhf3rsXIKtYTEwdksSXJapgX80
OizXxt7Eo9Hute0kvwMe8zNy9uMWJ4lJdAiuQ82DWSvWbSZnjsBc0DbiS64z
JMz2mMXllU6H/lFweTd2aFkzIfGThepG8quoFtqeTVYxF1T6eL2EImYrhtBg
z9ZKYP7R++Y0y/9U9XAFYsXeBylOooG/ESZSO5Vfj68mHBhS0zRFjh93NYly
6Nz/InLuvQKjldyVNeA4A28o2ualF3K7jehN/R+SIzNoAL2Cf009Bz9+4WKz
ijJSnhYg0n+Ts5E1FN6CPfpK/x7//jThNC7M/zEGIbNJK63AkhfrCRLot6m8
Y33bE6g5CyHyYwPFFNi5uJClMB84T0niHYFHjkPVw1xrQINdyQZRz64kKMK0
f4aVmj8gOq5EStF8gijUwH07z/eyJWScFGXtzWfMkScjKX5Uww+pwJvsJOXV
sLVY3vigysmNdlv7BCxEaQ7hJo/0+v5EspAVcIzW/r6TOTnmfiAmpJIeLSTo
57rfcFnRNgW3UbBPzOPYEykOfLpKzavjtRq1vIYgNKtVYEweblG3k+IERJVe
0y9FTtA5Is9ULMFryyUud8x40JuGPviIEt10IaFBlEwcjK24SOuuInA8A2PW
U/JAAy3w3bMavDDZnUX+8p6k4y1LeDHzg1TxMwP7O8tEy7su50+T071KdUCP
BhNxSlAHbWYmJniIrXRlPfU+/Hl5hVnq0X/ucefdtgsfCwF7OvdfPflJ3qSI
1YJQyr07M388GqYjdlfvFngoYlgvENECGcq3vAgGDdpceniZfukC8uzzAxqG
ydALDDUI6gTRuNsw2yKagBkbcMasWYA3nsDcur1bwg7xfp++ova1s6bAvhbx
sF8NYYtCXc8Pk8mqQb7sAC03yixnrfwg+OaHfpqO9XEBM23Y36iEdXvVgflQ
j951yFCSKBBztVRvTAQFTafXzh7bIijz9o6grizzIBIX5T4V3lOiBnixlK/a
696yJwjykM8Uvu2MahE291oupd1M8hD6SDj06tz49IBxFQ+KMJEUzN+Czh2h
RCv8uqCPCOjP85+zd4WP6OBzjXDWGtv1O7Npq/d86yEpem+Mgi24MLe4JJb8
NGBhPqsUYjPYMwaLMJQUBsT4PSzxvpRqHgKgPHm81dUDEJz6hipzm5X5Diqj
CcVScIQBVtXIpNJxdXBqrTMBB6L5/OOjQDzYixM9gVHpJiHmGkzzc6kpwPQC
qQklviGGfXxbxYsc9/tn/56R4pSoY21VBHU323S8JBpHNyXHSYfMz5P+1q3Z
Ndx1hrcLpcvwqcdsXjRVy6okL6kjlQEazDkkalQ6IZWvSuogu+ACyk2OdPlJ
NA3f+plkdnpf/UICujrkm7MBw7GwT67aq09RJIm9ki/qAWOSfrq7hPo6ccWO
kUQTxdZ/XsfjlWGjudiWFYYUsU5LlR9Ab8Tm1//U4/e868lacG5o5izgGVkV
te4J4B+obU9DlVBIraKHiiTCYQP9uKEU/6M7LEL1JsSckrQ0OT1O90s75TjO
gAC9MPcuv1ox+SytF8YXOFAsLaC8Fu86WQC88wNHYFdnr9n92jZVYj1TL6uY
o7f+6Vs84j5C4DibuRTzzj9ukLnxPiwqEojcKtTtPTAudG2MyJ7UnzuucxRA
mvxka9Jg+ezrJasqiO62Xtf9iM7EwVDCGDRVmmQrWUtfxMuzmKC2f6J8sPuY
E8Xj/YA4C7haeuu/X1sakCXOAB+eiRyCEYWuFya+soZixdcQUfOGqnqy+9eC
8yUZBmhASd2NZ4kQe+jHGcDhdlCytyIGNx678/lMjGLxV2XRMkt+uNdzaX0b
ijwROgx62hoNjMJxLjSiDHpe7Opizfv+2wA3n12bxo6UI4LMazSPHCdRwcBx
Ux5Sr4NzWgnGzeudAJ8taM/68fRQ/kIKEaLYMroJv+fYkA6doJ08KN+3jw0T
jaHb0j2Rc6sxd0kmJ7YGnoI1Lqx64GbQ2BI8rOdzb5+ijg8IK+4bLOgJIL4V
oa8tqS54K3NRaNJmOb597NjOgk/hZ9L3J14Dsiahb1w+gxw0zQLXCM4VU4IR
wcN+zjHbeq6gPaX3Ve11KMCwzXAMX3DA+Z2u1gXtreNE//CgrFemLohXcJJM
vpJ1UEcNYalTCFCheXEs3jiwuX69wo30u0QbQRZssQhuEm79Xe9yvUurV9G0
2tplq4dANkWrSTDVWSkYWbCOAt3ES98Ge5Q7eqmA+QBcq+PnbOaZQJrKxqJF
PcWLU2cAW9+SAoHfZneI5xqs9qsVZMyVmGkzL97jZsUnNIgT0O1isJBVlPEw
FaaNrTnP7cC4Epvp9KYSiU8iEyvwswRXJ/pCFY9sk1VBAjy+Ojb/EkJXuuh4
rG1Xf8QjC4H33fodP/PPRVa+/zhUzo0Rqe8iMxqfIeFfUtokWvqdE6Lw+mcH
APsiA5e3PL+g6kZlKI7Hyyr+O/zmUb5s23Q6w/49IWV5rJSdk09kHSd1yuwC
1e95HUzBdQ3p9LL/LcQw08mSahG9a+ZLWpkSrc7npEkzTpLHw71gPSjIHOXv
z9KQilKVF8RYp0vrqbyzRRwJ7fWfFsxVsblCg6bJGAT2eni55VES+Y0dX+Wr
7v4b1dMa1snFdk3TLeHnusmNCq/rbDzRFl0qajCMLJZAxnk807sJ3H4osDTg
LG3d1IvKEkxmX/CZj7fRho4LMDJTY+oN4wYxzFG5qIN797vfG3T6sn7xmnzG
n/dagQIV//5qdhNS/qP471IqRkxkXPpagcNrtEVdqxGF+BiqaVTTAyk1jAdc
zXsf4ysD3MU32TLW5F+EWO6zLMq6UyYilST/szWOx1oSPNNq6C+G0hNg/NuT
TMGnOXguopqlkrKxZ7oxgeM/KoXlLrSzzxqCZGfd1OzsJt1IuYvr/IWz5mYX
Ya2Bw3rE29w0tdEo68tpOFRumO1XbGAs6GXNqfXYoD1pDzY146PTqzMmghQw
nCqICSKm1RouShwxBJQK2lJ/nKFcxNW60sef8OWbr9UfL9ay0+LgPMTX9EqV
eEKVA2Tfzr7fF7y9kz+67A6IADivy88u+l3wgbbCkVOvi6oytO5Az8j5UB44
wX7z9/wJdp3IZprmThg9TT1qi8gGRGNL04I8Ru3FYU9j8Fg7SjIr/YeZrJ/r
ed8eoq+vP2YSdqdYoZS5ByB8DMeTLnKLQg/j/ON1f/b0tlJprRYefl0vkZ9c
1VsFQ6ioCbvcZWH+7pBH0BPPgTQqBputcn4saCsqra/i+PxiAiTJoid0PBDK
lednYKIKy1gEb1tJyyJ1hgQZalTCJaMS64eXoyAisbPZ6BXU9nHh8zA82Zkf
BPpBMWPms0p9fRXSrgdIzZ4TsxuwAyNCT2aP/jUlhvv8joq8i9h1N2gs8R/O
i+KiRxXTpdJbNE2cWTZoBnau+IMlGXKFqrlB8msZtTCfLt6O+vLQcwH5Q8Ns
oCqMNN9UzlHjmyhq5Gnji/dMaQLCi1ot+wkeY4NrGsPRaf8wk85yrhme4+na
X8EgJPlC0MiIjze60F5O/JTEGBOsda9uyyuNvWKeVI7XhkAlPp7V4yzIJPOX
9ybF6nJoE2JMyLOPsFuhOkwMTCHZf31TKzx3YYCtTSJcVIFcOKvzn5jOFC/k
ZRF8tg+rdC4oTG5gUKfvoYJU0M5yV1ifzlnoZNa3wDyxtIJzAPPUMig/C3OV
D7v5+fik/zvc/oRLBZa145siuekJYz968Eh8x8x0Pl02NrfmxqvgYkpgfEiQ
ONEMWZyUJ+tN/8kQu57+YCOnzXSeapjCGWg1ah4V2krTEobjbGSl9EAh70Ed
LC5PbRkdl+VTxp4bswS2onIrpDhk248OvSzPLfNxpUe545UBcuk++atmv9aK
v95Vrsl7FtcDovCPVA9mjG3+DSFwRWeAm9Sqtq38I8hb3YOFVvaCXo+vcYu6
bGafR6we6Klc7HL9dwC1IS6lfHv1vBs6MCa3cAP9RsNSyA+5HMdpzb9crARG
5oQxiAMs/XEZI9KNf2iiVc0aYYZ4KB3YBKEL56XhUWPiid5ABZxnOUpedvVO
UBwKJe4V4lQMt3juF9qrFMKpwyqqCvHGoYViaxL9fDnamqyZqLhQVrtdNdc0
bi+WWKnrsmdEDJx3mg2Xy0zf/hnHuX9LfNxfFCLSR4RKW+4DNFAyMgkoNdVz
FiK6bbGi/sE0URCvLFL6teQOK6v31ClWcehK1F4IOXa1m0iQ2oqsuGnICS1X
REcC+W+qlumPvM29vb4AT8EJRbe77ezcXaoakfpYU9TaD5fKM+iis5gYdcWN
IP0dojr/O3sPpzoCZZU+tA7s9nqukynQPl+Frvz75YQV2KTHQPKZcBGhPcx/
IMPDvqxM+E9pgGE+eM/Lt3ufw/WSuTKo45THi4dUDvTWjiPQ2rpq4a9V2Ndj
tuwW0JRGz1fAWuEeQLIZHxszpaB8bf9RYyC0NA1IRnHKtCinzwUW4+X0lnSU
DeICrxSum3sAtEoL4s8YDO/DIF5ra8iacABjy38iKYdm4zAmoW0Ng+28ZhgZ
W+NeE6ZgrfC9NaV9Z9N27/MXmu4GQROJcX69j4BL3tM5BmQuIZQgGWoirzzI
ykllhr1/Q16wWBNen8RvjDS+sCdE9q78fbHV0VNONYDzdLggcmQZhXXZM95W
adleLtf++KCnMJ4CPEVYhjQZ7rDCV64FKAJOCkDKY8W4Q91EILR8Lhnq1Dbt
eaEVyphBad9MF+oOTkYh9srr6ZS/izJj7P/OKrz7u4Z1u7CvG/uCUpdfFg3l
9w7zkm2oTuEF5YMD72Nc1zpDx8rp6kDtSsvRqab5xEYh31Ymk7fo7KVDgRNc
edYRex7Wgh2lehQyxSYlYKAc2m/xwE9H8h6lDd3h7M0aCTcDqfzc8vANcBZr
+/b3wrNCYpBjX0OWgASrIK4oyRODEK1aa7WNGcegrGUShc9ad346JXbFlqSh
/ir7uU4OWTfn+GH3HBA8A/ECnvrmAnVVK0WVa1yx4Od65yDmSfutynU8FqqC
pkHCtdAZ5x+xvEzNt57cVlFiKZ3KBiNo87aqV59H0QooxoIqoZhOHKxgzB+z
0Q+a+Yyaxmd8PQToMYRfTPxF0QCQgfZa5rhqHAOdQ9bcAEh+Jv3SnZ+JWdw5
545o6t9n2SjGzdUTknz5cPAuEw5uZJnTMMyrAKPaubC1MVPHPO7vHA/k3gLt
OcNnqf0GNPv/BHDqZ9k8dzAyXDfAnLCJTSdobtQUATimb1q96Tg5OMibFud0
8f1eTciLKLGU4rbqC3Z4K4Xhg9VTJbdBPDjvgrT+0zMXM0HHKqeXJazH6Fa/
0Q1U06CrcJUqD4kekk5NoeRPG9g6O7Cm7cU8Mke+ApNP+e4N30kj2Fu6n1gz
jR0j8j63NzmL1eimqgH/CPSlD7e+pj0zS0bsLS8HRDEmPXIWM9H6E0h8VqWt
p4KZM24+cfDNh9/g4Q/hzu8S2Cg8hMfmOs5sAkfb4MaIVM1keUl2z3DM70Ln
GsHzLnp3T6zZHRT7GjwFj2Y97iIUz/XZhzhfV2Gh1aHhMKE4WxCLvceh7DQ5
BZxWvMiNMsPDtP3opa5ldVnQ2Cbs+cKPOs2HfJSveP1fa8+FAKrLkgsR5mz/
AIPwqFcNf0dKMxNoTn/RG2spL1vmQ8wBhc19RNWjW6ebGb+YPD+x7sQVPkHE
pCs16fThuAQGFCREuQOU/gjNf6+p7r8IPwp9UfVwp3NvUylwkql4An78MSPO
d6eVQahpWp8os3JrVqgiHNWgcl7TCJWcgwTHaKxwkIZiDbC6sfc465BqJP/n
aS74jIRsgfCVGV83/Xl0/LrvOtQKR3VEQA2xNGlFkkvERJ/OIeq/IDQKmq1f
cpWBjX24EuHXaeV/bK92ljBXTr/xJ9SIw2PIbAXe55yqiHZ/hG3i14znIEgi
nvjaudkT7HF4N0ltlMuKYL2A+1pEWvGPk9ixsMIFYGHRzsNkRAl7iSyW4+6F
jtubl8DlDHv4F9SQqSgWo4OAiNCrINRcPqbPQ2t1Mc+BPlClfFLAdBqiDPDl
wLU9IK1X8s0qbFmsq9oQcZbBrVTrXkiqckwcismStxALLtxCvpxXQxSjtuGO
FI0qlgMdB21KO6wCmA2TSmjozkTTYmreMU7XaK1auJBoFhpnRTPRzWQevlJZ
RcOlj4WD9AARb8QtMI2/KSl07i+dG46RrdtxwDHKTx/yfyCyZnbPf06pJ2ix
5UYXzdjB6f4k0AH2b081dOowbxon8bg4m4le5oB+hcdxzGG5aiV6MiyLbdiH
Vih8AHcJ7dPMKLXITRimCN5kEH64T9mCS0BHLwtsP33NAfSbRcu6uf0lDUTC
f5UwUVs7ncrzlQmzsuePUghk6ruxyoPY0rkXCG/S1KIDDXl5LJ3uz22Zly+C
nqGWNku+KslIIXRe+gm1A3fRs32IuOwwlku/26wt7fWccWS1ezyRn5FM+dil
9CIPf7cIlKHKAGIDB+SHzvjBlGXZYt5pfdfvoS+UlJgTxh5vXGTiD5GfFDDY
w5SfpKhnaUIhZrhuJ0CuX36Cpf5Q0fiR+OE32rrHdtwnHvIa4rlzqFoltOpw
N6qI1CGL1E1p0ww+brFK1b0s146umKZRMHRwvBJxiJgImunGCtFPr7bD8Nmv
PNMv/+RJ0iypKCa3I7HOMWc5OTgqedl83OHJQ4qesb63enyv4UdMZ8DL/azY
dyaX3xDceXSUfRJ2lbiKbut4NGErQcoxDh3IBxY7/U6C54H++kGQkfvO1pZY
Zb+Z08x8uCr8GgNPnto2/V2VkzTUbNTfXoFd11qB6vn3YiQZ0/2L5nHuN0Tx
23Sh0hj6bomIFgAkX+bZICWRJp6n0PzRB2dPBm19rLoXWj+2k/TFh/hW4SkH
D62MqKfwR37TG0cn9mHZ3bxWXjq0asesCft+Sji/bO7ummOrmbi0NThOAZ0h
+D0Kosiwvj55iCwvk2wS1GZFzrlS7wUSMn8UxIooLw7vAkt3LVXcaUEYYeOv
7D80ZZgubAkDRvTPQmXx+L89L9qqBy8JeNfWhy+CM+RQD4DibK6aw+jXODzm
TxhdhmvmFDaCjboFt2mOUdD9aKwLRYKPCgnODQ+NC6StPsPgDmsdtv4tmODs
rh/mEtVZCgV0uv4lj/DqeaAzZCUmvVE1J6OYboVlEOce/o7Q37bqBZ/s+3+T
PuQzVXRlX0TpDJwim8/WcaZzRgW+SGjAZrL9WLF/DZRt5B+urdoI375ck+Qg
5PYfbgpQoL9hhXxx8rxBtDgnYfZ/7KrHJDNYhseIWGnac4LzPATaDtNLxl2o
Gx5GfEE01h15ZDDd3RUhOLXsWVkg+DQEwUH0L6G2Luwe7Yo3uP0/l07bRJGQ
O9qZWW6zqjSbb3RzPSo67364f8IWHrHFAyo1cGldiBKp2kHV4dfbDAPsYPt5
YE+Px2YFDOoy+PKqzLLae0pl32jdNMu3oR1oe4u80Vdr/wqbfCsqb/p2ev/w
jBb610MIL5xRAKgC77qnLec2bxjKiJIaOXa3AMt0zo1lZM6RfEIn9QGJrbqD
pw1JzuwWuOh81KRu4MhN+eaOxR8wXCwuuD6JvZwICbxG6NOGcKPiV17JXWp5
Q5oA60Q9Yr0n13JoqRRtclmWQb/ecQrluTLr3D31d9mfi/f7HQtQU1dMhjNi
CQ5PYk2M+U/dVsE/yvAoJWfk84n6rk/6dZb67xgoiv+OTFVjBs3c5N0HZBye
JDs+rLDHNIq5WhBpE4Q3DIwGAGXimoOin9BFIXAdeCED07coV6j108d+lTnm
Od8Qacq7gTQQ67OeM6azvvOMAPCVxy+tL+0ByMsEt9lUhE8CVI8Wfy+ketuT
MwWseSNgDSXNdTMsGqAPltMEThKnxqThxfNNCAoY1MaUADFlvKgv/bTvOfc6
KcNUge221SZCdNdQ/qCt0sorxey0Hnxr+rcXvhK10Te6/aECjzv32DcbfLjW
LLmMi42PvRivqMxhFx7Rj2WGVQaXmvsci07+dj0wv1KmFImiInUUcswi3VMT
ljk4qs5skQoqafTew3qCR9yP20U6SJHVUNTPBOpGNF86ih6/E9dC10xXBOPV
gv7Hm7BIErZ+YyBFSzXyq2mvNQJwzoLYdY8MuP2LKGr1W2gnVRrD5LNEUuim
S+rSBz5x6IWvCI3RuVTbEa34gkNPHu+b25eFj4ptrV3JMsUY0dYYdJFuh+8R
kmTOIZZnU4TFygLf1SDh70WAi6ZYQM+aXE3n3rWEz529F7o47iRhVZhfgqrk
j5y/PMJ/MNYIYH72SRIVlOEZnrAl/YVNsTby65iDg7ithA/ilACF4dUA37vR
P0Ah5InBQ2uRyEnCvyGCz7TDN+PxbGD7iY3MrNFqcy13uu4WgnpXHhP4guBv
fHW4bh00XK6cDjva5X5zcXbzlDP96l8eBd4fuBtzOxr511ae5p3k6+ezwKwD
D9MYZM222hz5+fhoOUcI3q4bCLnt4M92KLAt51xLeJeqzJH2WWY976dXq9ID
rrBxxYFsKN+418WCx6G4OOYaZAy3DEPyquiMijgJMOAfjH01PSmfN2GCyXg5
Zj00o+Z5TH/ipQzduXO2yyfIUoglGfUFPb7F76/9TmdWI//+DseJF3NBsVvS
uu20wZ9Koi/XZMOtAvRqxE/AxXBwGRvUDol2/5GYuXmyX16Wgih0D/4Uuxbl
tfPuEZXJxFDjPiZzfEOHrnVUy6rA86UhnZ7b9wol1+lAz/jOZQZ52F2dAYbY
VEju+fcGdf5ZPrukoEvXWk7RVuKhEvVJuaqTpKayFPL8RvFnkNnNj6QqIExB
yH3XbHvOOtcQqUJVulRJyd/FqL91NZRiQoyzGokMf/kz+zVkFrlA6G3tiN8Y
5kXY6Kl5Kt65sNoDwlKLVsbArurY0+g8SvIe9ie6ZcDFbXBpk3QvCBHsq8l5
1Jm3sfrOvbUU1OaASOd0xQQDNaIlbmnLGgfFXCmbsvFNJ5pjv5IYTFMaYUX/
PJ2DtPR2m9IQUb+hm0BXm29qTfwCQsA6AVtxtEoThxbncT09TI8nMKTwVAFR
w+mtxZPPtb5PdL95baMDDZjT5Ou6RmLAL2tbj1I/GRitzgrl20nc/XEj8StK
vGNx9h6Dh/pG/yZie/Qlutc8Ij/VIsIohan7/bAt++y/QefZLvT6UTWlVA8+
okQetgCGdO1zhW1MpIrxTZuZTXQ7QmnaiOWWLvuGRJOEiMkRA/L5JG7dHfbP
UDmgfyORbA5S3GjpS8h1u1KKlmO1jAyurLk+GoisF4UDQ517RNueIIK7RSxa
BFumTJxWyxzUuBVQIRT6pw+MUJ3k2X7Iu7qsG3r5XFJj6Rir8iGM2atGVVeO
CDiGtNrTRx3nUOCxxRskV0BGOAp16ERD0ZpsxqdhQps41XkooBuOaxEYP+jn
ZdwgC0HNOoK0KasrDgdFjZOypv071sOohaRJXRvR6fBrCaZpFa+FL+EbE84s
E89VGteYaC9FoazeUxMTSHzvubSd8sNSWFR45khZBNVAbk1wEE0S29zkvWhT
FXke6UNcdUi916/unaONokUlX7XYqPTogR81aZTVRy30cE6XeLKvBpNd16TR
UbmnK4I345eiCa4uXZFxwPlfwSsXo+fZ7TtpNyWOhsZMeDF2m+C5AAwxJ5mF
RiQwkfhOzNAPbq/Pt+OPSxo7x6uzzeRM++ybB3eHPo42Y7UoxKBe6C9c+JeE
n331BdyI18kc/1o3MMdVDwOFPKw6k341wy6DDbFsykl819zQoj580+97Pvpn
ObBPkbLE41eSc+739GPCJXL6QJEamO9bUELITEYs4XiIL7k+TxxXV51zaAIx
fBEcvbXyHorgoBsT/rrLGkRwZ9y9fb7Vlx73SCJZmiByx066ItZ0A15k2yAL
XEZLWCKicYKzAQl/5cSvadX585p5KvvFlK+X50OIKFahtSrqZXS6FgkS2ee/
evmhHf1zWZsLRtShnsb/bDCavAqCJ3lg97MweCwq29RoB7fKOWtOKQQhq+Iy
VW1MqqfmZ26j7kXbq6aauV8Wk9PvSq4nIt7E3e8b3lA+VijMELZ6YXzXletE
8b/m0r4WTSQ9IT5GdMbUBPu8zCaqsOLtPv7DEQKuS6yAUMMsCRqw2Aj4BpfA
o9492YJ+KXIAEuD21qYFgLcwCkGQHZWw17SrmhRgHh26u3hC4aIsNoculfic
AK0yM3HEzHaeolxiPI96PrhKRLNgb0k9hwdpaDoaiO4OB7rol/tIMZY73hf1
3Nm9ALD1IseR6HNUXHL6nNZUebOmBxZeaULs2PGwvGrznPOayOvehn6vZm6M
Ga6MLK9gyJQXWd810uONoINLHTX5/KczxFDRluZO+6UNkJP2QkB2Ksnnsm6D
T3mQoKRhcp3kncDenSb/wWgwtoiBjrF0S7yVc9nWbPaCqKJbwYwybW5FVqq5
2JMytV1w7YXbSQ1M/LiIE38sZyuJEv7PYENwHa15TUy7kKVjEj8qNZGfZ7pr
KmoFIdhGFSyPBS5YTE/qC0Pz5MSwWJ19zvOjBYLsz7Yefvp5GeT+ZgRffl9R
Tjyh3XMGIyu39yC0ASt9HZtUaOR0bTNWvM1WnfFvUoIzAIYa475cxxRNNLdd
l5eZtFA0OlkNxahDMvo1rXxUUVKh/SlqqugcAsVzUNttmzjKKyce1MUWQ4cS
DA7x20pO0Ff1OPZx3VHObxuYgNB81U5JSQxgrLrnfDZJHaEyyChuu/wwm3bu
iXDTs08RHLQT4aodJYBOnMgsJd2fx+YtHFqV189AiPDjG0/rBbenhjwQDRLR
DGlh72WbtsOK93mHt37XWvP7ufJadJc1+lmzsyL9+3xgFi2vQVsyYk720Twv
3UkIIhNDe/hf52vNTdK5SpmJQ7jKJO0gOxJdxHdo7PAwq/c96BHjh8As1QkC
FF/Uq0K8NJWw8IRdBbSvxReelHAc157YY9yk2PMbsDVknUsdnKpIpFDmC9MH
CYQQHpnNLX0l2MgoSjEZp1qy8XAFJZaC/ymgWDGimc+9lkHpslWooAmeAlaR
e3PPqD/h1TLsv2xfk1udIf60KOlfFkwlJRTS8FDBE7nELSZrrfcB4vaflQUV
nxq3iuoWxc53BrRoXfK4nosN2e5lVFPDKgOfJLwfzpmZ6hl7caJEUdrlyub2
aj+PFqvuigCGlc3LlKZb/5bOV5xOD6DVYt1um7Z7/CZVbSdpw0nojfjN0Y+8
7oa4kQzpt15vlEJN5V2n8smdqk55WuUaB20oRJ14dFScH1bsIOmoOe7udmlj
nkgclLboWqBffJ6jlavgK0IylxTk2i76XsY4Xx9sdHSXRtnxU/EEad1tLuvV
Ik3JlaLrKoDB1Z3k7OUd1XzjyMPhGe7Yxgh8g0ILqH9GXD7bVcrJJx2AbeJG
BSh4+j6+4AU40iPYCaXOWJ1CpVofUHZQHa8/Y61DZZyJtXlHULqeUTXOlMav
cWTH7NOjKGS6JWgi+AYF7dcbMj+7s0fWPzzlY+AVFQdxoB5p90RxYFHFxk+T
esbvTPosSeK8y55+x4oUj8Q77c7PRz4E8J6iIxuDS1kYwn38uSTk97BYswF9
U/HpsNePAzorss7MIEsGZjgbd60L4++5lV6nXLZxKk1rJUbd9qtxagnP6Jy/
yUD4Ze3TQN2X2MK/TJDRiD23smVsAI6+Gqyf5zkFaHx38nNY5++X9bUnxRnd
XHI6XKWNgNLxzgwivu3Ei6IDl15b6vxNzTw3CrFpaWAoGjoz0LnMap1ojeAl
JQkRt5z/Qd64Bnk46Gl/lY1dS6iKQu95gtPB4qwkGAzVMClxOMkWOe9Yr7Rj
dAlgRKmLQ0DE1VAP73hNUBWCNw4ZXxhPJ5Dd0dJHELoPjZj6v3qQjfNNU8Sg
CKAjRrG234i5Ko4Tur0NJHUyLICuTF2PPqfAjOv6h+Lt+nwvUhS7uY9oirfB
c5XjqdYnuoLVGHQRRJ/zOkN7EgNRlvd5n7S20JriGNNXuGdMmDiMEmn2bNOA
GD9Vtu8G5AtK58uXBYH1ioDeD+mrztgPadTpxnN7jAGeX8taomE/NYPLHV5y
y4uq+BrAMSpkt/yQCtwSG46sKTZMnXICYs8QrtNpIkn9hh0yS5Q3EKscb3uq
f7B5tyyYUI3SZ+XWy6JLwPnzcLgRL4HB9ywLOmJEr4HSiZpFtJNQVUQwoqsY
MonwGb497PGPkxm4dYI7NAlmXbqjW1j8DTUz787lRNiMIiuSfM6QDYYOQBoo
id1mE39+zpqCoNcuPz0Lk5laLSdI30hyZDT21sooQwEwngChWSvXUg2iZk2M
LO+mpx2hJw+QS5LqG1pcdLwgJXxSAPFaHdm8/BqX6q/dfxbnb3wMEX1AlvZ3
SISVmr9s1HY/kWCauaHMvQ+hSXUH5U9twvQI3qZaUdRiR4EozaRSsDd5jga1
sPWsv3sOp2NLr+LGKsPQbPO4y6xSys4/b4cTHACJ7Ii4VetNQR1LP130Xcgv
4gmwUYqJDrz/eSIQmvIbItpH3hCB/fcbu4xzi4ibR2qSAFCjINctI7k/arEF
p0rbJGzc5sIBpXptQ8/xW0AatctxRqmHxU7aLNOBEaT8ppJZrz/WdAb0Xi9N
pEx9M1ZDFWWJ1pEbA+2wvdfBf2vmwkdw+KwS0TmcW4E1fUR755muu1Bbo5ej
Cvh+2YbrVSYewfvy78mAyAcwaqweawORT2nxrLzZmReNc0aEqVeyLUbZu7eo
PtloDtWSPzkBO9PY/6i+oOUw2UIoeZjtSfQHn4rUq81pk1iTmvcz8Z67mfDb
QuynVeMB77ZHy8BWBL4dYQcBAMwmK174Bm32piVzA/sN13yaQ6PzCL9+KCW/
Kda/uNQsbwHoZfRegHUyFBZxSc3Yljh4ojQu9dVSEGuS68rhq2jLboPqzSUB
YmoLU6EJfLSyZBdMYouIhD2wH/H+Vb4m8HD757ZVZZJTiHr2ejuc/qWe3sqY
K/NL398Qxk1kdGgmrWw5amE8fV7oYg/qJSaS9TeT7wk+rXhwAwgXS7uOXK7o
yON5vzocJiQWAtVZARpuFaoim2tyKjT9DxistcpBVJAQGz33WzSfB8JT9aAE
Td/kaSvhanpOeAiz8JuUTjAX71aN5VWCcA0UV1gxxdyHcMcdRrQtxq+0Tc7L
bDVHoCYXmGmA0K+12ANTxfW4px3mR59VuMRoI9nWqZd9HfzJkCYkwt0aYXkt
bHPKNAifPvvlchQOW/VcHINw07clQxMNL9v9akleMbgIO7pYA/u5NxFe8NEb
9JjpzrzUplQJNDNnieI08OHDhaaELDb692RfvY5/byKFOkI79dxZf1ZRd76D
LU9vQ9/Vabgtb9DCFQBy5woASXPfYEK/rqOmVr8exJFZsTzspRmH0qhX1gSa
Ylnft2ZCKMcGXzKnbfBuNqgjzCNYprJcpyfV2TiWEcn04ylYM80vBqxcHJPC
4YYqP2wlHckH2ZurVmCaii8ISC8mcXW21MJocrhJSpTnTgn+R3uQSjS+Zdk9
OaLZjSTLaOyN4UTT/h2WKY131mZvuLYLJVMiK6QjBZwTPN/Ulf+nov5jyjIg
o9SExB/T3NRT9TardtEvwnLDqykO6gExRSqDvlSrFJJ/Ec9dIOBtbnYqpfkQ
xlVbQWwXSE6gP6M8oXiwQc8UZFZlCwqjfosyDxQm0azMgS8W2TYZM0rHG0PF
2PCeDXbq8vee4hfGiufQ0jJ+1sQaQVqxqlfXv4VllSkrKjB+LifbpnQ7fQWe
9fFh5mPzUcYPgiVPBb6JedWqr+humIKQVh1yHu6C1utMXKht5j8+KeHTXAgk
wOKGowNxsC21rTJh6tzUJaN74llf+A81wIoIiJXvaUPvEW9EdA7ifTREEqg+
+IwVUgZELN3+qknY1xNrhTm1SibtMbDGPXTkHgX2yLe5qLKFgv5q4zRF5tvy
/IbP16PWNM5fX1wlWzwFYmhgUdl26slJO3OKeyUZ4JNc1R9SO6tWSNAAzZKw
fL8iDrihcsBuFVO2YCS5M1N6Kel2FRDdt6qD+VcYZmttaH1Eu8N2E8D+MdAU
aAHV4MeClXjO32clWQUJo9FKaLSmWOAfeyPE7zElrHyF7RY6LCQzpGeBgco3
H5JiBv9++i+0cpfRvy3ZKlVZ0+BDMOSyb3c2s0uMPe8Q98MJm4eZphOL+/Hn
huuVebwEIEjS5qUzLPCzZP+f+Hm+8JXpXJvoAi2C24LmBjhDD9X00tlVgI74
tZjQuDY3t7CX1t2Yn1Xoj7KBOc+S3VP+8BUtXBLQV46/N6VHuTC3O5zOaF6H
FTOYo8rNPxnrkba7N1bT8qc6FjPNf8s967pL7dlsDO9+J8uv9lsHSja1TAua
qsPjy6KTW8B4Hf3R3yJ3JkpwWxsDOVS4822M1B8JUwpSZH/kZz5PF087MxWD
wcfXHat/qbPdyPtGOcwBvxvYE8zTtiWTPZwUcG/D5ZOWUei2AaVu0PAB+dtT
yUlRpeWqTR58oVBs/PXW9OosPlVmsnubIbHMNUNttP3OoDDT+l09KbewGt7U
WRE72oa3dHSyq6QQCeEdwC0UAOyE//yR49nd9jYOvSOwfhs+MoqQvWYMGvpd
nMzlVn80mSbEypzjFcXI+sCTQQ/nCg0MIRKXcrP9RAI9K9RZzeX+J/oJ5HS+
V11U3sUoRNpkJ21ZL75b5y4uzUs5HCMDLXmPNLFFe7sZlUWrRAUPeZQb1z9D
ufFGPQZTTUDlm/qZ75mH094CHAN38PSiFR32EdZjvTc4ezpOly5HMV4NmlrB
gafLPTwHvzu2UCKXNTZeBLfMIDokeCEI5yPg6TBA5nbP+HuQ3m3CJVfKGCIi
suuT/CshJ8Ax/qQZ8mZ3hvk+96DMKxmd8ivChsU0XKhBF8wY/sLEllp70Z17
QI6ThuO8QBuaZhM640jiXEanco5QH3AH0MU4F3mptfyi/ek2v2mpD+1KDgbQ
tpyq4gzZwxZhKoXviA0V9NP1AEZR0Hmdjv1oLfobRzxWyCv/GGvzezrO5vlG
aEn/w/rS/kbwmTmTcsgOh891paPCF2Sy2//bNztfigUj+99vftkCYBOf91/U
pvT6IhHePLGaLf2y28uXK8Iy9L/szUuP+NZxjhD21JJ2pBemI6jqjUDkCIBk
nscoDjeySh1WIPzki30eeNr4r9lBiq8UY3woChZBX8UGWgbCb7Z/WX0cmtNH
o852I/TwXCsDSebAIt8dewJNGqkaLFzu+gYwQhGMbRzdXxOfHpi/vPX4TnzF
T+jhkclVGMRUsDiupJZAk9aycNUvQAc9/ckAM/g+6Jn9SQWi1zHojXwl7spo
teq+FlH1um/7rT7I40PbYHj1ZseyxgVmwHEt3igAFbV48eeNENyECEgRkGCA
WkQAy7EeyvJWPDetYxAEQJx7EODtR0xusTi0V5ThHiJ12UVwmbfT+mzTJSIc
ovW6hSetydKWCZkBarydEvlvR+70nlI93+z4kzWb7rda1qVx5g/P4whiFwfK
lRv2M78pu6SbE9osjNgmM1ulrRO0o7V9cvWWQ/l/cU+sJE8ZVo2gMz7cE08w
8JaSuru9yrgmoiaAD9kr7T/V6ZhFZIPxWi4ZwkNRQNXZav1JoJRfi6auhyUf
Po0cznCRm4JicJcIXquV+Tdvvl2meA4DxoV1AGN5lRi44Aj3n0P2mdbNhhoi
ukeIA+6Af5OcInxDdcRUI6yE2kMVCds4qTi4avNBwhnzW+XHfyRXPv9XBCv/
66rap4bQY10FPMvgJiFKoKBdIONf2BJ+SR2y7kRapnBSB3Foh7Bz8KOjyUj4
yYIxa0k0els4r4ers83GygWH1fmdlGxLVNr21WGQVkC58uBUDM/OAVz/Wp4g
G33gk5XIm+jmsWGGC1oF1DmR1zNKpD9qS88yGlMdH80n54geZCqPx3RMcxZ/
t3DjM/9I4RtLQdpOGVf+uBMab6Ap0OSWI9OOBfiXm+MjP0UuCEsjYEy53y50
/l9p6P6cHtoRliQpnKIxnJ1ZuKzZSitQWgCz0LW0JyIv/W0YnA+hB2tTIqPq
XX+Eo6Jx/Aiu3cV3qKOn6prFwGjhyLUVFVqRxYUTmFOAkJnwa5mXpjJKzZlH
XZU8swz0xX/T80ZsCGB1j3AWxzMh4ij+F9ThRiOQ/X9+uPRrFMEnONryQVnu
1VSa10OP9GvfusUmWbpaZM7OVT1u7CFlst2TdNIxe2zrFeF2gmkMkz/cpFbr
XQ1pEVpQQugRDVzwgOpJgQ2ZZwt00C6bvWWTwK9dT9hrgNaW+SB9W9GWRAsR
046ObgfpS6wxaadSKuaeFqCxxYxYZTqQopvAAMvYY+BTQDatBkq35n89BrnE
I+nrmCbkOqPWw7BaoQblq7Ar/5GJPajdGp5C9qKYkLVu19ix4WQkZLw4Z2Gz
7GRe0S996pQHM02H7viSGfMQdWHbUKIAzclHIL7E87/zDUt4y8mhXBDsaYFq
osU+gDUcVCoo8+0OIs/wTsV3BQM0bnijV9tuwhcx/q2GahpAJYtiMHdqHxyh
K4fuc9bXnW7Y7Z1N6EAQkxpRbx+bvaIP9r89vFRqU6GmhBxDdMC3h9uVknkI
ddSvZJDpBhf1Jl4jw8LSaS0FZcd1KeQoSyjhGMW2dNMcJp92kNnSFRcOgwjb
iOwr0Rg/gw2SV1ywDNH08+Du9aYQ79REg9ZvwqSrGOODW9ynapMjsOd5IfTY
J3kzWhShq9cQkuIBGPDnVMRQ4KZyivPy8uA9eABE4GBC1Oo5MuLpQWBKl5VU
i1tvtg2fIunW+ZCqT3p03sbkCKJHHPgjdN4kSnlucjSlSaXh5kbMUsf9vRV1
gE7107fGziU16AL2JZlrl+OlnueQrVtKR1cBSB5JFW48ZT0ZNgJ8A1eCPsbm
8W+s5XHh/1JiLGD8GRdB0ZbuR1ZC59KZ1WVNcxL3JjvBYf7Jh4oc2KkVt7Mb
3/VcGBNhtXNzR28ouNjEz1KxloMPjHFNKRbwsHG/WFQqUdCn3jtDqGIkAzMb
aE8NJDZuCAe4wunKC2PpMqxXRcFxLennh1pdLXorvP9go2T1zE2bGU7a/FXz
6x/RtdlkcNgALRzMBF0u2c0LrbRqv6PDrcF1GBny22BIxdaXxAgV5q4XhRvz
f4j9J3SHLwVIJzn3Fs6F8kDUxzp7KdfdAWnLnEqlnv8WqnfERqXPf9U/MaP8
m91cL3IupNeaqCXlGL2rJPI6WlI7YNO/uZnedm0EL/F2LFcuR2LyTbEkJARc
245AYSDMTrtQViQDpQccuOPYT6slQRr0IJfWsuRTswFIZgec+vYtFOTXKjnG
7JrKRJWHhKzA+F/sVT6iUssVFVixH5PB9tHKKLXRsFVSonX1gVxdNavQaRh1
jkwvD8rIKTRylPLn6L66YvJFrN3S78Iq9SCTOvXCF9e+m2cScLHO8jKX/ew6
a1KPgOqiDTac72Sg2kFchnAgW5jM8iByRuWuAayGX5l6E18z2QR1v1UjLDiO
CqhTqo4AnL/jmCZenC1S2l696P19rsw7uR+uEyaB44r+C1cVdto/6oPyxyE0
MvFllsuraiZb+5WlLnmiPVYDdh7eHOwUr3h5GpLA4byE0u/AUHH44K+jsp12
3F2rzbH/x6b65OQgw/susszvnJwK6utlh405hdA9q60G6B3nob7GBQ5Iu73a
xDzFOPmcfkbQlDx4rkdQDTnFWn5cgyrkrEH41/NRGNWNPw5o4jeJnJR9tZwr
ZG8KL6I5ftrdf13SnnCFfwemxxIeXCRkC12R

`pragma protect end_protected
