// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jL1VKo3VaOmEv0yW+3fiVTSY9qF4aHf07FQ0edzW3RV9dOC/PdejUyLDuzyG
phYdKxMuAKnxTuZ6wDDxLfMSFkm1Db5oUGl27h6IgnNUvieQjonNb2HjV/hh
e5TiCVnl9pdKk2sTMRm8Xn6l6MYQ4KOm89od2Ma0Q3MyTlBx8DskWRbHgyOS
VyZ6P0XT7uSgNLbOUz8KeyBCPTucmENHN3J08f9QoZv/hnS23I8r17LRqv4q
nHoiTJXinv4RGEEJv2DoD83xgG24MxGmedv4L4Bf5idXrDKW/K8CdzxJnASX
agHqkwq3bn272zF3E1VvvbpuJQqUkMBDWuv7DU+uyg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OHhw9mhtDO9j12CF1LLuS3E0i3yQQ9yIQScxJ5HYYlHiyt74w35KdAGEPAvD
PwAh/dfNoBzH52HOw3eX/oyacYuvQH4my/RHLvjukF6Pwkm4CCiB0bWh9vAy
CNRFnJ+HGU38vCqzixQ6PLtEYWXW2ooUrvWOiNGALSUod9eJb6tLxsiytZ0i
DmbjEd0jZ3BqPv+fWRO58ZzzqtKHV5beghABvjNd2MmgyykAqAWoplaz0xoL
J7FAy8V8SQwevc8XuEN1/n0kKzDAMqqEPSWl1bHjh1oE/UTUVZv6wj1fOCzo
BmT7ueh/A8ZCPLyORg1fCvcwcfILOfYL5/hgmUiPCw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pttd4L0PGf4Ppa9npg03ZI0SW66O5gSyaOKy1xnzNntLDPtnSOJIkBLe9LrP
/Xgtd1+gZX0YLbHhSp/fNMj1LSM/DKVe9BfbpYomUlJEQLRXeMO65jWxyZof
1EszFNv/a1b7qGcOACMFuTuSv8L5Ksjv0nei/iPjf1qis90aZar+0MO/hIC+
my8IdqONKkZPCt65wG7H51uzOlGavEQobMGOSaRwin1xNiH42vwpMD38aVdp
1ovDmcE/OkM8sN2hIUZ+A3wVlY46oJxXDYz3V/Cu3+LPq26I+d/Mqw5b69kY
l42x3OpZCZjNmD0JxVramPEFMbD9XcP6dO11hZsmVg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LJ5ECSm+bsvNlaFqZlJf3X/gM6ws6uP5ioC120GdpUvN2dKYOOuLfkOy7UjD
PrkZcClYXAbbpBPYuuXNYICDGiLV4dQWZm6SlUyA31Kh48mYr6DayqlJgh4P
hDFxS5JJCi35Ox7+1knBAf5oNHCkCBxAevwXrLmO6/Y9pvLURXU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
s6NuwV5oD6wOeMLALCZvdu8C2pOqj3Yta4DpF2PlB/7rhbzSh7IwJDIT7ABV
yC8JWWL17WrUVlBvywN5WCUlGSi08tCjIRf88Wesop8cwKDMocsLgtsC8IHZ
puOXuSXC+mpce06qwgNpW2sCIPYkHV1wVoNjtX985ynWKYsGvMPoEPqL2PYj
d4n+TNfxWtImIzLaVx21ntbzs9K4NbbmVv8go+4AfHGeHhVuxiglfUo6L2Xq
asqlFiRqlfHXwHg2+XdBAZEfTsDSpCTAT/Ub794EfP1Ut1/fKsutIZQHOmH5
veCoPlh4kH+PPUMoM61vumG3WAx5PrT8EfD2hKsohs6qwdT2Pl7kA4RASJ0I
e/XmXYiwSV8OOdnzvPw4f61yLLBXLrKUxu/D/6HYZHZ809pGC1DE3tN2xdBA
ufEZdQ/srdEOl9UlsiBjl1htQ16XO64N9pEZMY0yiPnZQR08GQu2HfQ3rnCM
PDjpbkbg9+mSzSW8qpuqeEwT1aUQB9Nm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OpvO/KJkyLK4BzgGTTVpHdo0H2G8XVmWEmLYzTl5rnF/XAdrwWRF+7lgZBXm
hLCh8hnDeHkwhui6IrxKz2Uud0oWSbg65DNXgjS9bUbtlfnDgWr/a7gLsM7c
+4LuDzC+vRDFcz5F6FounCl5tLUCAIsFmXFbwMBSaa/E1TeXaf4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bmN8qjyY/wKoXDb9wK+u/CZ/kdfCgQam18IDvRns1MpqFz1OOVAPSXcy9tVb
s4SnCw67YW2XIQkdqVlq9/m7PQeSmzINM2YBIWDoeR7Xc0D1t77qWX5IQeEQ
d3Ig0fowHp7Jc1aKBnlXt3eZVKGB4a7LpWrpWfeKENAhSYtd5xo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 91632)
`pragma protect data_block
zlN71m+Gx2idY9iKQWlaZ9OnttiBizczfyvavcsTq+1Avj92R4743pqUz0bY
k/3ymOmz9MPE0E2t6bUrR/GO2419VlLJmm7Ww3Db936832NX2foWSwzEHZQc
+LLoUCLOPv15yBa3fxZMKP/IpYJQxelRb1Fnbr56aXC8p3MKO+jnJP6yABIn
HAdLapnzQoTiG9T2D7Sb+OmN83+siHij9X/q8p5ComSi3MyRPmkOe9bEYHu+
mPOo3oh36mFeiRqGFvBXKdkph+0S8LnUo1MHKP9dm+9H60OG7z4Lv+wTUKzM
PwJK91TKh8TeceJHT3yRY9K+gQvk7/rViYRDqSb0sj0ncfqfUd5c3IwoOrso
0kBh1+WJva39DaJElIma9P9L0W2wXJxI2b/daj4t/Lnz32Fsgnt0Omo5Wmcn
iuC6qucH+8J9vX2+UP7otj+CFRpqroqpa2VOg6N0lfoMhwwlYGMPu7w25hsG
wIFGKMJ0uTk7MPHcXRWks5NrkGDB/9v7Agc+AKLHknADemUikHS3gOHVotFq
LK7zvV680kRtal+eGut8YrxPz8lKFRMHvo2mxBGINlFwlFLANyCv4hWIW4bz
nftwLuQA2BXnuyUQSmfy9agYGt0nzKVJ7qSQdwiO5sc6nsWE0GF6SDdd72Jf
y7Dq2JatlYM/d9A9R636s+K7bYvtcqiaQXucBOyo6WDMrc7kUDGX/z9xlTaB
KJUy2k9ERL/5LQY8V+aQOPvNaMAExsNIIECocWCeMFIU4lXGAlHaL/LODQV6
kaY5SLYB2h9XaTUTj1DywE/FeW2pFYCTMGkLXznqf95O3XuU5DJtJt9wf9Y5
K7q8j4EZzX9e0JXrcxVITIQ3mzZsPoRUwjQCbejMUS0ryyIYqLiyJdBUeqzh
FCIKP8y4VYSBqmqbleOliOl62w9iROVIsRf7XYxk+3RLxYAzO0iyjAyoaQ53
wMm7PvWeJIUUR416dHcdgqfLWVcDLoloN2NAzJ05ncSnca5lwK5W7R9Nj8qR
WVEWAV/mhhW8lMPke34yg8myxxuv2Ud6yCRoFYfRIVxpkE5+GfwjpI2SoqM3
fFIXl2xaLISRE7GbY36E5N8cUp4d59G5gdDzBZYsXZHakQuJf9e19Wm6AbXB
57CGVLGmDVTe76D8XaCY+NENl8TgHczKPElxg4Yo+Nn/vV1MalWERk7kQSTF
YQL75lLDM6QpcuCZSJNIGbXW/IAQFNN46TULMdoifBmKZVp4/fjrJZ5KSVXQ
+q4qYt2q1VSSaxEWbcw83iHEhsiobKYNezA1PLiszD6htYP8st7v3G9qfmkO
Gr9dH2vy1zmTQBztOpZ8JGc60ub+52hq4XxujWbsixQpMiE/YfVqDtTVOSpd
cHmhgEWELx223kbVN6uDE03UJNyEZXd1b4u/GbnZ3mejX+yIj5wyxeFprNAJ
6Dmfuqk4xiTkzs7QaHWpxLtKUxnmKcMi5GoCp39vXLWfDHVvivyXR8jowBSM
RHfwDoN8KvkKUAhBgekbQPkBFuvh5lfrxEjZHApaNzq6GaDs0wFQfvIolpnm
VhsEcNWrWRQjhOvfy+p2p+ut6Q0bc7fzd7eLDoFqV4mSP9HjoVLZCvU8JwXe
zTL3lvRubxbhyPxNi9+fRv4OrXX3L28KUofNzAf1HhMAk7EwVLsOShVA0Kk7
VqqMDCHAtdP4VfyvmEeJ2F5+qt/EuA02TzBTuEh1jsOblHLUZquKebDwnqvN
FucTKKFH2wI83Dq7LNAxykGDmc+CZBzxR1Mz+M7DXALqAcpf25mxctb/rtjK
ZrGfGQyLg6lDf97hPLehHIySX41sNKDjpe0qD21fDQMk+asRMpmNe3y7pyYs
9in7/2jiudyGpQo+Xb+R+5oPwWoh8eGCvR50EU36ryOzmgeaTAnglyDVplUA
IS0Brl3r+BUcwihWDvuibx2bxtbOnHpkL1RzAjj8hUg1Uzlr2NS2WMEtJVv8
CuRlrx1qJQO3STis6QBj5qyvg4ePWwSKG2Ik+kBi1UuY3Ldy/h5HZRiXPxKx
YaYU9S7FfTittveHRa8IopyyAQaMJ1CapejDIEZKYlZuRzUKBOMEjN2CjCGV
SE6MD4O8pddOs1a63p1I0/jOM7z/em7FfJGX9IBjpTHB9dtdV7jEN58GowPX
/5yvS1fi3oFJzCV4+ted8euvkeccRjv5cVb0yczhtZsApdK69YvmUtlQWPQ5
HGLYHt0+pusjngD2gdj8Ym8JelnWfyxs4+8NbIhUL73Ku29nDHsxE9CRMj3z
OWl229GW5BxeNGDI9CRfWk7CJNaPGpveYiaLO3/xX1YyiyAlFw0kSNQVFwX3
lhsyiZgVCV+9wEutC3Nx19cdrKIs5oR9HgNnZMDb8f89T8pHtMoF1c9y53aU
gnOyTF5Va4vzKuVSHPEmrH10s6CMIjx0noQ9yYBGK1Pjt5PKNQNUkltmeapa
1A+XLLkHyvMUFFOyhBIsZElvqxj5TnSOLBnDXKS7jzjJRbbCOheLdxAbmhsV
S+qJvk1UjYbUkKrP67cq9rFK20R96ieufqj5+UhxBw9/8g7PlxA7tGcgqp3k
qjTT/+qZl+DPqeRPnXBE8Lr1ggQPTZ2VJR8pVnz3aRZoR4SSy0fmkDacIcHP
7PTEI1AcEjJoyhs/GjcW6sh8qv2ypVfVkxOZ1aYkZ/DeYTpfMIVmPVGQqDS8
1Wqew3+056KLDLf7PSEVbmHFs6KrjwTgKZLIgVtBjIIcQ0nnNvdT5D2Iw7ED
4s6FsHPhP+xr/xeYNG9cOOfk14vij0EIG/HqLQp3vHRs6sZzdl6JD3nHZ7Js
yYkQeRA1k4x1Svg6Yo4YPSOIoLzou6mmiNG8WV+PDBOnIgGWVbFZFWl8g+Pq
6nk+oD+tXsnvAX8Fjl5eIDnZYA6+MGjek95gtQ2hB9sycCgw4ML/hUc7xi0/
KYvrucnhgL3YqLvK7CmU1khb+AH4gdtuGGAltflra+DCcbkigB4K70wIC2gy
xuIQXkavqEk0qckqA4FBzNxyM8FMmvkczz3HobUMFJb+vsS93w229GXjMzAx
QNBI+oMmIFCltowfQPDyAp6liecTk/dlbgT6Bkfbhe/FOzLV22ocNa5ZOpOZ
38OS12/R+KKFUARvWq5sYgC+dl/UVrn+IJ3adop5+tRf5dcVWv+1AuboxxUD
k4YO8CL+T6D0sZTLryYsa+2JyZfoUqgFWnKCpB6dQjwNZho5rpDKW7bMGNaJ
MQZleh452c6545JXJSw91wpqRdpmvDgb40uHlXSoTQB7drckMlCcckJ597Zo
hQF7UXwUOUdwSTphCIA4qVhZFEobVgHLy0zdc2sufrc1T9OX21oJmYnRkWwl
qK1TtIwQg7t4oobTQDC9TKJMtEq51ZYOt1OPb0FTq9x7FpU/g6MBgvpvHNQU
1T3i6oCheMuEi3lrvffAcm0uRf4iy6Z0dx1wQMZUa2ggp4aThIr3AyLE56DF
nWvAvJbz4RXNJF1LSoa/uBmmW/MBtWuiaWROHahQlgZhsFdtjZCvjNmCqM6O
fgkV2tupkCYgCpnEelPTHmC4DOSQZCuUxVib3Rb9Ghu2ijN5z1sxAgywJGAG
jJ55Sb25A7kG6H2rIsEqP/J7HncAAbKldKponeZcxHox4gUqw1EhMsC47yTV
3S6abxkhvTwoFuih+BxePO+a2dAukOsizZdXCTEQ6rlDY88g3ZjrWft7t+cW
hh0G76iaWw0UWc45ChdO0NXcuOm13BkWRpIbdw2wr9tWuMOwZ4UYaqnoOCOZ
jhLogVQq3Q/2A5ght6QDzi95DXr2/wkhjY4wAaeCve8hdLNTciPU551Kkbpl
JcOJtiltUnYHUV7ZMsOte3IdFidQwcCLwx1y2r13JXXoRZNwuQsszhFxFEeS
MlwvfrOVLk7LexCkTEG+FzpQFQMoqgu2TDsg5Hk9Jdj1KxQF0otNTq/KC8/i
uWMigiZpghpnOiXGVirzHEHuMQLHxMUCH6iQ3SyUUxnvvZspDJv3DOG2aBx3
Ay0nbRmU2+hkSxN5YpvJ3/Ya71b1MOSDAu6f04LbQfapXzz9yhtKJYRTtHLR
drqwmO6+fUIR2YekGSPcLA9atqwWFjq06F8GgkuQgZCvZ/IKB5TEugSIZzob
G3gYkYcLFLBIAtmSbDxjeZiBeHmySzyFOy5YNXaR3Ww4nOc9T7uKKTzqbRho
6fReIU8Eg11XVKraN+F+uyZDSAyLy8vDYIaLa7SPIVVFAeuFvifgYArR6V0l
a876kUlNK5XhfgR5jbTlPUVU2VMfffChISz31jxxE05qqZrvcjfrcu0GIzch
TxrG1lIjiqwQcopbgXGeBznRJo/fFxJjkUTgkJM5bk7MDZz2DjepH/HR1f3T
kwvGIZWFB0SoN2dr8BCBZBj+T+LDBJvkG1K+d7w/7qiNIeaZvFgmtKbavCoz
ThoIEHeD+56veIJEVX3M9c+PKi3zgpwtp0BNEOpOE9klKFd4Iqvdc4pLv2Xa
Lfzprf23HKpvSX+sDoNjXeoh1EZZu925VakIQKImck/nSuuVGCmpqxWzDILu
5Q0KKX7UABbuBvbXtYRY1CuX2uLc+fQTPjXFAUPpvWk8iIb0IW5rzMzAtyfT
SfB4PH2jor3QP6zTgDkCL5ZWn5+Qo5nSNeKAcHTdQdOsnuFYNJSpXGGl4kuB
z06FgY9T844tadlyWSqv4d6kMySFfJRqj3i2KmQfbrWbXG1U+zMBb5jzVUB7
9kpRC/hu2rOPeOXhHBTKzamct4cv1Jz++//sVHvbWIHWdjsqgvCKTPc9+jNc
+E7vxEYIqNu5JgwMo0V7csvOCTvzD9DFsmhkDZMe62I1LYwQiZmwsCv4Hjk5
2ec1oaNlYG9GuroYqCFRyH7T6x1UJU6G4SCO+G4wNokZaAvBT6fj5Acq7S6i
dFJ2doyrP+FnNYdELdLV5581vYBxS7GMcdf36FQgAPcQ5qWkUJK1DLHQ3lHc
W8sbgd71x1WvdU+yZWSTpH6eQhoLJ5Lc3DehuVstZ377odB6Xna006wKvwkN
fGr2GYtROSgJPyp5tY7bFNG8OtF0Wl8tuyXOiRnuC6LxYf89Q8dXfRvhRQ8g
jSTs4n9bpbQWzJ3ouwemFblfZf4uHtQh/YDYlpvKMAiQ7hhzeQoZmxHeV98p
XxnI7Oz8gg4ig9GK9OdLHVVtR59gmFM75eIb26tKCnQ5y8SV303qqA7JHZAy
DKciVbH3Rpvi+gXpINg+nMEISaCwvh9SGzx0t5lQGvKPrf/k9jhaq3li4th6
a74QqjietLiHCbPXP7t03s1Q+12Ai/z+QhQRvR9yXxoW8A7PPBukUqGPklGY
HX/VGcphlQMXSZGvwP7KpEcYxISTlN+bVw6GufdTtIWbpZsS5Ak5ATlLdjea
seLajlfvriwNmusD1BMZfEUOS0Dh5u7Ciix/96X/ao/k8ANp4nSzb2oRvVWC
WumPLLZIhwHIq8BqdY1vmQ9QSj7EChF0kFmfIK/xJEEf96X3ODSwty7RzI3/
rCQ/D5JobZGRVo0rT6uo63dDtpoMVo0sAiIGDAnWmI0QedamF1tUl8Qhi91z
YV+0ggj9ZbMB1Gylgkx1snpJ2jbJWfTeBom+Wa8Bewak5XMH4kNsEP++bRGr
snnAQwkX9UYSS6sDkfQA1hLBb5fP4706GSvMgbHeFjmPLUA3gvARbcz9bkNP
vhat5ySRRXCnJPEZjJ+zKpREO2bA56cz0+6+6M3hs9nZez2XEmYq1x3rImR5
LP4GccClXpw7yJC0PPfcVHQur9/4EoEPCpOrspg/svvyWJan/5X7NJKnq301
S7W2FmlOFR1P5oYmU0T63tVcyPwn3rZTgpcgAH53ffhw0QVuO3KuUEJD7WvN
9CU/X++3Hs/LVKIAKKPUkCdgHQTXOJNuAILifn0ZQDhJULzUoxJIl9JspGY1
PHKVpGfZcbEUmmNO8XaA7dIeCOQNjWCsMTYEFkRUS3bXQPND+/l5ekKH3eGV
HD/P6Qll6o8oyHlJ1Fqfu1SJgk0/+46kHTVzSdcCIeIPSmJSG80ebF0jtxwx
CqjX8IWM3XHCMN2NnJmW2JWO+evHAREqZ5Jk/p2sJDS6vydJZalMid734P39
dVSHUoKbIRy3DiziDlwF/t4qA3O2fatejQNlTwdvnXsMg+jXsLbtYWk4THfO
EdGE4M3jWLH2eBq4q6cwM6hut5ldOukv8mGBcZl+Ib7/xW9AwYQaC2OEj9lC
EzBvLYSEP+1ACbaKH10FkCgMVEvIxT+O9YTkm1ZwYlOjkO/iEUFIiOzyFBCO
jd6SL1F4xSO95jmIKlTrDenF1LM2sBAcTLqQgXTntLKyca7gaqq1njnc5dBj
oYl5YCrVaHWnABsDBK+lgXAVF4bRObenJt2yc+CzQlcss7crVsdYcex+q7Pp
WCrPw24m83M/4HpA0/KGUI/Y+kld4KMtqn1O/F2X3cte4X0t7dFZo5I42sMy
VGtik7RMwcfh2MgnLq9ir6Q+dzWz+XEdC5fApR0Se7RyzMfNq7LGZn9Ig/OB
hNucfLtFH6Kscs48an6vYsUC3DtnuZ3Gw3PPoxJfivUf5oCc7KP/AXoUMqX+
BpTivAAXCOy29EwLflTjy6B3CSiWtC1hALiL/urUvkTn0+cZzPqeklI99Ef4
5JL/GIfsj7vd3q3MRIi3YVkUz63nGeseOTvEWMSYDhf1Z46r2y1DCSjvMPD8
qX6IRWTfQBTMha7276cMoLkoNjB4hzFZb8RjgkfBEtckkLTG41sMHIboClOP
HmxYKqSctEcEffxqu2SKabGbSzz47NEr+MErSI/vVQP35DU10hP7l7JxD/UA
cD6CIurMrglYFj89sG9mTiSPemO0UZbLInIbd6pN6GrlbmlKxFSUVHt3wNHV
fq9Xmm171O+rfEk2zlzAHX9+GL/3M4lud5GM9BQNG2bu/PU+YRybKyE7bv7S
kTk0Srg3hQqzkV4mJlQBd5ZQI8W9VscRVmQy7pZUbA3T2l2aYHhUK6Gw1OK0
MCTC8AN7wJY6l+xF3kKsBCNGOug9wxWgoU6oPezFzj4KzxdnAvq0ayXcY8cX
uq+8mjPrxmJBd0luHy/Zr2uYZyK4eY4avYGA4hVZD7Cg8Iugp1Ziu9B7L4uq
A2YdpS6ltPgwHx2Z235i0tE5NqB905lRr+5tG9E7IgFtJTRQoE6Ie6j8UocL
jOLopqT6+buWC7sc263x6UH/rufu80KlODRxC8c1ASf2etNj7CsNJX7s2epC
/AcMEjJoLuTprUKwNW/mZeHwsG4Bxy6Z3Vc0Nes3yECXPj4XZcY1DzQocXgr
sfCgg27A9cohn9Xst2Te3Gb2ZCB854t59Zl6pSAldemv+LybRZvW1iijGy63
ORnUNsh4Yrv1vGwWpMKyb92A8hPwxV+QPRQzAKcj+3+tdfNgW6eEmFVhNPut
T9lcCitXM8ZejSCqtpvDP5bo6QDP7SDdSvdW7lzY4IOlcTQTQ3ZmAdGTlb08
7X/cvwsa5tRuGhTqZwjWUp6i88jxAq6qBze5/Ht+0XjvgMSysYbO8U9j3QNv
FRXmsxFRW14Byie0dPGlivm9Mb/Jm0jmw0Mzfta12uU5gadQoDj7KyFa0jB7
c2KsuLtL+/L3tzvk6jepebZGkjJmV4090kPolmqFaBiLmnZ4O9bGoavkMIY3
GXpYgFprGJdI1EQ5NczvDmDoo5o3P6ZQgaCm46QRS4Jhlo1VGwba1ODjV1i0
eYUX72Q/QAd2PD8QWi1U6azqY6qX0Z3BlGbx39CREKrz9ZRnvDpWZgXJhlOJ
C307ZMarseXKbgfWWiF7roq8Q05b2P6SPei5VfdDh4SAJLLennSsko6XFumB
gThMpti4ok/j7wS70tJvABhbd2iGANBlZamdHjZQSlztaQm6dZuOwSvbFO9u
c18U9PQ54eZc5i8MK2lCCx34XjN0C1gm8Nr3CApx/JeC5KjEQ08Er445Bnko
8dXyKmVtowSbZ/sJKfVN0JHhHH9COqKOaoG7vs+FUzocjXZQiNkMpqtY/R/M
3Q4tFI7gg/ayJ1AhDrP9u6wTj9r3vQMEr45K5t3TXOGrGTeTA12PYnTdMwix
8A5GK8VVkfZrMb/8S4+7u3iEwavuv2Cs3HBYCVvk/Dml/BEuSa2VBaF8a1Az
UGclBT4bUDJJMEY3StCH7blXlVCDfgLIbm5wFEe3odpRau87iuliIzYPFfhm
QdMncK55FYejiT6Z+Jp6EZ/xUrMv/+OR9qM2iWB55NBiINuqVJ6Dt/mnem/c
L79q6ICSxKjqPeXcNBnGV7WFlsZ3AX9+EE3Eadh8rPMQ1LiJJegf6I0BqgsJ
IoJKGTYxGLSEwaiuXbxgu1k9GKOr5FoYWwy18eXToB23bWjZ2jWNmJx09rr1
JdbWdhr+k3ozDBZbgf9OC59Y2uZAkFxdpek6FG8paMDi1Tn8LxVDeah11bO0
gRVkfkiaHjsFk4x6NaC27TJbUOfd9a0rU6Zi2U8zzdrt0cPleM7ebSPXG/zX
pIwzbdKh3SYUkDiE6kwMeEJXbuUI6sxlEjtLAE1Tiw7uyzf6Fi9+bJ5m0Jzt
qAEo7xL7ISxeRozfhhtl9AJf/8iawgTO4jkmu8F/N4ujokYmrfje7E9nV8Oi
UKaqjpTSpBIWaF8mkbhFFUqoaNwnEgkDXGTdi1M7oLXEFiJ3f0CyCAv6UcPf
XbnW0Tue2XiNR1ijBOfvAI0A1EYH62X3mhqpt4IO3MsPPBcUTaExOftnNIHo
S/ZzcTEYfTpLgVqSMDi/ULxd263jD/tuDu1400U9+nFRsof4eYqRE/HA+jyY
s6O4uAMe2NXZRTszS7H8Sv/cQBs6p11+3RrqHqu27fYpMsuJiKtss3jsGxzc
BJYAzKLfceKWxLrhfAxxIKp5+ewha/1VF/5TwMVMJrpnj8/CaneO4KwQk//f
8ChrKRaaCgx04hTlnjxbwHYEVvf7+uDSdBd8Z0yVUa0D/CueFq7sKIvGgeHN
AG9oota3NovT+4ET5jtfBzAQp93D5qv7weW8+xhzew6gb9J3cGxK7KEVPrNj
mrFI3Lf15nXDqKQXoz5VwLli02CHPGPGHcDnArd4dPZRhQzJ8QDkZJupWWQC
YYrFRVEF1GsHQ5CNQ1LCIKBODrYMQy7mxiHGbCoKw3LTqgCQj7AfJvjp88GZ
ynnFJYtyQqCRzLDriIIefEtIebDlzmzd2lPx6X0BTNanefkA+4HZJBeb7ia/
FMLhI9IS1y6fAsGGwJIF5dn8GpyV7SEiTKQDbx+0JVU7tMue9+iWdLYJ9CbB
NppWKH9N1S25Pj9Mt0TaTNy0zrmYPj9DsYWLkwsXZBwJjX47y4P+1pA60ygX
3X2wTFNQ1oZqS2PHZ1XDRWME+GO/0rrO2aEumVNuF2w0d89IMZ2ZgyA4hoLB
q/0VZ/sb1NzfCbQHXjnxBQKdhyb8F2h9kaKMc0ladHKyffLNI3dQspG4gcXf
rGpHqNLB9lMY43TY3xssSpmwk2rfAfUvsVb/G262V4Ee/HwwuGW5P6GchLn4
5peNNRShbbR9P7rYQL1/Q55SZGWzPOf2r0PtgRGbthrsL8CLxFtG5j+jCYq+
vOGa9XuGuxXe9Wh4VM5LPu8mWP+lRDAkBs8izvW6uDJKlc0oyeiWrNCYR6IA
RhOsXbiqcw/RboTT5GpmrmTn7BGsGtXoJA1u2R9qh6kkHxmPcTkMQ8TATggu
K37p2NVL0Dvafk7a9B4jzdNZye7QfjpOfCfMRvFZqmRi1fNkG9wHieWIsY4H
6QCTcK3x/cwVKVCzK8r7ygVk5TpSeLhNNkkNxTrN9UfJPb4zcqT7b3/tjHdA
lJtNtEtlUCgSaB8/RA1Jn8T2XifnsRkdWwdxaBMzkfdYUqvRDsq6pIuSxLcx
ruvGBT2aw3dfSuRvDAGVZUe1LF6gyi2o/esuQU2SYT/IeCWXFqlp0Umsj/zW
kOcT/Qj4BeQvLvZiKBC8cp5YyucUL4xNfxWV/yyyjw5nSCA+mrLYYU059gz1
7szXTuADSr7OoWPXQwXVA6U02rvoZnP2mHueqsx6v5JVAcZ6u6a6w74aWw+G
2IP3LgoaGVBlZYWyvGnTDNyNXfTBjfvVwSwGAAXAaNWGaIAqqSjdUr4JoOXw
pSdi0B2vAblLamTXO/WJi/og/LRKXjOWNtgLZGFi0iWFV73G/e6j6/sNQlUL
dTmB6qhiFbpFQi6Gh189Fv5cbz2cCXNKof8G20e8QHDUTClOW2c791rAVLN5
8yCjm8vbstjW8j9WZrR625j2yHoO/ObhtzGH1O3s7OpUfHFfRkUO3dkAVa96
UpO9Ko2Mw7rFaKbLv/UyoaibZg7lg220+UM0csO15INXYetz16BmdBDU7Z9f
HFoGjy6nn/bPqYELaBIL2tEBaN1K7aAjuvvCa4zAAz8QaQfVoU/b/beNdlsg
7a/xo1aNvRbHsBSOqvWQV02UM4OK76WIIDjNkS4JRzs0oN+m+5vEGesVgFiM
Qr4ynYGDI0+i0KYK7//AlhRRT9D5oscmWcGzH/slAkbUHwgToH0RaQR6sYWZ
kjAKWGFxkFA+tEX7T+gObR2W04GRMfW5/vx4qwJ7S3nhvtVsVIB4zMGEwTmR
FhTmBR7qC/ywsdUbX27WeW0bR/Up2MfP6aSP62fBnw+B/Kal+zvk7VSn9gw4
fq6QAog+kkAuYodJxsVFJYecLY5OHyBQXu5/Q0yFn9UVpCENA5RwqHP0K8LZ
Hso/J09ZbUQz5XO+woLFBhKUWpvrxtZUtVQHrEfOZktVQE2hRxzrk/pF8pqO
AyzGoIK4ga2XNkCS5ynfyL0jra2dq+wC1Y0i2zyJQXwNNozbbV1xZeKkALOM
5gw/bwh+rkvgyzTTvHuwslN1cKEekAdEUM5qsXDO8m4KZw+ZT9NClxrZi6TC
3sUAJX4Y0HjOlqH5glBl3kPACIiOjbgnVykYq23btVKMC6eUTxH8YQ+niWd5
bJVbsZ3INtJFBqXBFmZMAU3yvNHdhX3muPZasWQXtbHWNgqWWWANkRu/0hCp
zALV785/FQJ7h+F8YMKAwZfeHSYCqWZdEy/hEJHRhLXwrM0OWmBzoK33qnGK
JCwlDdufxxlaFnmIaBjMHXEDBzu8lv5dFs8hTX4yYTQBee1Q0+qxzZTlHiXP
tQwUY6VVM8Cyatg5G+xny6cHzwnmj9L0iKpUiZpU34QKq+dUvlbM7Eit5jrI
d1tK2YoBMepxYjTt11wTnFCEBVi8LCx2KdtGCsup1lAWHAqmxD9ptJ774han
R2J/t+Hj95Q3QmLMVT/G3LuvTa7FZjO5Izilr3M994yrpP8hgIS9j2Mh91UG
DrNFalroG7mddLU4lvu2OI0tLAaF03AtkxcO9uhtuKYgmYkwQ6bYYmqqOxNr
4x0AP0IDA6Cfil7SwKNcxZ3LpN9NQyfzZdvmmZEeQzCe7wVvznJIqn9t9tT4
b+fokHQpYVbIG+J7PL5yVGeqTblj30xm376opqfIVyKdnbdbOWO8GUAZiN2C
NSTgyTnzxnPmztQZgGZf6DzSQ7Zcp4EAyuk6aTyTELRwVouW3yBdsPO3d2IK
FzNBYAEqKAowWMcmisZzbrHoBbi/BtFXQCC4YOjfl6ASESCiW1lS9W/TF27v
qKIIhN9wgMLsUB9cLO8BE4dt8rGmKQKY2Ge04l58LlbYAXTn0UT0AHl5esDO
TMKt0xsO4lygiXmM++BTGW6CfZ/mmNasyJUW+Fp/lWBBH9MVGldD/eYsqmJk
f8lWT7/79wWwwtyZ9ekCUl76mC0DAZ95fpgvBag5D50vcQrN7oRMFYMZmIgx
ZZIkzuXrYe9FNdkXdjCegyp13vO0xPZn+ubAfZb09Nw2Zwa0Jhv4Y/ZmzC7V
ziJCowEZQeE5M42Fwh4G61BGidNvTYxLO8t/ihuQPj3eXwdOdwvPWsNVZkG5
CrxQiSxjQtYIpqTWdd7JT5GuiS3tk/de9MaOczGYKPtKgvU3XvfcufzPXBLB
SpDBO8OyQq6hQ12nGUEHd1K4mkfm/ccLrk18eajDCqy03P3EC1Z+xcbMrjDk
3AaKYhkCfkA5FDb+PSZp6yQCH3ZsW6Y5TVOYQiiHpiwxB3Cg6zhA5PMKIxN3
OKBw3W2jDdUlbw9JB7du9kIbpgMlzgfHfQKLPuVJd3B2GagRGjXHwOOY6RuC
aUGZCAFU/pA4MYwcdrElOkiAQhvIzUL3DmHIcsPqzeqRDM1BgvhYOr2YPsA3
ey5VxpGxDArAYko/a/rWusgCcBoZ3r8FdOtjkigjwte9DlxN1jZkjAOlxORm
X/IJhGo3wro2CfrWe86p43LxrKFFUwwwgNekG1e0inAN+9+vJ3MzwqXBKi1e
XeJPfcyCN9s1dPhcrWHKE91wCtMIpASuXtNnB3MARZ0souWn62lKE7z5QN0M
mHK41hL6IkBHKFDC+Swp1fO9famSKWOtlYwB+1yJHgE9EJf61KnsolrnIGol
/FyAzplZq8HSytYLbuPrscWdJ/PyadcQ2LY2SzsVtg8FnNmAfje4IamRjSnT
2L8YopDht4V2yMAEOv4NAzml0msipWu9Rye0QXmeNia0L+1sicszsSBWvoJZ
jR3jHS7k0Ie7JxYIiaHsCAaVuqog08sQWUO49bbYPwBBWJz/ja52rIYtBhR2
x/btVxSXkz+nzebah7YTSrLQDm7uHWPVi1ZevTpGKgvYFiYdqjZGWB1Rr5RP
cIu2gRCP5IRr54EgFbKwQCYfaiacpivXq0/vLDplK7EU9Gb80rE9pd1xxqdx
KMvTLekYdDqAdC8WS8Z11kknJ1v3Xc2plQjYUhMVFShESekfMYwCskmZUnm1
gsmpTyxObw+iXndRnb9Fx+JfFV6BN65Q190WbZz/V0rqvpB9DfNNH1WM0Ky+
xbqWER+D4b/M2YE61OaXErcJI2vGvgVLRQmltvyvYu6XC3z+G7jld06w3887
G6VQPdtdNEU0rvgyZ/R8aIIVPUii9kuy1AZLlxXUFQBOOHfkpL242P6DUYKo
Kt5VR3dY01Frh4uINAv+O9livOQRsqEjgcSDAInkHHDun/YYmMaduxlPiASn
0cE98bhOFfmHKDhEJyNTQltUIJuXz+idDH25bbWwWYe7NYPEv4j8wK3mtcwe
XYbIXgmheRDKqoDDZ6EbYjzfQpe5WqjEXBGDpsY4XwYlPIJX4+rAN2UE8ELp
Srm2pOcWGzQ/79REhBlcT2ySyFQR1ZYoaEE1BTce93qhmds/dfUqdlC97d1n
Bv9TlojcNWne0pNUzy1YdmzmgcbgdCZ5Fnp+3lPMtGnhSZpDhIZk5Pn7Eqcg
y7RrlpPPVLmpp5l+Odmfqa2wHaEIC0N7A1Z2Owjpc0hzzEarEJJKtcdLHYh5
hHGf/+PW9YTfgMPoJ/8pk3Pi1bChMUchlchN0+YlrFyBNDbv5y7gGqRDZ8KM
DzBIOCn3iLHpmtyDu1QpIUwc2fNUMxGmG7O4x//2UjlgrOGbH3ZXTKxLe3Mb
XwV8aH08XnIfwCu8OKSLXiw/DbZSpbSlLAyzxCdXHUoxOlq0bfu/pqjZoQ0q
LnRkOFxwrtYCuajBl/uVQD9m8mCFycRXZ3c2TACBFQOfQIzDrHuItIkYY7Th
+cYxASnzlQmCC7rS5TPO7daQWu326brMNiteTunf0Q+FWEoZe7zB4h9+BIXr
uSGSKmzlG5PfJQSXc2JLMlIPJU/wTlNRAp9WvdbszgtBhF5qymiiCnKdZL0M
bhFz1bIxfq8maWLcgMcFnAZPoDKW2AQRFBqo5LhJSHsbpBoosoU36PHu+B4t
oiuYSUgHt3if3YVGXNLegPKwXYkrRHeovqL1rODDrhZ9fJKhmBV2/vRs+SCP
d4bH19qFCat7M0aSTzv+r3jnQE9kOT3uGcmAaZdLuESL5/mKhhcPiz6RWy1r
d5/5z4tmYfndIF35z8CbAQISyKf9DEUapCXCqE8dOMw3DbKoWhGBsEGVhoUe
aSx+gXemOq5DicmHWfc7XqsoHRxu89JHBbJtOrU7mjFGss9RSIM7j6/5tED+
GnrSGhawviZ2X2CMdY7TChrmRFCa2U9W3fuFMcuUA/r2yELXDIeP/HKd3wdT
5pmwZ5IfsNFhqH/qiVAEEkm9kSOk1PY4yhBzi0Bc0VibdDklQuTAfoA2sLRv
6Rw4HUgQh+79TilDaTNuKNKV7079VctTppDQZwIqKpWQxvk3f5vSMmjr01jK
3H0QQ5zZqG/CDyjjyfkC7LLlncHRIrH7iXxO5suLEf6k6txwmpSsXeXJpZNj
m9Rt1XUTDQDSZJRX+acMDzdEg9LXLlNcW8PWyJEUVy/FmAwueBsk84jbAYgB
RjzZh7SBe+7vOxA+3RKx/SFS4VSVydirFDy6FvVP6H/1MTAMr1zhSxbDsn6y
EP2F6kiOr8E7UuxFpFVyL2+o6thnm3ybI0XbWNr2GSyWcNEaUyqv0eSNkUgH
WkLHZ/W1fUFxzWCw2eYvzgXG0KN1LAETwJoZlU48SjziQTNax3Z2plBJF1eO
t3B3+UdmHaeAuUVgdZP14EY9tWO46exCih3nDKkgzOBy/7sxjV/1U4+rCYCq
/vAE/xgIrYoc377znYNcHYTVG2me8BdkHyq8gP2G2S65RXXHza+QmW5Mro7Z
9S0Qd8A7Ze7zIVR/LICi/2883oh1oduh3+cgnAiar1G+VmI2ijidEDByY84t
n+wRUUOE0LcGU/wiThSHXxso8Zmn/y/1HhmUjUONDfCLdUfaSERTBUa3w1lj
jVlvSPfqhW2+QCqvwzwAw0J/ZyrT1Aha/fYeBcGSKHdOZHQRiBOYW4JBGeNt
9Upyl+UpJO3TjvE01uBcCNMhhNK4rAFY0C15AsffFF7tzDYuDXiTNq0HmFDM
1dDt6/RLssaekfqkqKeHIqjqwQw5BtjUfbOgiqCKOlUGeVuQ0RKwSkXmIVJb
InJUURNToBOtq8IfpyMABuHsDNuLow6A7NT8WvJJvKMu6B3Zgq3DekeoOz+r
MdeFAau7kqk9KUXfQlvmpcD0oUiCPyWMAkCOp439RxHGO2EiGWT4dy50QXIj
Nm9Q4MWXgJIoV1eoChkY/0fkIbmJpI43RT0brvFfWRjCN0ZBy6ARdK6SA/As
ChVX1xyUO13egY6ue3/jWXWJoONuqWZ1XBR9ipeogW/ysPr2uZlQKD+If9W5
aJXpk6up6iOl1V3bU58F5qENrSpJliyJAf5aIXJI1cY1VWWX8lk54OHAV/NI
zjoYzwTnWlt8qlfU6YXg5nKcKhFZAnqaTcFZsd3/ocCmqsiqyCeVYz4frAeR
Ulxd323d574zlUizYEeBcHVebtGjj+9wk2AQK++l/PcEMRlrgsXiyx4U5fa6
3qC6SCEDv+D5h1I1iI6c/rD0qPLPn80LET1MJoQ6/NpaFY9jmryWt6bnQ0OF
K31E+loXnfHuHRK1sC7Xrxxe3/L9SV64zFzIuhv76s9XNecyEcM4jfHDzM9A
btqN25TZ+hfs+xbKmrnkLaeh4OjMeilz7QulrVpAqiEzQVxH5mDL6QS8qGEg
3+H8A49wARLwlCcQQUUZsePgnAJRGUt8dyDT9Rz3oxGPfjey5g9ypTXCWkXI
w8MlLLUQXMuBPdFIk+KjOfI1+f6ikLpXM3q/o5oBSJMvOxqoKkBsQPlkwYe4
FSjDjIqWvrF7Ed0kcHc4jY5orC2lwtrDA+WClShS6D30fjDzunaMVvwKDoA2
STSLJ7JpKsygdONy+J31i//AurNOzHq7/rHkXQveyCxGzjYb2DJHH5ukvfy+
om46fgEO4243YVhiupqsBx0ff5NKmAiz8EWaWnIh1EMkOPUNYMyZ2elPbkHB
XkslW9mzW1QbgTuD6LtwX4puB66CKm40ocovnHch4pCJ+drPCW0drLJfaKX6
mYeJvaghNYBRGYFzFigNJHP1DLq13Il3J2zPNAvi9YwnLgzgfyIWnbl+xmHs
Fq1PGLnaWzga4SbKLDpw3Lu1ZwHMHV2cBiMKo9HReB4j8c+5EQkc4qgvZGCP
KDAcdGm9m1wEJVr/A2rfmiNM3HwjIBq3L0SCHGD9xgBv/54uEJ5ejMsX7ux7
5esCwNVhGs9qdFgUo8q6yC4HefMxdgQVfhMJ/Ad+cePYTo63qgonTmYoKnO2
tqNHyLhXCDMTcF5/BI7JhGnNJk9U79rAHTlB8BqjcdLKiRysan5yHA9lIqf3
9MVXE7RHS85W01JPI/iZAu5AgQEb4RVfTTwZFNidTbluP7ZEi56pWNuNgQLa
m+0Rfr9YKFrwfAjQLbzHRjLQXlGdEVNlQ8alrsXLT6/js7Yw0vhlT5IhMSs1
2BlxvY8bjDbdhG1qZ2Ecrq1zAzPz9bK/iZZq0gxyQlgxwYhtLtHyGS/ub1AY
/XOjL4uARkrJLdelni4x9JFfib+rWInYqp7Mfmn7+LvOFP8ryqUuxrumcgDR
NBcyE66h4VBmnLIq5WpedCfBV44DD7qKpcEtNRSUMBsUdz9EbDqSX6kTUdwl
YgEivQVmlk5g9baICx1RsyZhbLOsIRJ/e4tJVIrafnDgEHYa3yUMajqKw5CO
yf+WgH5RIo2Xt845lB6+Gq+Xe3LPEj4y2qyzk4IZZ0v+BK4FmFERd+gaUnAA
+Ll7nq2p1ELzGczZA3SLYwmFeaXE1skSK/gDJ9WGERDbncLlCGyZnV/Uaaft
VQR5Jp7jCn6+VFLQ2SG2ncWXN1G3JKSxuzZrquEd8TXPqRd6XVktmmFYErPW
b4WZ7VbKEMAV8Ea9WDE3Q6K+oVTjWUKcsesWFOhmxjVAwvLZ9mDUez32QyQC
SkQTfNyB4qwoPR+NgvoqhG9IZxWpVsCcnYK0OwGNJhdKy+cFkELm2ZDVIbJt
I+2BwCxeQP9KjEijjONO07428PE8PXM+/dXk3bFodhYw66Fj4q4WcZ6iR+Nx
yN62Pu9ED/XZ5Co3CqWYTM4vkTuKA7DzL5dv8px/dm453VQxBbgIxIz0Nj9E
QL01Kkj9cTFk8aPF29Z6Qrm96linoiNw/6Lp77Wxqwzo9nQ+s9AocB5t6Shi
Ja5HjR7IDuv8uD1KBibhU5v0Wu9yzQhhn5uB12ZXKnvizt3pqg7upnPJ6myV
39EWtssG1Ag2esdBcMQiQlf2XKK2+QWDGEQxrf9mq1+7JRh4Iuo7Krx0jyKC
Ev1MEUdOXPMJHeH/uCXePpbEU67UUMQm3Pd0APk51o3Jcnn2R7UESNyDif0q
OhrxA7wAg5Tj+jYEBW5qI4NLUBO3rEKbYQOrlICCKVvgXXFTXxhCNQ7CJN+L
ooDy2JnnimpxxRfiDJ+gBo9mXnUB244TZezXo8IEpWBN6FmNjzdAK5p8cpWO
BSRwTTzEoHwBxvG2SypWbhBYxbmEggl/2fgpGMpC5QFzTFjpUFUa8XckIp09
GLgvFe9GByTbMXqo+zISlbYx3yEbK9Od/6WJc+VEuiocQUJBa5MhwZZ+/88w
DLDFMvXx0H8NsDelV53l2OX/brMD/9/UTGu9xlamS/w22pVUO21VAzGNSw34
eXsrBqfWRud2q88WzOLNpgkkjdqh4AIPjGHjBO+jB92UcKxvYMxRHuTULT9s
4SdT+TCks3lk5nDcXUiPZigTVuPsLRFSPHKD5GAULw4dQk4ZHd8/0IqDXDNP
Ld5arkD79TCNhtxJi7z/e5XW8T5eYU0i/Vf4Im85V1kFASlfQxzgNQNvHefw
i1RpYdctZvyWEX6q7WLz4Ia97Yabpe/5UxFflTdX06slxW8gOHufH82bKMd1
fFnljf+y4jY/JG3kLXpWqAMvYdish2i1zOBuws+iH5chtS7tTD/6c6JSXSUD
IN/fXsyprKOt1hHtLLiCJoRUzY2B8P9qUxz7DiKII2P+cntxPEWzeDjwwnI3
DtO9a13mjJXF+PksvlX8fzrtTVdNpoAhuCPrz3RYlyOVRABCUsGhXY+9h4Au
Q8+R1jmjoK/ZspSpYLXPlH6mnaZCCgpD3T17lxYMAqq2qhW+JbOheboZw0wc
iF7EEVMYzUw95jl+kTXYzoSGK5w7FOs/RrN3q7UzYLNmoZyas54JnWnlYru+
MMM6ffjlDiw518kdNyANobiKD9Ir5qs6v2rtV3zKHl7U6xDav3J63QbG5mjT
bieh3ck6AVh2RswZrhTNnROFR25rQMAlbGuj3uuOOPCyvTHlSS03V/9PjuUV
bymisFfuAb+ElyZvDNaVbdvwzvlBby1utERgbzMuX10nNLk9Viynadx8f+8R
7aKZ54Kcs0KOB6687yaemASegCgs6Tu94T+6wvI0GhckKZ+J5aFHU2/abEf+
/2xK2Ogifa+KIkHT+JTyCsCFqY+xoTjPZlez2d3XN1LXNh5auYnk9nGCd+9N
HLgmr7SaGnFWCxnUI5QbcDKEuVAfeLEM0TVSVqihOh1WxBhXbY4oN9G6kZms
dQ7+Kk/v3a1+3CtoouGHax4n1FQU6KKFQrgRXJxLBoBr8ZXF+jzzF50YsPdB
qCJuuXqlfSReq503ugMEEHqR7rz2JYsL3RNqtdHE8iavwPUpFUHanFpWmBxq
n7osgAsNEKZM+73lFvDjZDulSDXmGkaBdCec03l9alEu99Ic/dbyGcurMVzE
e4KLvOE9KnK6EAksQSLDFQ5TTeipzMh+EnldQbx30xFoLLXdCveFm0u07Gdm
842wvC9HRplVlTAfwTfPxXpvek56clkXFixi/3lfDOLsbZRiUwaGB260kwK+
Qe36VqODP6wAeM6UuqlZUPJ2esHA+270mHb2ZHCddp+Zgozc2EJYMMNJoqEZ
8gKyMENFjmPN2faeb3UhAbvcud5gvfaS6cUM9tYXGY7wX7u/T7rB9x0TSIfa
GvubE2UA6QJWVjSc7uJVbqABmlMHfP6hxX2txtC03QFGmr4SBZlTgZnWTV97
vSWmp2hpiIXRk6cM98hOwfLKP6+2b8be+5ieG8LnV3lqjNMwyL69H4a5mFxf
1DV+1G/+KdOBKlr8Ed3Nx8+ADwWH8xX0/pUf/KdpKraSKHWsw52fXq4YrIUr
5DVQ8/zt0lvXbIHcNMOCfdSZD4xvpPpWDOdiH+2iJ73Ay2skugdF+YdVYfhQ
O/v+wjFedQpyAiGrqHy7xRWYPWj1p2wRc3Ls+xBX4YLi1sEE8w4/XnzxUbuO
DXQoKXArFN6WqhXHJdI6knHlxxO9R0TD8+5KZLVk2o1uAxh+dJbBFwk/x/TU
hJvESQ3kWtC+yM8PItw2UrZZGkXEAKOTqlqd31lVVPtWXappN7QhSPpS/B4E
LAQaUU11TTaBJBXUY9M42G/m3OF4+UcGpPfT0uNM/YkOteFPDynnhwWcqrJC
7+guZNfiBKPYp8O/M18gNu8Nt0/9zAvVMfFHQUy1k+IXT/FMvYzni9GBqMqa
4mVJ+y8j6cy7xq+P3ISAAX+lUADDLPA+UojPEl7uSGzB54HTlI/fFaUwDSEK
sm+1ZPXTE1yX6wdusN1Xo2s5dmDIAwFq+Tb172RMOIM0V6EA+H/77LGCVW7q
jhl5qbGGicLGYD6GGeNoY9FOp0QlGbxSq9dUkpKF47ZYPHwA/uohErETXLwF
HgrO3ogm5i6rXPDlamk32s1tfg4rjoQ3mFvxZhoz6VGqSAPKA1lABtxk4zBs
IcO4lBFeldusYnFKR61igs3Pm+b2OHcqrU5ROZW0W5Hdrh4V7UihT+azJyIv
Z0WEsn8fA/DeVjTT3N9tv1qkQuDHLe0ecPxOt+qni0dFlg4FHb1n6L08/Pny
3QW3rijx19VrIhcnndQMCm6wJXCmpUzWOESDr/FkZaW7q7CanEitVdeDU326
i7itKeU5D/UbYxjkcJczTdrAh0yBSe4B+bGHQ2YxGhU7DFv8XyrucBjxcsjv
/ACch1M3dTE0g9aAnam8kZEYrop14G6NYu0rhR1Jy7PahJzW8P5g41AGw50E
IEK+VZyVMo+8cxa19r1AmWZtfbnnJegkM+YWsE5kULBpjzg1UDhFS1Jlg1Mx
ZWhs/QhBtpR3xTrELEmtk/52oDlWLgPXGsIBv2B6s/2cphqO4gkSgdnpHv5Z
VuY+GkUkU0Df85WDKojktU8wWV4X2UXvWIbyAZSuYfrJwzg779r3Yr874FVS
Ht5iuyZM8d7BVd1ul0ao0vY2UtonGq8hci8nyMzioIEohjlCxcR4u5BvfsLr
Klum7ipH/nYmHFN+BU0XsOZ2P11kSXPMARkWq5z3RRKc37SOCtj6GsOrNIVY
iynPOOhTUSP+jeQKVYnkK4sQ6gEjWQRSmt/74hCjWEVWCLNAEheF+C66QwK1
MlPzFiJxALFlPZnxmoQTrDLwyWF3OJ7qaAB/ozjpo2mAqCWmqWmaQrl9XTh6
AKTGNM5EpQ5xBVAzJQbF3MmottX3f4HdK1ZlZXCH/a0jLecPWulgLpREE5dp
/YgPJtiwPJiQZe1eQdNE3ekPRoktdN18HARry5yXhcDMmpe1XEKT14ZOXoo4
lMwEh0atCiLcaCRUj79e/2X7WFS6/k6Ro6ySqaWP5kWWgiaiYjrXimqV9JIl
RlefINhh7GFGk42pQkfOFwYhMgfXVWkFt0QYDN8f1br/OG3mAGDZbYSzyuxL
pEuEwSZni+DG66lzVCA55Iw/SarVLNfaN7mJNPcQRf/rg4TwkSqVYa9nC/gW
GfYWgQ1cPhrYVKEM1I1oAoOvGbohO2U/kbfNQ8ZCRw/7hdptgO6149AoFEZz
YhuJCiwTTXNH0t5WKtpC/NKlyJAZvnz58QngeQsSDGDBE4QtGiLLH3bh3lDw
T7JoTHil4CuHZ3tlFjZ4syfydGUtz7MzYYtL5nSCPLgG8pX/vvpheK5ETicp
uenIUWH0D2NNtpQkJZ9rDgaC7LRC/po3h998i3nSz+aKtqfRGXmPJcz65wUc
2573/UZN9zCPokniLub0qRiHASxeLQZVownBUeo7MSv2ug6gY2btGliSVYJo
0ayo7EP9oc4cynhqzF4WBEaBlP2UMOK4udpE6lkabwCoiBttRa5t/b+5RmB+
ONIQ3laIpu7JX61Xr7yiTPFQbWA8rO8mWsn0xiNCW+QKz8cphkTcoUtX1Cbt
lRmLL6vdl2V470mI5As7RcUpKKi5weLCJRidqRj3hv90QPwfVfukzOBqkp2q
Vn51iuE+XAj0vjdG3nt8ACVDdoqtJIaeKfAsr6fhvFoC4Hu9FzPZ1U8a2tBe
bRQzjfrzeihcY/RzrfjFRQkB+fFmpLwC6SQSQn3rzrGNXLsqgJwa/O5+3aYp
KFootSipqvOSgfwnS95bF3MnXqwpC3x5N9mul9z/tmOrkHogwgEtO9UZT+m1
hBW966XTg3K+sxVRr+DzATYwIFTTfjCJD0H//7EIIN0dK91XEwZxwWJWa5Lh
HWckYKAsL0meF6OvKL0lqWSf03xonS4V3cLNz+0Q+50zB+qNGvf8OnVbt1Gv
TE1GNNPYYVU3uKiSbfaCJFuz3HEreU8j4KN5GlJD1PTDof8xgiPLsGZJwfCs
T+zR78IWzaMHNYRGfjbjLCuAtQ4X5dZFhUsYPTNL38rckczjdHb7TSDcrzbK
q0kZZmUuuJs63eKfN59OrWb3jv63ymOFO3Uayd52fys+8JaWamqF716hXNch
wZmyAVq0Z8dwCN7SfcrxrRaDzD1DJzTBvR8p5lGNfDodl3EYouQVnxkgVjjl
+MCR/WmuFXrgDE0dH7sqEfaS/X3QS3ngVPVl654+aJASlO3Ioy6mNUR+U5xX
z+T8aDjI5BTsqbKahJnWvwJgdSsSMhWbfEgfNP8gl96SpcXAVqmGz/HnLbbf
e+mEHqw0kDQ+kaxVLHDiOLBXNgBE0C2JsOy/ejw4bSDu1JhGavZRll5V6phA
jBT12hMk7mxmvMFPcmdsZ7iYy3tgPR8LsjpUHVfrQPh+v3GfHbGb9IM2AhF7
Ll7GzjvaWxDnvZk8rQDCMoAteS+tBStuz1dHpBce9UDwHBe+DSqsrGhfqrNU
XMty0jZl5U9wZF7hkwVLkvOpCzqmKdLsNpo+G5vP2vTVigAgrEds5ygokAsj
R/5P/x4yxyKdC9a9ZdexzwW3J/oJT1CIuuTcTwT2V+DbbImw8xHcKje31CPa
N4ppkH8LHs9rJzTtVN2FRxotlYXC3Zkh8cIjhftDlSYay6kzRmK7aXxq45i2
ibEE5/hMNfPSIUNzUamsNqr/CspZyRm1WzB9GI03vpWfp+VJXzT80Vgtqqla
zzdjieqjhPmLmmsm9J8p+yXHzG4vHpsfpLaYwjh2S6+uGH5bOhLweN5qvWAR
fvwts6iO2pT3YBK+FGT7LlP+JfNXVcjQk+Wgz7bqP5u9snKOUxf4T4WefDQH
aQqdnbkq+v0P0Sb1Jucyk52FpxUcChqoDrvRlA6MnQRJVODZ2sEZl2IXwXXz
Ji510/+WTy8XhekvKOaBTCIQX8RbncfmVH/F/8XYL9ctwu4Ts4eOSoGVCYx2
zsvAKYFOAt5qV1JlqruGE/VmKkdlFamMLgJEhbULffipW/Q6qomMSoP6qo0T
be6VCKMnurT+jdPlVFy+fkHI84O56739ZPmF/VfVNnPo4HegWPk9+Lln+atz
sp0qYadrKbXVpV0GYBloz+oQActCsFx2c1l3LQXDht8FKAXgR3A7+YbUU+LW
1yUJZIC53zx9D4udlsHNvwmLk05xueOtlqoHeHAvwWX3yqXgxnd5kmFjquU4
CXdsM3S4v0vCmUOBTslzyCR5EndJOxhlZQ6/MXo92wg5qCfPy+I02WhA6hW9
CZ0Z8/cDGbvqcNrx4pz1X2sMtxveKEIAmEHqG627NqY3h2CNEuANw8LrJIc6
dZww4tiDlZjVgQgIYqFPp5o/RQCeg+IQ5+BKG9sKUJFuoqalerYT9n8A7zOP
JfxWMn0VI62FQ9kZGytCxMyj2Pz9ljkfy5tkeRBRbpgmhV+3s5HAbFaI8fbo
7Mpp6AiB5SqtZV3doTFba5qkw10teZ8Pmc3yZa+yEsoVJroMUJ2Mt4U+zU0v
RbeDJ9sI8vKFRqXrX4v3T1KTRRRsNv9kHwAr08TAsJKneq5Y/qTyGDLUOWZR
Hl1MqbK07ZljAONyNq3nQqOAJdA6n0NH0i7mb+qmgVWRtRQPWvtROsQ1Hziw
nB0/EkDbirA0ROxKCCF8O3cVLUwoPJqZK5s1MzybMdnuLV3ZZ+2Hzv2RqaCj
FIIjubBuoV0th1Dsn3b0GNpas73JXSweO3jV/X4ZrVq1SHv2XTsi+ogMGEcp
PBKKbZv9xLrf+zv99+B4lpBQ3wFb3YkDhbaVMKUcEs7Mmqkj415nqDy/JrGb
MtJPXzhgh+UmuZHK3sTWxpaB1Bad8DLThKrRK8TgrErzgL3KyY1rgR+kXno9
9wug1vsUwGsksG0Ht7Lp2R5a3995541LBb34Xx4jaVTeqJmmbykpsAR+nFzp
SFIvJDd7q0dnYWTGvF5tmuJyqDpdwEbhs6p/p2Tx77d/m7E+haZwAQIIWvI7
UDCqyFIrbnzF3FC9syPk3rXLrIGbSFvO3MMJqOxgLgQP0IiiCpoi+CTzjaQk
GwNHTDxECjCl51ZTJEMeAnjU/FvwFPTThk1rLrxDivxGl/nK14oXQ19fwRpm
oleJ87jMLm+xGzk8hy9bV4aqRx3ac+XulzGp9msiyj+L8O7GP0ChAqwj51Wd
jmkj1NMMYMiWUNXq/ezxTOzyjj+8kjl3FcuJ7ZH0Pyj0zSNwYsn4DQRe5M7O
LMYK8htf/s6oen7GpsYuj2mvVLiSRE/f/d6pqekmCcVspQRK8KqG891wIYHL
NGIq2/2S2723L+/tAbPnYCtHKdE5IerX9IAAAS1Bk3qU4s0flgpzV7+EP0yx
BBx/icyEJtQuBR8MJ12RaEk0dmtCLynaZgcnskKbGel08jQbgtsptEAFWrm5
ZrlWDujtIqoKrEviH9zOMZmVlsrFZJ10/3937JOQe6cZqkSMAES4MdHWzs7D
vgbUi7o1MM3x+jv1KBmE2+QGUThn9fdAhdoTFt5rG1zbtjjrp0cGqPA/ZV+p
EPbqp0jDSH13hQt1HlB+ohVv8KOGrekwKVJgLk17Wq7i0+/hyT4NtgGQEBF9
rNYVIIKtMBIIvisZurBzCmpFSk3bHpcZW1G3yegH62r4CeeZPZRL7EgRpwrN
mP8eieACo8C+4DfrSN/buwPQ6y2X2iUNmprEBTWpONefUirAxgqkhnMXEgEZ
biLR5u4AMLH3p5u+B8h3RH7EvZsV8J08GpuXXKlGTYgfRCsIglVlIBh3oi14
Ge+Gp3spvn/l7mIE38FhzMx/ayDEXlhovMgG0hh4RWRokQJWOn856/3j5IVo
ToZD6mTR8JNzLuWYJATm5J5IIswgjUyo0odyOczzIUybx0r5lUfYm2wXuJBf
/MVInQkWk9zI+vOIby7/pVyxk3Mooth/Rclgy83uPBf/SYjhWvhlyVqRaPfA
jZfWBfTtwVK/olkCT512rncu1KmjNqIuFgGfL4AMOEayqeFccB1/3dWafirv
awUA7S6rBi+67E801eqTHUEU9+2qUAZM0646WCf/egQnznWpiKfbjk5XMg36
yWVi7jkvv8Z+qB1bt+1EEf8Eq4ZZsE8P9s9hyl6wpBKSso5dYUY+YPXmEZr3
xyqjZJKeulLdMaSxxEwvmTqjg7dSf/VAaEL+xYxPw5a4OSYVJyyRezXDuX7+
Q+lgg2EdFn8DkMcHJK/ZuGqkTvdjZ93fvZBTL0HBKLgmX+juMM6xoA9ErV8F
NzHsMQM46GEIFhhz8c0esz2LDQBUyKBWqjXroqAe2Mwfr9fE38rcAvCqUoFh
2DOqRk7lbOSv95luPh72O4E7pBHSc+Crtfey1hdRFkoMOl4DW6XCzmMP0iz7
qAjrOH5p10/KyMe0eOnpAfH2dNqdCsxRhhYGPURFOPh7mXkoNNxkMpO51uNj
9Xp7zrKFQLRjt0AJCm67IW7YuzARbk/Ix4PJihEPTnr7t1W4wWgKwxRsBA3k
/dPUtpbxNVd3w5wajrZp25tt3LCsL23bqnZJFXo0uXIjpzG7qyunAtHx86d7
2t3s9ttmOnQ1VJZub870s+hdp+ToD8zE+7LIJI+/RRSp3D8XMBn7qM7M5YsB
DNUf0g9fJXM7o3YQX2mT+5wJr5/w0HvGp/kgTcMZgaNQjNAzcmhm6kyQ5khW
fSUNs6XRaUV+peAA04S5g8A/9KdsHW0BLV60gig9ri9RNdEC8KavkWSCobGc
DRV7MA+Qq18nCAyNaskGPFVz9taZE9ESQrGTJkVZTfpS0SIdkid2AO+d6nFq
DfLDqnZc3mYTgsyWJUrIdR8bCmo8+sB5MH/EeHVwYE8dpgNVn6p2oWjr1LKh
kWtfXkoFN86EP2TPZFq1Fc8/43wfvqqaakokfck8Ciy6nDQKxR/f2OnbzZC8
qBW5I7bPFnrp4Z1NkOBwTkju2QG/hRU51U03BWxYpTpsXw2q/jry4m70g5vJ
u3uL6wjBzC6vZgYrktSVIUMO6nR0pYgHfKolTtRtlH7tAy72kSbdJJsVMVSo
R2segbtGss2HuO3kj99Iw/slLbExQr6d88z6EcG3lrU7U+uW9541VBxht/Yf
WkX980Me8R9tJgDCFG8MG0PQq9mZqI78BxlfRcV4PUrglo4C2D2GiE2FvZA7
JHa7O/ocIWAebFm8lUI3UuU6mIIppzjqNdvoWE4NygRSTlsO5yWmOlGkXYfW
vBGeFGcC8zdaoteWFaqWSaFprXfoe/Wjf4NjC4cyKAG5zp5EA3qg7W0rRDMD
dx5IM8HpisHGoCjZtT4ZuR2cwo+3EWIBcQrGpFS/wq7SV7nnHLwQjkhpkCwU
z3SLHEEmjDTlA7eOiadch4S2YaZ9tEexZGljsK6m8h2BiE+ve2mDD6YTnqZY
wReBe1pxytC2GVFSDuLkdZ5vzCSrtVXKU5jZgKAVIDuIbL2Ic6m/mMJEjrq4
Jx8V7vsKs1fShDTwDX09t1BF22Pj1h/pWazoKegEt8mX6zpPZGWqgIq5lNQR
FJ8SpbO7pbmJVy7pEfr67+EbaSuEo+abaZ45j17TWJSOHEzOd+wMwyMsmfpp
fslBtEmNlnj9j1nIhsNsPewpfNYFvBJf1FxmJCO4T9pcKBWpiPoJJZ0cwfUa
hlcu2MV8gQV9Sj8bEdDjK0B6z8y5PMQHhCho1FUsRhf5l1fQj+j3iYLafAtA
Nsr1v9eppBmmpvVD98cnWDdhV+und110tcjTxgMsZ/1grAHDtGq+dE1Hp0Sf
CD2lSR6o1++4V5RfJH0OW1qHtpNWwNYgoBCMhlup5QP+z+v49/ramr2kJ3aU
tK/POXQyg2dK4B6K8+Yr1S3QehxfQG7SaZz3F+ZTPyroeoPUnSPZvHw6bsr5
YEewGny8UmvCbI0YZvhG96i5Hwsm55gcFBdRAUeGIrPwUzY9ia7zUVteC3mH
bA2LKv+VB6iUiBVeKPASgGBEKGeuG8Y8aYX8HYDSk3GfWX9ix9/cRdTIaOer
6fnoceEBzRVaY+vO+Kb1BcHE0Dm5yO1Z4MiiRJbVjKnNbxmCHG5blrauCASA
6XqCjMPivKNyC2T7wIIkMkwvng5M4monfpvwNnDUkmHwdO0VtM/GzMzlhqZ8
fk4fe0Kvd8gShJR09RAgHACKU3lzu5rbLYPwgQrvAwZsSIPJTqhcXNnr/d49
LfTwvgH2uXwXaw9R/BOMhFGKTtFNyxwmswgXXiC7YI/Cm+s6BIfL5PWJdHwI
mKfWFWWtR2oGV4DHbA9R5Np2CfGapfAAmxclvuMLj1TaFrbrFH8mvr976JlX
kiDnKWBvNQZzaHvnJ5j/uB2kYBL+W5zbj0u0iSIv5etZQGxcEoiSbUqMrjqQ
D/ikI3XfY0oncy0g3osBkXRjtH9N15IJ/ZozalOPLiVc72zHR0YQBmLnG2xW
xauD7XhZqP9Zg5u0pymQlQ9F0Hbboyeu+rZKCtqK2YMuW0qNThUiyAldRcbA
ugHsT8Ci4mjkMKOVpalzS9AksE9ycdJM4NvPfSDCFYR4anSkvWgAyoHbCemH
pbf81RldFK7gMwd+Capyy8ySzkNOIHQIwik/knwhNyY0dTMRblanvxD84psd
DsKsOxOh2060kG4eNBAZaaqevpdZBnGoFJED7u+Ip8kGsBJ0QBDwS5WYXaO8
CeB4fm6SOCjzcjm3J3QnOpLsnjn1qjqjv63cAktGuTdFdBYklZl6PEhtEivA
OslbO5WHBzHLTjN4VuSAoagqUDuxCxkfip56/Y32SzB4t0Z6WyC8qc9VisZa
9EHfewE6VR5YX7jWT8fJXzYlD65c4v2ljyrpqckX0S2HdH4g+WFKIdh1XTZz
P/BZcVkLtBL+e4EvzGrj0MkBG7fdbmrXSq+xfjgsWxj49L2DcjwBsgeDRg60
hTwwf3ycrKaPZgiFZcief08Q7LDkoGeualR7BvNpv+u9FUaTxMg32ayP0HR+
ZSUOs8A4lRD5yFETEfZ1mL1AD4jCXWwM3rWHm3lVBgYF/yvxn8GbaZKh9GLA
YCEn2wBHRD0Kr60HbA0ydSvrhK0qM9rThrO4l/jdb3bNq0yt5lvfoutnqllg
jNuLgdIefj/47uolIN4Oko7CSe/WlAc8uEKEN8iIXX91Tw5eDjl5UIJ41VNA
RDTvWS617yvbAniXb6PxaMQtgNVV1es/wENTFqIRIA8wI/lDAUGxMWTK4kQy
W1e/Hsgjfuap9jNOtC1TFxqtNBG5VRRZ1PpZCw08+0zvQNuWmZia+524VEUG
4gkb1pRn/9deiHC38iFzA/PvAc8eYGa4Mc0z6Bxs9CAYYt7aVRmIcvd15lHn
5J9aBIZTlQKwWcEumPpXIMpQTSfuhqds/LkIMCsAjDGvbq/0pD2sxm0TPYr0
oNi/Alqf8NqG3I97BeBzGKWdGJPQYKI0rfsO+cm41bAvDDFFlpVsYjhxiD3K
WVbdppdP/uwEjf3YFmqK9FFXIl6Tend4KGBeE6rpvxaEzk5E85CVpWZEiuZr
VoVUcjG73Js9KaEM1jAstHyNlV37SxEEEmeMAgTVytygcOOkpzdmmsbX4hyt
CxUcbo23tVcKq9vGvIUXSk7YddBXxtolVJGwILIJBjohRZhpIzrvFNZV+3h6
D3Pu8n6EYSvEHBm0bX/HwZg6iqpB1bzR3DSbhjD4nWH/fJEyOimYnTcq+8Uu
kRqOhx3T6lFiGMC9y0t6ojcfKCzpEnQ6m3jHORn3c2hxHNLOh+7qb0ePmPJ6
Og4cwcdkAid8PXXlP5X8DRhXsMVc5+XayuQVwjolImqvmhKjxPkDxCrq9IaJ
BImHXw+62tKkVHEoFT91/UDslfM6s9oYCkNxifywIXoSw/cOgZKgyHZCN+PZ
VBlfInV7VgopKoTU1GxjKHY0V+9rbfoOCvGzjjUqq6Fl5uY/aeMLL+bAbUvG
1xmVme3HgXtxc1bF/XzRuDiKk5X4HVakdP4HtFSi2GC5QyCTeViamzOon+qM
ENOWQkV16DxGIS3830WPRqZgvjzxijIeoT6Ox8X2BlTmke6J14Z+n98dkUCD
kcJj3MbZkIbTUgGzCxstKkvqtURK/DeSPESERRtOVS7kv6mszHVMsqVxzJkJ
W+oAzwNj0qdrzQtyDJNx8GzBd/ONgjmMnFVbeloNW67HiGWp0qW4cxUgd/yz
X/Wudje9SShSi8K7xZXKPF6UQAbz0i73S5COmyKm0M1xjWIK9V/nKd+JAGxM
jzCnkJUa2z02ZtPnI70eKyTEleixBDWw3QTFzLj8dpqepEuqVbWWsoNzYbBQ
hG4i3ERaLwQGMa+CEtjih5zBdbn9Lde5GUqTjMfEYBcPc04Kt1Y2hn7t1Plo
rW65RChGrN3O79daNou5JOJpRbVRj+3hiqkd3ouOOzVM8BDLtwpTyTuQoPNe
EJ2jO+trxZ5wG+KagUHvUh7LWy5FnXbbUkkTnC9bnbdlcu1hnSHSEI5Ku+mt
+89vlWlnbyk/PGXBSL69TtdBHJZJgiRW7YxcYZkK1HA2YDHQ+6o/6mk9PGkK
/gjpKEVsvkrtXL/rA40BTjEvDXrZEbvDe5YABH21XqtxZ6NWRSuLjCOOSS3p
NzhwaexjxZ3A220Tv7ev6O+BBjmJvGOBLYJJkS/OYnKPD23iNWZUjVK1Wshd
0x5UNkv7J1SABL5K1WGpCQbK7eFr/IYGpu1KKcrSzBtUTRJ0B/cS9H9vMeK8
eIkVsMJ+8MMxu4mkCvMyKddinWmXAPQboAgRr7LXvm3Gx6ZdOBCFeUOLTGkc
AXOVR46vTZRf3Cb4Y52ZOLyJ2mb6hwBVb3nz7h5SXrPMQj3x74T4wnkcstJY
GyPFvLcHh8BQd8EySnr62zXmZoyp/399qVS6Ko/CsPt8YeLIEMoxGjupwUFl
lv6B3dlrHsrzC8ekh1tFIIDDFoIsww54rnfPAieXkVQyQjjkfwS1GrHioLmO
1+p2HwoIt/3j6bVXG4M2O6mvVV7X7CuSHpIw67T1hyM0B43BpI0Vuwo6mqf2
uRk4+KsKBhwiNmLZKKdNeqwg0hUVzTqQUEhb6CUQAHwPNnEcn3zpM7g8y50u
+hgR7UqMNu9W7XZkTgmMD3/sXFFgHFmoi25iQVSH5y/FsbTi3RfawGhcE07+
7qN55v0Atjo7JhqOwdxovrHyaAvxlS7b9tXZyQJnnZ6YDy/AoAVnvb71cfA8
TI4BoSAHsaFtlSS6PY/g4/pJ6BPAf46lKD6dO+WgFU3xvXTGCtH8KI4vzX+q
X8CZMAUTLntXcfxQzflT1nKzB3Hizyj/bW8IIjiOQUEN4maNgHk2/8U5rDwv
v5KbYHDqgHsdNi1nLfM2jkT4uRfquBvjD+144Y3gyV/oGtCbcDRq0j0b+aIg
sPf+LvCJIn1AOuPNaAE29OZMQJbjSI+AMucq41Haj/aBsjxdidjRmdSEwZx7
fIN42nE/tCgIyUUf4M489VKDlV0UsHVRKKYV19SfYP8CR853gWd0UK+Pf/Uj
MxKUZAzaQUQ2+/BjHSTptsHZwFA62MxooriHl1x5dlxr60NjLkQ8L3r7tiv3
36A22j0Q8arJ0SB75mH2ceZ/COWsVg7hU1v9ukcHm4ofD7qJ9BopZ9fvl+S8
sVikY0G99KSQZeUOyogBQyXHHBRpWQnGeJx5eXgt4XPgXPPKs3BRDHsYmqyC
ZRfVVm3+AEySxPgYUdTns2z/1SRYdsPNJiqzdtAqBKJNSFt15NNTOMQhYt1t
FMNlGpUnaysJJxxECU8Y64qlAuw3rr/oQirgZ4guaLPvDtianxTJCX05plPx
VLMym2cbLez2t9kVawulrh3CocsgT8eqCFGNhCAaATdy3qO+PFA55rLvdAYx
Tl9GlykICKDWZgPGEK0CF3oMIgNWYL0qZzB0LGL02OCafhnyqWIO8FrxBJWM
hqIXzXh/O2ljL5zlxitaeSlJ3L4aQE/ajGj1rM1ACV69BUVWSa4uOkIVFKcG
SyVXeARcxWJta3hJim3gvZDmq/wgsufOuDCZesRvld9emDHo5YaYsLEJigC6
tU8Q7fWuIpGNbb4RURkxgP6pjSBd2Avbnmk6p0P8XcWzNAkR1tlihyKoZcrl
pe/W2pRHyUJCJ4pFO3KpVoM8G5wsdHEqHTiotWfTFL5YaReD55LQeJSsTAWn
xzxet++rL0zfbwIOhtrOvsIEkrp2tpky1BkOrPSWLf3+MSLm7AfX3crBr0Il
CgDkB5Y0SwpGjSq6dAOYvjSBFN9ahY/xZE8ZeL0L9FGpI0dm0Gk6PWSwkMTA
3Lpena+qi+eG77DExuXafnjMMU++CMsleWHg6eD8Niw0Es1e1I8hY3h+mNhV
bNCxN1acLKkIIO0lwqnG9qfyzDoIt6Wdc1JWpEXdbjkyBvexJjGmKXfOrkZn
ODmqa0q8EWtMGLpz1quSYd5wIBeUzpQ5qKw7qd1TMTK6II4eap0jCq8Akib9
WTmTya/6RRTQQhSEQwz+bLLfKIJVODrnRC4aJlYbS6kVPEpa9fSNiWc1GIV8
o3slSuq4YdAPw9ytRqLa2IvChFE+nkf6uqK2R1bFkuIyRYH0GYvodfds8zFH
bTR2UrW1c9XYrwUUVIiYAXD2mJdj5U3QjEyo56tYMzwKqkGryzGi/E1vE0CA
s7MhhVbYkZJmA7WK8MuapdR3ZOH2lBmlij2/WKdkAGURUVfSBxMj56ggE69L
lZZA8RAm6MEqyGxVw0UU5CMK5T/7W9cw1YHGSAoYLNVctnKP8b/iXmfdvFx7
43MMC1kI0UBD0KE8133UF6BRDoK/DcAT3cXz+h5n3fyvKZh2Yn6Io8capGvW
6Zreh0mFkA/dzYuzHUULDLRZkN5qMaxbHQaodPxwwPXG9hv3SoERIO1RI9Ss
hf45Wq/aTZwFFwhHu1OUnBHe31T1i39YwpTeu4931uACu4QvBesNYgPzjUDD
k90PyEAbuPaZZpymmVZvU47eZ3CD6NO7/fNcnuUNx8ag9+Nn4Dwmf/Fr7eQE
59QcZhssM+IRQdRjBPBWSUUAfP+HVxWBjoe2UslXI+i18JqnmorI/A4gl3ju
0NEFJUSid1Ondgb4xb2ujdgCNdrObFXuJyVDjtifmFCApMK7xq/PVs01zH5b
Mfr5l+CvcYVedsIuKpEGJE2flxlllNAWTMvBw7GgSLMIwTu8M/mfFk7msp/2
jFQVvG3pb/fIJpmqHSYeivdBFv/aCy3K57ffMVuuZi1hB/Q74isJEt5UJUCN
nzLc88QXmyLVb2A+zf7fckd1MKF/XqV0Vk5+9znlDRLle6f6SgG3jHrmZ/kN
5zZ+EQd5/4GnY1b9RmEblEEWwfUDYUb+64MP2xsA8A9JxV8T5fXNc3xXoeM6
G8VUMPbs6F+MVjTnwISTHVQMDIIERZLlXd/Mj5z5dKUciXO5sHYvpcu+1Db6
qDULZOq7AZVJQEO4q9zTJE0b88ubBVBjXJ59I6dyHY6X2GBuDEYsVZTHq/3V
/mMnoaVWBiFTV9aptVwCXa3Tq7uzNtN9Ww0/RqHpxIRU14qk3moHCDhMlyW+
vQjygIGQVpTuVGIcV/ce9U6be04FXiPsH2l0cxPKBhwh8VEK8D5/eZAB+och
yHQV89738vQxxV89uh/frCiz47YQ61HhXT1IN4P5CsamgDH19NxXwyQ0P0jn
yfj3hBU/pavKNLrpwP+w/iXW4aSVijmpL6oH9zIiDrjrETZbA7SQG186M/fP
7rXWgnBazuFUYmpeLC9UjEpSzoKewuztjG5HYGuTc/u7Wou4DtDuhr/cWaIZ
rOiCosljP2KNZmUUNGFbrF7SRC2I6N+A7VWhS/UVUwhlcYno9G9/Ba5DlwLr
8RsvN0xgbbqH/U6IRHQGvahH+q0BBOjbpWYMVxdYx1zb4uaV3izBkzzHvbCx
hFgECPYBhMC62zeLYsGrlw1bYiKPPdjh/+qgXtdFnm6OJo6tadLVGmpP39jV
HwfJrGnR3IiA485Yz8vW/KwTPzI7hYR/f8zhXF14goBxMaZQ3iRPXRWFdfFb
uRQnnJahhkQuA+y2c+rPFj2LqCAulZy5/3kI/yhJB+R5JrkXWnbOUtuNZjT1
Jm6SZKrAqEVVTjKS2o7pOuldTRmqXN52Db77qWjc5JmEmNZel/x8TwiLPjgO
+JmSjrgdMZY59o35hXsTwerXtxyQEE06UVTuh5pJ5mmnU2oDBEHUYDUijt9H
HNav0Lkry7cmypm2xKffJyEBdAdEtBXQZySa7MPCY/CKf/1Y4Ll3JVy586AI
rUbVNpz/o+FgpFJfFZqVCN8KXb/z3tTByHGRum7BUoNKqc2WwkR1v1QCUCqz
z4qKBScCnPGX7a6zuZr/fc6Z66m60zHMoUuJeviCoAAsDeNsGfVVqiF9dois
PtSEafdtNiNyhLNXs/jsj22kXEdlQ102M/FK81Paew3zMoqBL7z5ULb63Vg+
3gAuU9EBvMJId86upiVO1ooyd/aFpYjL7+mL6og/nXYjFfZldB/FHk/IxSfV
/QsiQkAJLExT9NF3mLQt887I3CRAaKF23nbVONe1eDmCGZA7SJF5lSITuySq
5j84adqz22rTfo5mDc83JHLKglBBKiGfr24BwwWrA3m2kOQuW2mVobFyAxp4
XKk4dBR3H+/Y+/QiJOyVOgH/Fq2L/E+SZdyC8gI1R1Yi2ml0Byo6X9zBaAja
MIyHMbiHFw645jhT0aImqBFK8iE6+Est+FHuOcqQ6ZMR9ePtW25lpXH2ig1P
Zgsq2TwZy7TUmRQSi2eUyQiNO587HMdbxFRGl1OHVrEnYPGfwouIUg6ive4f
awjKDYfrF5INKHMI5Q42xqD6k4TsyZWrV1KmeHTTz4W//6cu7bE6YZ4QBbus
Rm6Fxnv++qVn8k/Ty6nG6K7nWETQcxJWT1tdNVIoMekU8aKucOqxDaPZz5Ss
fTJPhxDxLNQ/7vwr/ywpsY9Lmkpn9ibnj3vzhTl9oiEl50R+6umR+zvJSWdU
8lgBnJLDAb2t9P5fOS5hAT8SZlF6wh9DK9F3JteJER0weNYQ3UjfM86OZP7N
mQQZFkt/WIbBWKOxzXPOTG96GK/bVIDBwHjF1ZEPl77OeHM28el7ZLkdau6G
U4+dGrhDK5pNjSEchyn0jOuoLwTeev/mWM9TasOpFooV0tLE/zbgUc6zc5Nn
L7HZGUrtzCgmaMVMird/1klWFUi6S3mW97bp/LiCOKxOJ7jobjQqB0B4GIgQ
ZNcqt/vPKmgPGmFjzHYDC2b4Sc+335y8Us2EgUGs37igpFbSNMoykVPZ1BC3
UCn266SYf0XM57942IlpwOD7znq6eks6MT24CDoajAKihJZ8PXFfDZXtac2D
7DFO5Eq80FjCc9ILLZpzxoYA9rpLsdHeEiQqRersnsiJv+inpySN4344SgkG
LAxVUP6HQEPC/gdNyVTESjkAj2gMYysyFK14jVEDJ5SeuJaotKgSnbH79kfj
rPQ52ZOsEbJvhvJHcjedvzWus8BPH4kCqQ6HCYjH9eJ4RFifu4WDrfUnkgOI
1w6uTRuDSTotoKYA7lwB5ikRWprliZaW0GDtnT8E0dTT6eGk9K/I2CowR/Oa
pWXzDI956ArnxnvOwLT5l0VzTDy+zK7F8HA+rqKxEWy/EZbZYSscogLl/Af/
EGvt/dIGXuu3Vo1ervWGEYTwDc99/WCoeBYQjt14Gbt5gkPP8FYsXfsLIUVN
aLT/TZYME8GirePKvHcLtFpa2Zyct/DDdyllyDdpT2NAWSqIuSQ6yD/PdH2o
TPPjP8ppGCIfMAkZO0wyxIU3TCw5S7aq9W45wlzT9qiCQX43MI1TNoa0ZSbb
s3ZYcSvio9t+Rc7BCKX/3c9XzstVqdvLE3w/nt26r1+0hrIZarN3G6D5wznX
HS7LwH+eO67wWrHERFN8UxqknokwraLI+8ViXfUPP7fViK1rybedb115t3e4
i2uzayDMOyufTkowsgt7JZuA//2lmRCY3E8GmcsJrtdxUDgoXfP9UXUMPIgE
0R8I8jMVPFSXGr/5XyWX5wMIAMmsmTaWVAbQLsZTO4o2e7IrSB06SqoPddUr
VZnF0ycVHY+rA94TPbTk1C1hci2q3LjvCENJhHzCEktufz8/8CEwaKXTrOeI
WPH6egAp4bHZ7zb+y9iCUfPPMbYVWqLiUOSywpu2MaAFw1wwXnfUqIgtpgds
YsOMSPvA1bXAbo22C10j7PaPE1SkZZLbwtuaKzu62AlgCblJbKQnJyo2Mex7
5lcN0X6HdiJxSFPIffWAJdP/z4NrkUd7FhGI+3Q8HqKif/6Bagyt7qgm+AVV
5S4U3xiV4JLuj3zNulnw1HAqq4KRX4pLfSWQu4Ssr6PcQweA4O5UM6aG0M+6
OJmeSnY1dKG1Po1bReXocAtNclIH39KuWezGri6X9NUZDH6SwNiPXvdiTKAg
68GMcaV9BfKgfDdhQA6UftNAdvgGyTAOQHxvf/VG6o8oiAFje1vHx7hWrkwa
O/y8TxTcL4vmXGFv68W9BKcAsbR1WQnbN1t4CgkVVMYtelUtwBQQWMqwJBpV
D7/M4E8t2xqJz7K8PLbFlVsTAwi/chYfkaRcFYZbCaY0K4y/LLZ8rDtSOqZ6
TksGp91UkQskdnel/g6/pBiaczSQgdEyoZFqdKZ1cYTlQb1yFkiRMUOQevqD
Pf0PaOUwwQWjEwGgoAXNHEauCQqjo53Tauj+8wx7u3sBwW2PMu1VVhDnHRH4
ybGszR6HHfugNLqLJatRBCBZ/tAIL8+9yAT2IeyurhVfEkpr/hTsTEixNEvt
cPCpzC8Fxeascw6GQyOgBb+e54aUv5Ur0NMR8a3lYdZjRbkAHvRCw/6RFR1h
2Y9hIzp4L9Ozm2VpZ5YzLxS+qgGtw8kyBqvXvS0G4h1I6ylWSbBZFEaqemKP
GVwHiYkvf4Es8QaWRz1JaNAojrinvbXEyTkjEtXvQ7Uy8P+NiUsCwya4VcET
7y7h/98MHamg4xs2GpRSHQ/zQrtTw/hXBBegpenmQT2j77/jMSQTpCS3QtD2
bS4JXNbGYtIxVWyEBEYo0vJ0dt8v/zsT6cOasg3QftuKcwNeJKoD6uQtZKFK
rrNI9RHi+HCizBRcjjImYxVBW0Htqkg5MK2SukyKSQt6RKwxk9bz4TwIBnqW
2nkXlxJfwOxZAWHKdCD4HWkv2+mXJfNGXx/+Vwlf+pO+eD18pGf8olnduKAl
DvjJVcGMOZPhmY2r2Z9887uS+5AJfMD8EngEnjKccOjq1jqmKTbkjfBFOwzS
twplHyyFC+HeZGgoYnlwQXBkjr+us1zsS09a3tHWSfmU2lWsgLtTj8Zzz9Ed
h5e1DZekP34eMjKRQ2d4K65axdGdEHczhbLB7jKoF3ZsA/TyFD+5Yez7poD/
aYnrkd7tuMIpXVZ0my5E57mpCBl+Ul6dnFnLQs6JBuLVIFsZLb6gNtnrwXKk
Gq7jV+p0lIyVyWqNGELWYrfiqNNDJjD9jaWDK8BErWtCO5jsm0MZ4NF9Nqge
IEgU6HCq1Fr71OoiBUxFZWiN4Rxoz1hoBD2e2YVzulw5UUmWFtE4n52m0DwW
fF+Mq+Ivj9Rq4s2e0o1v0XQCBkaT2XyGCJZrSBj5G7sg9X2aD4hvpkysGywe
8s5Oh4tRgMDlnxKbbsCbO1bwMGFxkTdFGHQnPvkwmMWnEp6vaNtHlotlTJXe
WGRW8mCPTvsuIo6W4zuxsd8jAGI5MZFpWcSdHC+ZTXbh+CcwZF3zc0KET078
2wBAeR06QkrJ2H14tI4B7lUHSnnm2zX1GlWbPGrtQ5ae1NO2BIdAX6BLqX7n
UyfJ881VfE6wf3ZwTAV4F1iY6Si2+JrQ8mx11aT9Q8dikYlHQdqOF8rHC2Rs
1ZlISmUPO8zjCvh/cvlzxMNB84s60ZabearWx0J+kIs91aAGI2D2YAupY/WE
XyKODmoOCtjiGH670nQQUOhLPS/Fqx3kNMy6OVceLuuJeIAnV6/r73qZNem+
uWr5h9TDSClr4/PjqjeJlRHxZiPNBDpKhFurafuBovCcWybJlhvaogxh22Bs
8fRWLNdNaVsDWZPK3EbGFPsrjrARUFncjzgdV8ZeR2/+/a+7n87zl2RSaMAH
rM34FFNgGo7t9Pltj3fRr4vcGU+8R3jw4rrPRCpwI9YK0bUEoQq1dmTYtGLE
U1p0ZwJ8Q/HpDauqM7qjEEfYGmKV4OfjLeSjeQv+sgBP0eb1CkfdiFvnsVus
VvsMD6q2o8h6JGEaUWEhq8oxJoat6NnYx43S/9MeVlpUYjCi/qQMcbBvkIfx
eEYQctYOlm8ZMK8d449lIHf0DGIfjMgTLiUsSQ/o7SVJFrKfUu7WfAtVRCLq
rxjeblzVElgyY0Ps7Ct1uFhAFbZ1AjMTw75GS2WzF0SOd5eCD8i3T97AtzVB
3VLlHzgAc5DM7wfqxON/cXCiwlRl3dm61QGw69/D2hqlWPmgONvwhl/SHjwb
jmloSP+f2hSASr6wSx8jdgzUPG+AwZksATsdHShZhdiSHtoXowfrs1uMsPfr
rQFOWZL24izZCvg4Hz0bmmHXnkO7gvIDBZxM5DYT7gFF/L1dresB3A0ReoKZ
i5KadFWAwfRo3/X6r6quN8rBDH5j6HKMud6JSNCqsAkSUNWN1kHcOmqoKM1p
kAj3IY/UHcLUmHniZX6p8hBqTBEMLS1Ypxl8g7YV5HfosTjlPlAPPqcvhGMy
qlBuwpz0uR8/g9FN61QQvEs0jx84zDySMU6lGtVdKSOR0QvCtyGfIzxl+cCH
opgjIsoqVo2c/MpFRCjmjJqsbNMI19DugSev6cVebEW2vGBgnsxAOtmhB6uv
vE3GKek3hF5EP1ZuqLPsA1JQGkPir0UslYTuF3A5N54nKk12Ok5GSfany+kv
oDgJiUuLW53/VupAz8oKB90zvPJxy3C7SdIaYo2lIEd2tJvTY3xm50RPxL+K
5ju4zNLv9Nvx2P+0kdknAGWF2vQfUMH9srENEtcYPoWfkbigUIWONxyo8AGQ
29SVIfhM18lLy/crek3oLF+A5sHBJ14g07X8EoO69L6z22ekkjUWeYxiafwN
za+YYUkqQzkRdA8IEHtK5vXPgMAPFpQDw8T0FId209XnMPKtYb1q1g5MOvm4
2HsLMGCaeuqj+0MJGLjogwrU3GL4yBBSQy+9191BQ8/r9JWWc2bDC4Mv9UwJ
QwGEa5+adqQPlwhJcQGG10PEArd/pmEyrBAVQXfUf077q5NVuJRlb9xi4Dnr
iNgm09xZE/YfVa9MzVfwq7QKcw5Wp1S0NcSNmyPj8K4u3bTxDCxvqudCw4Lv
1zGNhNAelPzwyUniUYPsV6z9ygfbM8m53VDHLB7Bg3J4eJtc08mutYC8tCZj
eB4JSPfmDBr72rjks3cpooAfy6HPxnaTMIvbBk4lVfoqZu4kyN2WmgKjwwl+
NF9TsZ2dZFQuyO9fdyxQHXfGkEQWkkUctO7Z9PykLEtzb6GtQFddslU3mlkU
T7JEamlF/36eDNPI3dCXKm9wW3vIqDh+XmmR4WhNn/dhkUF7oOQPklJPB9Lg
8cZpm4+xaVQFnc87ESyXAOb7Zm2kpl35FsZCBdinIy16K4R5pJ40Lzq/twmh
Vsf0wGYn0a4iKMAZXVg/uIoYHpsjwXX5L0VTwwW0lgX9y8UY78dYqATI5vqi
ho4hC5/oWOr6jBGmxdl8EAFX1TGF+EFbOQBg7Kz2JYDCTYOVEE+mmda9OfnB
o/LiHBmrdqlmWbcVL3zLfqbHUDingQjJyd9M5THzAyd4u03l4iSZ0iFDlnF3
qPw5pTboHuqzzfO5N8HEW61szwZkJmyB2npc3Cosre6qphcXxn0OF8z6MIS0
wvaq3rsRygSsc+tf95maamPjGoVb9GG6LyUlOfF9kLdSjdRxIVYnFN+U4y2r
jeL6zls8OV4XQHj2okApbILZz4LRpNXroMHrZ7BPDOssDjZGDiBg9RekYmYU
Go4hqlNGM1F34gIkJWvzXQImyXTLK7uOnUBBc1X+tTa+AE22QCE7yFoqQuib
DQSjhkdu+YU3gd8xRufGjzY10NYSv/hhEBYJ8+gqQpX0ft4QNMJ57koJvPVg
s0lIF+7H2hchofzvoPkImCYbYVifob4uiA59UF9CZf4nWlqzc9b0S3UniKBJ
vB4dJrLWKSFGh7zFSiz5iqJWwA2RrQJgcmLWcuZB60ToUwRyuaXQm+U4fUiL
1PIxUPlUyl/4awKWU7skKvj+58uwngx0j6WVRVM1r8SQ1D17h8gkOjY9Xdd6
qm/TEIX4yMWNT/Aw54oj1IPdEusiPkxxVLNcz5R+FMHcSSGKSg0nkK1taW5w
vWS/tCM4LwpcNtmggui4RiPCRhXqh9Wwwr2cblz4SWXeHcJd+I6vVRl8mIol
xuRDW4IPz0NMJAynxl634F1uAtMPuqomQnwAcbtEhk+q4gaByiYSZeHSWpuz
7Z4bPqLoli7s/g1U92/gB/MjTVxr5jAeJFVubv/FoFOdtmZIzN2qHLJNoAfu
HeBG7hwHdANiS9LyP7NzjUjnCrVrkLcwYZW3Ky6BskmX6KlJNigk9dgeqDLD
oWQ4Qi8XFEbFJLvRWuII4Kk39PyYXv55GA3OmVT5Up82wVbIMYFskA5zdq9J
I0YyCRy6Vg7/JBJyr6qmg28MVdkd7BEmd0igKbZttJjHOpf4V85YrHRSldGC
TyfE8HB3PiwRuFnaLS+V4ZpGYaCgEAui1JF05DEovZfrF18hNpYmeOUEUokI
C7zOqN/vOY6wEaMeTz5B9myQaHN5c4OuKFzFE+LE4uWbfmelNhx6+VMKkNgv
zlFLyKp5nzULMbcHINdw/XOCmzMd6WEZ3oAjg0qUBWoPmSfhi77yvHviyHBm
aFrnnPbwxF+RG7rld41QK41TU609mjD+14hPXaYUI2yiokFblmEw3eBXefX+
NtZPnpiJZcxLttMY2Wj64AHD1kS1llABAX83PUvpl5w4HaOjHpRmOeaVg/cU
9+R9frGmHFu4EdAO8u0jt5rd+IBjGMoSTxtfLGhBooFWPMQNfyMBNe+/SMwd
QEN/UktMksusu/CEvjZzj1HHkrHfH5HoWB2q92i7D6Ud+vYvJ2lO8HV9+eJ2
6eMOFpQUZK4fkWGKqgvrmhqbEklIWGd10DjhaBr7armo5KADo+epV4fN8ZXb
rX+YMtjIMcj/PAKOf27oH5CykYsw1doye1WTMFDGmukIDKxPtlvntqazd/W3
6F4ler+LDHAI0QXHnm2inmNGvUCL6ucriWGV7ek7AsD/kkowefg6AU/7gk5Q
VoRZEw97SMansT1e9frSb6GGo5TxQV1f6Unm6S9LGwSUsD8U9vMApaBGQ5o9
uFrzVzimeaac3i/kDZBafQiIHEPpyFJKQzvd+PdTCBgKjXcudmBl/VcZ2md5
jYMRogPd14DHf7V4Y58OPQ1EaJh6sJ4qw8DWrXvlbeA0oB1jMod7r4pJdVEX
TTZaL4Zmxz90ELobKhPrKLcyWXomzYcF2oJtdbv4xjrD4Kg5nrGh0tiQxPHD
HmGmNo3faRskrJ8sBXLsVKp1DHgojOWIlTOJUigOY8aSCFswmNY4cy0uuJ4K
MSCjrf+kOIB5X2CJs4PqnansKmHSGZmKQkvK1S73htBtwFZ0SFgRsJDCvZcL
sdOrCGK/TwiE0H4OhNvTId9kGBPimQELVVrasqlUKE3RDNCnSk6NjVTmR7lw
7Isd2VLkbv5F2xRTp29qE/CVeYGKx84DgXCYvUoZg/IHcoE0736JPrDmh/rm
wPNO7UqFEXOd2BTGX38pEEch3OD75pPIkFzVEp3Tc+vE/+UarD8D01PbwQGP
fImpOU00aPeDBDIp1CS7VDqy/VzT3gFLk9AQGsHrYScUnQUn7T2xA4xHK6IL
tAVk44q+DKmvdZ0dbKf7234lmePS+qtITOW48EgCdrWOrbGwauSWukRUaiGw
EU9NgUnSMTlKPjlXqNK5AKL34EJddwI9I4vnGRjUwnr52Xu9UIRirWG72N/M
ceJFNWHTDUbmYYMlElTCFoxgK/noO3uaaZuf6ZDy07G3a8E65uiYgexHxHH7
79lJfLlcipOTEcOl5ZfqvKhFy2s/QxrDDgUbxTRZtNpTTmyJBpohgafr0JWw
qaIKjNoIKcewGFlfq/MQPzrnL5hIxJu0lF44gd4/4jRlzEa1FkxK+zfad8Pk
3uEA0ENM8mCX6x8JF/im6XOW31oSDFsL6VkpG1uwXuURaVXDkExR6Ko7Zl2S
/TsCzxYVqNgMUNttwtIvlxLy6mTGhrpJHHuttF62UKAxH2DtFfvEpsrb1/LN
RSSyMAKtJHOTD/EA+b3jWjU6n/nWWTcVT9V7yb2hTFdG/rabhxjWVVdDrcrX
I7zonxZ0e+qaFkrHaSwHOAyiw0o98NzGfDkYynbJaBYbSZXc8umyqE+J4/je
9XqHlGA6h/ehBPEIbohucekrLC0uSAiBzuKWFzWgOkDnLSDId99fLI1Jrg9A
nH28cYsPc548C8sTkwruIGT0KkulFzcSnwdHsBOUndmCSpuCrDOwIZtLyF3R
rEwwZnbHU7WfU7ifbyePmWbX03s85O1ogVLY4EfG0V0hkEHFpEmABujIlUpi
ye0PbBLAakOd4GJ0Xy8i59NvlIc9TqCZ76Ep8F8VVaqFJxgkecwISPKkttgE
/PG39Pr9reQwG2kXyXtXjBUN19CTvJltP5IXWT3ItWo/xKo1oZtukOHdZypb
zUKoMSDbMtGSy8eBZYNg3WcHo12vOzpAkhqG4wXGfVdaWJ+p56rpNpNPvmY3
T5QEVlJTwnCpSXAlwx+g4d+KYyZB9QGBlo11IfJy7JFsPk99Era508u7WhqI
4XOyH5EkeKQXUXvOgR4n5lXUN/vW/ZxflJkYzy39FezdUybLyTruGeriIpVi
KufQcIDBjbGsPI2He+abiqY+kVXzQKAKWlSpetnWlUlV/rReKa5a4VXi+61q
DGzSbzi8IAR3sJnAkuMSHIFwB1DO00PpD4PevnW/TiwNuOeHB+zRURMboaPg
T0i0PfDl7m4VO0mjiHpswc/7kkb6o/Bs2Uety3BDDyfc7wn7l+BEgRGoj3+z
X0KjTScV4Drsq0i3Hm3jrF+TYmaZ9UcOuqhcS2vVbcCxHec3/5So65noxM4Z
rNqQuTVqh/iaSPxxVJV3F3lixlWk/muQVpxocpHIMnuqTeXMbqEqwN0i8BNS
Z3TGDmP+4XleYZDZCr43fKxy0bRZdPtgfZdvZDJDLVB/CcX4vRtiltBzunUw
peFZqj1KxcfKU1BaKI5jgym2SDk7I74aStkcJvYcY5fWllxcPob8mfbEtDLt
xT1sDFQruGmX9r5dvwAE4UveBA9A0fqKZI1MFq8PPVoSFj89xY+uVJP+Uw4N
Xjrrx1qev1ejhqGcdeT6Mz5/yg4D+uG5FqwWo24kAeOzijYt8l+gAF7rDXRA
TXO2Agyy//CCjsGJtYUxIQEy3NWJ5UqaG83lRR0jdG/oKC9uLidtiR4RrXy8
FZ8zUhKyfDNitZRtCXvhFODOdDq8jwRBJIyvRzo+zoT9+sPUvv7NGVmkPgjB
UpRCqtNPA+5AvjPg8E0WJeM9gJjzmw59tH0WE5cIlh9oZ2EK5TWwazLYRlLf
LvehJKHO59Dq0bDdl9q2qBmoiH4fn0nWxHkc8kwmNe/C1FOLHiHxEOSDT4fR
pAKlrUrjhAJwzQU/Hc2Td84T9pP6T2qRgkg9c9j67aze4j6qrhze5UlwtlWB
q5z2VcV9SYNIaBW9o1Cwrhx+qMWunrClzuC2P8gI20w2ifM+/nEOqHF2/MEu
3wX1TaXEDWQlU99auiwdXmqGFhcFO0QzfLQQ66/TAPXIuV0li7yTmizRb2EM
04H577cpLLpiMkrrhZX6Yo5f5DXd/9RgE5M5Y50CG0mgLC4apgql1/gkQzx3
QqkJXWa0HUPRDtSVezbUVH4Wgwv4u5ds4B/hREovRNLzk29n4vWzA6N93Tp+
nMI/qbAJO7ARc29GyBaX+FhTBQtAtgPpZWBy8mBtxbtoWnbG7aoWTyg8ukCP
Ox/MzHJ796MnKxqOz4BZhQS29ot0UNaHOtRjmXaDHvIUEbjSIIFEaSx6Of9T
RP7rvmM1f1B15FiRjgJ5rYApOYKvdGf0Y44FyjYYyNVXB7Vda2N9TlCWCGC/
Ob/f5NUXykLAYrJHPRZcMJsqhErV4zH7eIq4+HxWGK5W0vtUOP859Z7Waghj
1vDPxnKKjBgqyoVbtZiY2c/5KZqEjSKl2I88XqBcKxw06B6v26uMHN8Tga0x
/7ivxteJwUUBtud7syq5ujMFm3aR7cuLUb6PMequHPj21uIxVOlqsQKV8ZwZ
qjEsRLdweQZVZKTVMdYjpXUjeScwVZ/uN97JtyKtOMOLXkKwLWVP29hO3XLF
7mH8pEdK/8+TMpXbvQVt3E/NewLnD1Zj5JDyxhnIhLD+vQB+2DzAUO0Yml6Y
rqt8x9oZ7hGmQlErfJhie38ApgpFKJQzT/3xzJOrPnLfAl42YtQ4Omy5CLb2
KoYVzTUNvwQoslhz/VKayVHLnvkrkSH8xGtxAqE5LYH6Wry9tN4VJAi7JBOA
CrgQc2szfz8u+iuax9a0NIJYQpydtHo6OhNhRxRm8qB/xoOpCIaMg1at0izl
l2kATvg9gM37Dgo0Cl1kylhBwZQwpZvJl3vHsM4i2pt1CFekmIio1Rdv42+o
7cp9pxfPGdHOHn/v6SPWosyycZCtpMujX+4nIaeR+zj3JRlXC28Rq6ka7iMt
qBei/fsNDZKJPhb8zcaEaFWoFwxcW+aNDq9DnrirHzYHmQ+Xqlq0cUrx6iio
zdUxdaiAvpj1VT7r+Xznqh6sjV0xzIn31yi0oHCOigVm8Qs8aE6TnKXZWUy6
hlTxLWEztdLT4V/9j8+Bz9xhqnuzsazRu6uiSHRGN9J6eUv0ccdR6WHtk462
3f2bdKbRRjAb1jaHRk8dQqtrrfVIfPmcsBXSse2XAAjPpwfxhpoYiuUNq3QE
gduLBZ1TPUqIoXlmd/+fl7D5mCz25O3yX54W5HavMCWEY8OXmVhYL+x5i+in
4/fXaKFXQorMsct6Z8wIJ/TvhohNTpEWeZ+SeZupiy7kpm0/6m1GccmbDRB4
cALgfm9uMMyMQMxbsBCURyWBaXSS8hn9UbgdWk2b7gvOZa54jZ8hTVGt3qSs
AqeEsLo1axSc7Ii+7/OG481mimHLg4Gh9AsoTNm768Ipz6vzmT0JuvEFLEPh
JAX30esF8tIdIZAisxl5QrHM7fsC9iMIP5+dW8981c7bQVQl9yf0aHl3NJIE
xuqpQ3oQO+Ou0eEFV29CUxCGEEurRM+PDrtVMBkrap2m2v8uyx2u79xgou6j
3nFKxgMTPR/NVUKM577QfmpqGDnOQ3w1RHvsFTEBjYxnl7T2WC5kHla4BFSJ
jMVgrUeivFG6UmMib79V7MEi51av+BgP9zDguJ4WjkZPr82T+KhL4MglyD38
1UACorN5k7H8EScCUKApanwxv3dDPwOIwFcJ0qFvEvnBTZq5eST3PRJYikvB
CZhIS+4cePcLcWLE2fpJhrpWZDE6G152zpB8HamCyUuaX9P6ZhydjUpZwymQ
SacbItVzZMVHMTJ5SWl+sBWnxUDBbuhSayX5Lccsuv5+J0cSbGXqIp1UMwFy
KlVXzdHSuIyS0BQdfRB9WO77v7lCPcj9lWrp+fnRV04p10Q7fqRhZYH/8eUO
EXh8RmnvZ7la55pqmaJbG+nWEPxwfISskJ1dXAjYvqTtT5df/QdOoLtsIBjd
nM5cxSIFCVTkPAYo7GZKJggMDVf/TbNUkksUyorqDe/YBhVi3KQ0b6p91qwh
kmsuAInxym8C5e8gs8l/UjQsPCfB1l8aT5Iv7Trh+v34ItMMxdzjjSuT+yP4
DMvqQPrVs/9+g97BWZQQu9itrb/OB4PyoCwtZjth0nS6j6rBH/wGx1V4GFNj
ckORGg5pUtjAyV1LlVlczaVft6M6LT0NWpQEku/R1XsLgO3ROpjP4Jf+0oTw
2xYWp0CBTSCi7tHakL7iJYRS3t43du4G7Io/VgIoj5SApyq0WVhDVa4Ujiol
cYyarhTw3FbQ0uk9tbbiMq/7sZqYt6Y72wPgjWDLCxLQBgWYjlcIFOY3gkQO
Pe8A8DgUts90jOUQtRd1i9vUrelq1llDzwYey7vNZCb81XeooT6DeFGTfA+x
tNdVCCz+pidaAJbpCC5d4Yw0KPzfygrMS1nXD2/SZA6aD5I3XO+o4wE5KrQ0
83/L4BFvxeFj81xTmJ5QwZaBrI9dhZBW/Skg60SvoUiIC1pS76ZCs8IGEixE
Xm+otgz5Ct5Ruqj9sTqfbFIv+4TveCMLJ2vuqL6r4MvDFqr3J6zf0C8emD5s
ur/wQxDposqomW0ti3/XBizFMQZ/hut70tNAosK+VZm1Mtee1/5l56lst/h3
1e0bJxw9u90jcbJOCbYCsKfW+yb9ycEcRXjPQVs4sY1lgXsBeqRP6ebRslrH
cQ5lKp/aT3H01YU2pfbMMoSr/BK51mGY044/OY8dv//mR/a1hfFjNARI1QN6
S5zt2ugI+lfFmVQ18NsViUCK+LEFElib718Hd14EUV6kL4uYOgpCerP0Z7/q
sOW72EVxVmswlWtClbQNO2u7gK2IPcHWMW8zBNVSVDLICbNZhI9TGPYgcrDL
iTtetU7qGd9BoOACZ8LB3l+U+gSm183zDxFTlIFQQs2G2LH/7xAEDua/5WfM
iqKq6tnxSmqxBWNRIcgJjC/njR0TWaz9ku6kBLik8DRPNWY+iMb676q0KxsM
fLmiIazHFCsZZBUhJfoDCPvCBf3goNZKoXKpcmn9LqjCOsT0/huFx8oiZGSs
l5B02pwWSxzIAssAnWWf4Ic6fEXBLJ8XZDHSp4SIkzGqYQoDauyBfrK4l04w
VfrcFSDk6pmLp+FG3LxyfH8rYJBFFB5g+IyOsJGfqG8FVZd7LWVXGsPOvmRD
Gfaw1O91eChrC3iM2A/B1nuE6tj2LEsx2SfUm/qLZsS3ix2/40MXzTLBDmbs
AQz2kbv1c5imMM8o1kg4RFABwY39F/Zi9lLynWBjRArel7AcEHIQlzWYD5pu
DTVM8MQj9X1lvybnDsiVj+rtN/ROferJALXzZmx3/GnZwIv+DWb9DTzVH4co
VGapVAWGpHE+AOBOo5nmVgIeBYwCJU+deu/8exTq7UFL+a3YTLeOkdxLOblg
rm/3sOMcFEGn5UlGyE17jehf/RP+9ve1OF+kQhYrQoK7lECQLfZLtrW82sL0
9M0DEZDpeG/+6zNbW8ybcYtdFvtmXgYJeSgOCq37fwetwUcQL78lPCN1nv1v
kxk4RV2XPk7YnURHPydyo/l6rBfA1ybg2LLF0ulgVwiFBNU7UYiMps7EoQTh
+TOytsd1G8PjxM9akRbBV+xAm7Bxt28QTBp6zGYgKtTEw/DP1D9GVMOjGOsm
FkNUSXpMin8pbMgqXEf+2W94YvZe78EWFTLakIoS7LWA32Q187hug+oK/Hpw
zXsvI4yLFFZj4M0gT+xM6RP2r+ActYs7qS6z/6dVSZ/9RfSvU3qPANhzmBJt
V+lOV+2axOghRlR3bSOSX+FjH+mmz+K8JrLXl35HXELgGWG+eRx292TLAhfP
qSzrhJ8ZGWX34WT9/75XBTnUH7QJm4sO//igQuABB5h7eF5W8kcucyiOk/vl
RHEY6fVVekgq49LoRgJzQX0pVGRV5zvIkQdUfhb/YsJTz8QixUUoGhbskcW+
wuhPQ33H/J9zov2o5+XbsTtuLyo+p1CFeSrvPy79liXwrCLpzhBaRJBgcIax
XOgFxSq+XPyWt4ZNstSj3z2oDfxq38TwknLxOP4LgmB65QW8uQpPvmz5BW4O
DhipdJHXEtBSTgPcE9CD4oi/EbupAf3oIhdRmiRad0b9zF2ZvrESpVXIUehB
iBUz4xmeQ8LvyRmp16oMUUyvTTJYmxt0Auxu50uZYptY1B4B2z5e08ow7TMq
o58cQ03E0I7XK0LJbJE74ar0T9heS/KVKGvwFggMLcOxfXBFqR15Sswmuogi
R5O0wB/jPEy3YSZvlRcK0oGzY6bA3mymx9PvtC4BmAFM24WivESQSLRpABjn
W92PFjQRaqJVsnnsJ0L2BD7A/LWAjFc7v1LexwYYarG3jtOPnNXuHYIVA84/
OfF4ow4bCGeJeLAtQdkPtaYV31x44/AFzBNs+/BPyJTLBB7NlLCPo6WWxBWX
IjpaMcOPESRIrwmezKJdDFIzEtqTOHhfOlVd+sXOcYAPbBxnhvh+I3P2zmZS
vrnVvDGBKHPo6S9ywmxVLp0iCHXqKTkL9vvqaauQdE1ZOUGNQ5Qwte2iaqP/
EZu+4qH1lq1hDuhYPpoq4d2sz1TmaJeiAxBlyrIBsMYAvXq4yLLSeIrhvxRL
TIegQBaMV1t9kqf6+esXBechYcel2oTdJ5/NjeJyuV+mQeon24jkMadhr97L
IfYe+8prO3OT33Kmbp2FPudbYYft9MT1fVkgZndMI7cdx0+K0dU6maWw2Whh
PfOzAHzHjjl5CV8sVJd2vMO5V3DyJkhtxOgzreD8ujzMnrJzmWpHkyoV1aCg
8zGAhJ4nnND+r8OiZqDFokIr+fzchwZjfd+RUIgPlEHaOI1ZNq8SedziYAwg
2Zs3Wu7CQPTRvRzhl/kJbw7ZbR5XYhP/8ilHT4AozRxLo62cXCZ7DzY+ra1h
lYLvFAuGq6Js75j7/ejKE43R6VS+at1TBPYW3ls72bI3bsKOk8gYEpj0dhAX
/NUA4B0jztq57uRtohFLILxw3xnt1WG7+2UBq/saHUZqPrXiqdqqrgfORhwP
Bg6qBVj1ts98w/ZLdbol4qewBe+4wPbYki7ba97zZOFm5JJ7/t0isIwfyQcv
e6Yg1m+d6tCGC6Ciy2R1O6HheviFsHfZQd5tSAFvqNVAUMMkiiPSyls6LBrU
I4TUKJPd3vtgfl1oGyOZf3uAuGxtQX9MjeKWK6VdX0J7o/S1PGDrG6pvpzw1
N355eTHnXr3tRMPTAx+MVn8zoJv0ef9PdLrRMxbPMBjKxyFMxRRdeU6Ae9lC
MmACzbG8FGwQ5oQ5PMaX6Dua/tHPfUh86PkwPtnN4NmLdQKX2E4iWJ7JsE3w
zJNOtaY5w8rRtb/QTWF9bnS+wvabi9pzphPoAlzAtxRx9k125IR9GbqpSN79
px6wGoVplqKHqZejJi38qJ0VoogS7LxG1jonjuVSxl4ktpm9L19cFL5fYzq3
BOgE85XzA2aVo4u4lkec6QPm6BgdXe9AqrvKa30dYlb/tbtiKKvo5cmb+7nZ
4QzfrLgG6uBN/0Bx1OitfC5+KVVf+ozdZ0wrNDCbrr5R6MRPHluCBITt03qk
V097M08KtpLUZKECC3kb/SW9RhW9LmI7woIN3TAk+gUGwky7/lq3RKrWOYmZ
FWOt/YRktgksFfk09LASodqsnUUiOajGtnhZr/r5z5XDZWZuuyz4VrYh7JpL
0AbHMPs3R/We6BOPcEkwKfoqBWfqSeOQN0/A46MY41snJrXRIK+WqAZREPZh
1efD6wFRJePGExDwF/hVmnIr228ewaX3StemUYRImYThlscCEQmJdo4rvWTV
ZzWeu5Ix1lr3lxRIpk/9E35m7PFxBrzmS3A7lCB76Loo44Tr9ozuQxXHq7QX
DcYKay1+8jEBHSPcwkgRK1vFE4VufOZfYXw4mFjlegVdQxX1W2b/lwf8FEdM
O/yIdzpdxttkwizcBld00M/8kAMNbODrqNXZlC4ZHy3+DOO/IyjZSfmcKSfi
8Kuo/2q70sItv8fOAbJfdei21NO7hVlou2ofnbeGqdPqvMVfD6gi8R2c6l6J
TWrQKF2eNq7du7dlhtu7/qvAgQAUuAQ+vytwFfUGqH9eEnOQ/s8bE26cMQU0
At70n8TRRrcwCjlg3iD3CWyzrDPOPA4/hF4l46X6kt6qZ7UClU0P/mkNAr/f
neA+vSHv8bMktRd/xIvfie3uaW5Sx0v08H2p4XXn6G5nTNN63go4b/jIIOYT
Ow+FBou21iTlJGocd0mKKMZ+zxXNSODQNICLq1SdpbDbrIv/JFe6wVESPX/b
YUqVgXjZHQfIG8lksP5h1Megys7s8bso6mDCWVylq9dnS8M6hBhPjsvkCq/9
HGLy5ohzDRScZ7iIO63rbc9wBdIbY98iabCl8wVMVqDgRmIKozUUVtQ9pSAV
ljd1ZgMg+/ZLkGG+oHqPbp0V1iLe8VaMrmEFFJKnJ07N7WOGLfpfpGNLOtY4
pf+8Po7QeaJDa7CYsA0DGWb+oCpearAVrGM5BWOYOuCO6v6aMeB9nPW3FzTw
YorRc5MnQczDei78KrdjXfYvM2DI9zE59QjYwQgjrzVftLcmWubsfXWIMX++
EmJ2IA1J2X04L8uitk6C9ySjjKbr9Gh+sDTZCyz7whcaTGC/TTvv7aPmdN77
+UgKWW+bt6hF3JsXlymCRVEwb0YjHeLOWmXoGkPRREKPtJIVlQY4Dhl44VFc
oCkjx2g3ui/DQtvWBSDSdPVs6hpih44M5LA8kVgtKHBB3PdGD7YHM7O7XuNS
e8lHdwOGnt3wb79ElXfpod5BO8g/JSQgnySEEKCdHePiGuZKh41pMGDjVkVI
hPbNXLtzmvfXdN9QAHBsHJXlKvAcpFUmpJu4oDSnbPkNZx8jyy/tc3yBNO0T
NesIQx2CN1emmyFvyv9v6hOfZTW8M/xhbOaGDasTFmDdLL07pfsfTx4dBOr0
qfViBWrR4rthOq5cRgVMbQywjU+UwbFihlToeJCDEEgufEOmgjSg65cLxavZ
kMa6I5DCfNwtP0aWUX0hY6g3I7pNfAhcwZ4gDN0kjpK6QD5d/T0s1FlgO+1P
GiK+W4ymhcRJiYLn+IJcB5NtLV9sUQuAwF+RE2UE3lrXWR8WconqBh/QugI6
1Aod3tvL0R6nrFy8BrX1Aigvz8tV5L/dJDH4FeyrGkqFtFeU9/P+JeJDPDd8
TncESSDNEFKezJzN2Vr2fVsYU42sMk/hWtjfHrHN/PwlDZ96xV4pgx56Ej+L
nPJ74k3FvBILD4HSwU75vfbxr1dIv2ZlyKlzMqdA68Hz/8cUpMOfoJfs0ihd
wnj50KMQBSTtvhvXlDltrjG0kphreP+beO1VDLzNr9mkyv8k3Nd9csaUKwx0
s6JZQohJ6WL4BdHexsh0ofCCQQgg4vPeCWBBT6bfZXIuoE4vv0F5P7ZBNOpS
s+rMD0eYae3CTZ/lEM2xKIGR8+ih5oTpKrXA3vdLu/aX16oHjM71jkB8ECi6
vj+7qZSNskYavXMbouT3xWOelcrOGVsz0t2aZr4+mJAreqXV64+rhHCjKoBV
VC+Yx2+YNc9AOXa25mbTCN6nx/+ypGQbo6UNmj4vttEYviw2S97RHPcguGBb
cuQnIouAJXDpulv9pGV2QKcDd+El2leBR532SJ6pSmVz4fx302Yad50zA8PM
buI5tzPWHY2hf6+drXaSxe+/X1b3Y3TxRs9Mk8AYsEr9geTeRVt2F8QlWarV
ZA75xMLxBA2WXC4iRIzq8Bncin00xA4vZNnyK/FsgLJJfRWTLN5fHobOIB2C
aRGDE0H8aj9IQF6MUCPoxkfa96Hm+T4a4UG/47/K9xwWVdm6cmrXMhxKqzMX
lbfBh3X8/6+MaAURu/K8h1DXw1w6QTRfEzEtzscMiLqGwlKRj6qdaeIoo4sR
qY/s+4SNk0ojA0UuSeumKoGU/EezjNriOIgfgwDXHjmn0fBltf7jChGjR6G+
6uOZsDj/vbvhA5RM8Fa1t5yc1Dq6M6A/wnHE0C/QsrKP63oQVjkmkfDOIsm4
M7OvBfhBt4MDtsVha72Cv2l35VgC6qEzooMuvb75S1VILdrmQbGemhsT0YnO
me6smWCCr8IatKb7cxMeCUXiyq9JMxlg6fQPeVi2JbG7RG+0DyR11IECbZsE
BTK9Pb1hXOLUY/LhkRbABa95i0WV/EcPJMFCcIu5PPElypXqk0TYdRsueC39
cxJWmbO3u92XECopoE1jCL/b1Exfjl5lvpLLXP9Phw8UQC9L9eSYctAxK7Si
5z4vdQ14SNf8rQf6kOVzhVTdRvDP3SNy+hWl1kOmoM1zpwafefwkeLWBM9KN
Dg19M99SXj2AWuTb67FcAJpTpAp9VAKGhi9lVaZyHZEGxGtiD+9YsH98VxQd
vDUOTTFUySa885YPVwXzvUpbfjUxk4vH7+4Uu7bvT5r7sTVQcUODv7AQnjU/
2NqOvEhTNDM2BmW8CQz4JWGD8DnTcEo3YXxngRWLK2CkfNqJJmWmiVNXJwmd
VuMZxUsVtM0Vzy09RATvWuNXJUdxgOsPrz0RUyg8hOHR/8g/XFjPxoT/wCGj
GdFz1BJ02sqQ5kdJMX+dVIThKj51eajHLRhRSE/F16H4xHWwDLmwjsgXN34i
CiS+iu6UmJ6pI3DR4mMhCdKSYc15v4j4c3bdI3Op/r4YooprNt9kDaEaY4CT
R5ugBGhP6LYTOiSEoop9Md70cPs6qO7BZfS5NZykPjERMhcMRYYltpI9/3Lh
/1vYel0dEPxNRc0+FgdCgVt+EPoFM8EvVnwmHNZSNc4KavVz9z/ZkCpal0EB
dxlaAenZ1AnKogPaJz5YfT36X5JVzBzvOMF8f9h88OFpC6POCuYtZLfK0oZX
VrJqvxe9klvY6JzH5XVRiqPba8IrURmqh9O+a63kDJmpyx2L2JT2Zl1GFSzq
ZAd9A23w86R5mWdhiNUhRADqI8H4x5Wmr4HaEYFu5IlwkqTKxryaTXUJATDA
mz1UZmEI3t6o6of92e53KFRPkdkybwWWsDg6eKcsZ8vxvKvJL5gLW4T2lqP9
qagynA4Y10BStSBxiGZnECQC3Etg4ueZSNu1lwwEwk+FyEKX2xIMQjowkgDz
TUTeDBP26KOqOyBJdOfWpnePMOHu3xoPeAA/HqRmQVSYAWap2xRg33XdhLW5
qvJz0/K3mdVHQXU7amQTLtRryH+beF+pbO/YQhXX6lrwQW9/72Q71tO8moXp
D/TJQcXVel/6iNhxuq9gQmtp81EM7jDsDNGKpltNpaYeFVhPc4a8MlPy1w3b
o0pkRXzyVYqPJogDyNLbnrvHu4OPMEARJGigZwRNCdKYW/pIuE/DNlqOuE+3
vRJaxmRzcZ0DYHlnwtqz4NhokqTA7ydvNZtYpSKguZzZMSlCBz8dxR8igLf8
32/X9fiEMBq6rdl3/5p3O9gO0iLZ4QAz+YxYYagDZTEbwoST+Lq3aN8TW7Re
nkxuImPl6spWhHwphb+bwcqCX7C4MmN42oiDuLrriWz4gfUzPKVgCk8EaDQs
2/V5tYWKRL5FWe87xUsfWvTZp8ZGnGm424hn1DdYXPg+9vUXZ0sll4fSqgIC
q6ybL4Ld3bf2Ih9ZcZAuhOc2uJqK7M2eBReAtNoUW5B702k8P5rA2Qoyw92Y
DLRiInd4ojm9a/fO1cT22vALHCVxgELfYkKWP1ok7/2Sl0CZ9vRAd3ZUq7As
XGGJci5fLA4SSckvwYB4xdq2pWvxNWTMm9s9FYuWoOrgMpKcmDVBy3KIDmZq
oMr59qmP+/uTz0Vr1cSWigz3JVkeQx5rkgEksEQYY5oMxNrpR11aeC99Qv0I
joBKxvSzuR7jw1LcGuWBmYbb1JpuBb4z4JsSW9m9Myhs4TyVcqPIu26tBsAg
SKJTg4Zkt3j0AzPBbLvAyz+fTu6fyrGCdio0mOnR1iKqy0xk/h6Z+18O+Ypr
pVjBXjpL9Td1W0DESW8JfhIekh2KUuWcvyk1jCAi/dvV4eIRQosuw6hkAfyE
Vz9r82fx57NS02sGjqshDvhc4s9lUkhp3/ak5NKAr8sZPA92/RCzifK15yX3
6l9vbKhSyAp86e+KSzHct6QtK+frUf8kf1XdIhyudCosVr4+mkCSeKGO5us5
gh6q/jFmEbBCu1wZL0+dKWQdgxd3ozNJsnxMVov3xk+3Wtqkg5zky93Yd5S4
a1oZbmciRlAjeJAIP2oivlSpmPmznOmFeoj76NEUu63peGOE8ohGJ0rrXHg/
tMlXxXTfh49ufrUIHa9MpmjYmpsikbfk3Xj7qD5d2F4aOFUlgbbh3WKcwhJG
fCkQdxHsi46CmEzxSHu0Upv05bn+Gl2ZKDadNIkGjg1soHjrng6szqJv/WaB
oOWDzVpdGbZrtlou8cuu9q1ZPM/2JoTrxcQPyT8QmBboKC9zJabdWt3CeKPY
WSB1tDAGjBY2Mq4zN1wO/xKhCHkSj4OFn3An+0ZVX5GiqG4PRH3Wu78HAf35
ue6QPqxaemU7frYnaXEixaFI0g1V1W9xtp/DscB90ntqv1AVxgJUBQiP4fNJ
vH35tJ3nGEvf4lzfFPn7G5ImpvTVpyKlETVQNGnFMf8J1WikNT7oMd14d4Gg
Yz3UzLrf9wqHB1VUoQyA+XPEyzwc7nktE0zeuQOrmDhlUXUWglhZr55YzWWQ
ycIvoaE9Z7B5vJixn33FlXEAzNxxV2NI0gik2BM2ryYLFZJGEsuubCoHksq2
xYvBdLWKh+Edg9bAbpAAh1KuX6Rt8B5BQzBrXqxlUSlDwQGa0Wr++VOMUias
ok0Hhh+hVSYbhlRyKFX5tljz3zQvH/E1QrVlS2UZXa9OsATkKgtG8AkH60ar
khucMBs6eiJ+g7oo43Tkh9ACXTb1CgI7ZdkcvaZbTIzlo8OrBZfoFO9wKD7T
UjBFS0fLAMc2gfKuxctTCrfqPxjXpNvT94QzyyBteStnhH05PBcvf3P3unNS
QXY8nCyvezOaoWI08cEqPuZWN/5ZhLfTflocSdgyPrUc/c6O1+FSqcWVN+J7
laiFW/sbRuRgAHulNiOOIdBtPuOrR78agModFFjP9imXvKcDkutcLuv6CKfj
Tf8W4iEvSL6/bsQdYbUUFeWRxftJWfOTg0YGU3+piLHkYyaait4xkR/Of1IX
z0ESES7HKA/U/yhyJQQJ9Ed0iH7ehf3ACVwexaqsXfnAEUjwhzev4VHiXWZj
VxEWuvsbHEUZDBGkjSft7yycbSEbueJsgApVoNeXJ34nFEnQmzcpwEpDtwR5
LrVdi9lzbsrf+HuyvmMqZOeeQp1lBXbU4po/HBRCmv/DCCyekkMk5BCJlxjG
bb+vL72pnJiWDK+oBb/w8C2UQD/K2KvXgdsgrwF3ejHaInZaqSOBHQ9ogsLN
H4d0gfy5dFevDzp1e1epoO5c7xY/1MRtumdkUIbri34AfHtM8dzq1TUV+5Md
pmf4oYX2HZi4lziKAzbvnxPKWY3s4iZw/bThC895X30lcKI0gAobYJ9Kjc4+
DZsR+cEWZlp/sfHsHPp/mWBT9eJ6DVII6nCGl/JATqeGmjjxyQTVHMYofK6a
ZH2yxESXd0qNgxfOkQ9u2XZyB0AFq2XHVOxHeOxpv9znqSx43EQPRtJzQnEc
2ESJYinhpz7G/hgb+6jes6XawXIFfMUtbJzNSKCqySxKyy7NRxaRKIihuA0O
rykZpmffCN6U0zafQa5iX6l47ZVsgAhFo3LFk8unD2umR4czQtluQRFiNFJk
Yh3bxcU+BlvD0tuhkGp+WpehBx392K0tzUnM2gL5gMre/KAX2MRMU6QUSdto
ci19Pl6Ccbs/2DaAXqAQrkhi8yrDpSSvx9uELS0czkUrKNi5UfJm4mwEhxUI
l7SFLDOVnmFqqGguAHpbxRc3BMdc2cHpvi01RHZtsTVsCvGt9pMAEBVk/iFw
ynTQ/LenAirjkZI1uWbEEQfArT8BOpFe0qTS8wfQNN49V3YU2VbDic+BnZwV
souJF8kEUTptJB00nJHrTpnNVvboo1mL3qnisKz5aCQUJAQrIeHO6ZYjRp/Q
xUFjNxu+mNN3bv5fTLwc1u5VP5849DoYWpKhn39tUemGIp7i9esuA1nIn26o
ChVVjHqCE1fT9VsG4OZIvAZHgN01/EKd+MueXLscDJLC+nwAPeVPmh+xSKhv
/6sWIC5mL4guUZtV396NgrNTXQZwUh3EmA7rm0e15ZbwD7o73WcctTGiGreA
l4+RGVdBfDH1qR4wnDGUmlektb2rtKkP7/4EdqPzzttVdElupUuk0sxK0aG2
W7pHgIxq7yw24HLVhO4REQXlIrdm+5mFD0AeBL2YHy8+CtWIM4200LhQRMZ0
jIZ1HV54ZFt7jyJ0VHZkEb70EdLDljBudmVa3tYRBoGgYYcfvOYv1GJHMWqn
WuerQ5ELQFWEgTuwxthn9rrdJAyfd3Pn1WdpS0dRHnZJBdn/RYyEGsO+ltRs
/TxSNFqSQT947Q8upBui0r3TsPRqVYFCQOvoUE++5HuShJHj7FF7krU4Sazx
WunIfAdySmdcmjT2veIH//9p5VOIrMT0TX+lr11NGm1AtF5F2PnIMUWLOoR3
auQq1MqT6hkAu6rCOI0WddO3PfYMcPmKH/W12CqHnHjVJGJkLUpTcwPRlOim
I0c+jkKeIN4olFL/qcMOTBtsQyt1BcX7laPXyr8kV0Fjxh0wHSmUS83ZUvXr
4Qh/igygh1XogZSivduIG1DacDmMN61D/oxJ6zfFH6Gd4AY6JV2UB5aAkkdE
yO0UqdLJdgfpb9FlguZVoCPVsy+NQRu/FxNO1I3enjMhqkI0oRHKsSG5sk8v
nR2ya7ZFnXZ9zZbi8msMRDI52QJ6I6hxP6Kt5nH1BRWEmQkKJDiXOypxfpd4
Yj/Hjbs4H8VeGu/zKwjjT/Cv8Qc7mr4QnggYVf51lTQQ+wnjSQtQ4wjHydhl
ys3dO+Yje6t0BS7KUEnNQlbr+9RypiieYMDo27e3ZujAzdAJUz7rfLOWPARf
L395mLxk6GwmSdBzUyL8AJeJbRwmfy3c+2xh9TVPZDkT053Im/IJNWDEFanl
8PmAoF8ErSh0dWcJTxAOxvhgovkxwo4SfKIObkfxF3tVYtgwFERyZVQKsNue
Y13guoDENHlI8AHf7C6YPBR0u36mGM+96KOSKHS3pMLDEfg4nEXGiQNiHbtw
7GUubjD2vvs1m6WvfNyMBsiWxCKBOES7q11ktXEnJsf7BGn7gDZU25R6Vnqd
2Z0YJHHm6ywNivB5nYfMFwPiIZoVBQFpNYBazokRRe4hXM4QPJJMtaH2okq1
hwEkVuzIH6nuq8UdMdar6KiC9gSrLFkkt1UK3dcBJkJIE7HLffzaPFq42eeK
GX8v5NugT0gdMW9lt+PUujUsCuD5Lo1MMvpcBHhVBub4vuGpbNl5+endd3lX
o7m7dNeHpw1yWc30okXc+7t44JvFT5i3QFDp9f+gLWJWf5mTNiidy/pW3hRA
PKqgjZLlULxY1cumHyjFJ1H8sWHtdvARPuhfSxt2+KjYJtKvEMnCB9M7+Xqs
QPl6f3EY4hc2IYWSecWgf6i8yYtWp17rCcFi+GLTXdGwLhPFY/dSTjCczHYK
HjCtZ86g8IGKS/c0015fHpaRQPpXQMGkG13Qx+JNPgoh43CDd/Q0xYXizvk0
u63cFqUzF2LdeyY7NG6SwLWIAtaKNeizX0KpatQbZHlw/oJ0lG3ylaiUWbU/
L6Rk8txWnQjxLSkobflA5j55lYJ0iobGqls9/yZ4gOFc2f8r7CIZVqDdkPlp
1CcIioY5A8xKZwCsmnTQoJRAeX9afta97Ti7OYdh+iC31SQ04xoLtSGJ6kHM
IZC2upTG2sRLihBYTWFRRKZzUDmVXo1gc4/LJU1HjWQVCE9aYE4Sxi4heA9o
jBmmEaKNHZDmT7ZrK5Qu8YzyZqY/GKxDv3Z4H+WaMnoxN0JxsxluFhddMX1b
Ra7ZmZJvRzeAR7turkYF2tYBsQchXOwcxZNckFBZRbLsHPoQhu31f3DJwpoY
Uq/iKeMOyDxgiiDu0zOjLky+YYQ5EYuQ3IuViEatx3hKF88f5J/BYJOwibcv
OnTcTHyAP/5L1xIFLGh8tinnWlJylDhG9fAmBZBjKGOsZK/S8X95kuJ5jVCV
ICm1tkxyrcuvMlokpJCrWvq6IKCBWmCLJ7Dt0gY/mCwmHKMnjzU7XkijlskO
iK+S+D0wwmVoVGnELHNrdtGFAQZkkDCME6NeYJptjSw5YUONJmbZywIglDGH
XWleO+eajr87YoWxmmdLzkREqzglWSGWX1KCNQbUuUgLM/cf1GFgJu9aFebL
oAAzOWpvRo9F7/TwXS7H+TnjCsqJmq859VzCqdcaX7+4aVPK6qyA0/C/KFsE
nPKSA0t0Qn1sbWSGiAdpxxFD4SQKJlZ+HJWgFJhsOb7wSbKMHP8qzjRhj7Av
Brq+BlR2laYvGYjIc/sk3a2DfTLo5FA9imBrpB7LAesh2lPe1x4aWlxKlW3+
THsDcM/QXDvOmLhnaZX6O+mMSvoQPBSH2PtvL1gCAq8/Dv1WQH5UYxuzDz7b
prwWLXu5EgxeeD0gGnB8cmZUkAphIhKdmwsRvD/cSPHiKqxkjrmbCmutsTTW
GCBQn5OequJA/zZ4FB/KP40rm133xRDNNFyt7JVU8fzYILWPa/AyxWMGK5zy
z29rkLD3SNpSmX4TeznhdqF2QDLvUKOHR4p3Ixz63P5bKAObjF7XgN0KWBq5
3n3TjI7CQZJArpMrYcmKbhRBKK8CY/XWxYpoZRIn5Pkt5oe1huJMv+kON6Os
eGexse6FEYWySPmFzBA3GPJBGdatCERteWqR7etrZjOwqB/MUhvhKUTMxg1B
m9vC4/G9k+iBI19d0T8Rq07xwi2a4LOD1vZFmKwXWt7dPhzBmsLfBRcL36PP
qzgqfO8TnZzPGx+PnLBrgWM9A/e1AonN+nwwD5TPgQCDLnLBmqWD02x8Y2ZE
vkm8l9A1EuKh1y//WaZBAq1lQXOCOdX8W9cUEYq9r6lz1QiFRT75ZCKqVQ5E
I+R9EvdaveL2OkbGTpzxxOs59wHbQeSuEUiVw5Ts/W/53lKTs0PoL+7MktJ1
YAT4uTRIR563/7EkT+JFvA+LwxayzcdSvqh/wtewiU/b8I3rRzeQQwbqqjAv
qHYtdfEVTYoMXB5aCkDLiO3DG8SzGlPwzoTyo9Vpp78Ob+Rt107CRs788dkD
HV8rjEesbZWGxtdQeJtcPJ7uatzWs7Siv1x2Eh0LXV+VuOhIPsLwd2IilIK5
seOgHh0rG/0kcMwuaONXH4a8R+uybKnOXK8zrjqlVoeDhR5RKb0/zmGrbZqS
bFFKwtO3ZruL/Je3ThZOz1MwTrt0MGlwjDL1b+Lpree8TWroLOCv5y9KaUz8
k80RlpZGEnncBoXBywaKi7W0sMlsFqFtxNPe8jrNzs9LJHeoj6ZEwhD3XAUY
l2hGLO2nKlyIJBZKxTOtvKfauSSgpVGh+XZBCBHZ5l2DAMhs3piT9+wUi8+S
5AKhyVLRScxbf6Zdb0I3TMn7Ayk60waq8ASL+bkrVo/b5wVQVokDLb/gBP0u
1h6eTkT6iCoF0kWGfhg1irNTEKBTrLcogFp/W1cs+2b5eDJKVluFTRFk/gHU
fnk6UHCsOS5W8Os/Hozea4WVGebYp4QlIySMXl6R3chPsZ8zcikdUX4ExiMG
ba9l5QhhLsP/1bqBbEbXjouFaeazEkVI+q5rmbuzNw0hGWzl3uNkeCB+vD+H
8q3zqKK1va/CdqKdNXI9J6u6a39l7+umolEejdUXlLTmaSj8TXbfLsDM8F0J
EDoniwmI3GyIVXLjH20X7jgMWv7WGOq9fy8a+fyNvPg6cuX0kzFjJg0DTWpz
kDryrUKoJEjNMs+97mQ2XmNBLclVy8ezZLPfTLnXRJW2zzdpkQ6ohDkwe7Kq
H2ThMIdrSIg6iTZ6a5kcKK56S2ustUdhtIoirv7XSKmrwwNIq1WaTG+Q0u8+
qcDQ6WyoIxnLN1q2Gj2RQr2WjAtt7AnryPU48SVIZ8OxfsOXVYvaxeda7Z+1
uXhrzFDPm0Vc2/MT+SiIMkcsAg7+cGVIad+xWKA8GXTqT7TRQfe9fvFUEDCl
PYBu30n05x/n+5VywB7ItiFIDXmG928h7nFPh8RxTAuz32X22GJ0OkfwUz8t
fkgEH/zf3GJnXtOTPkc4inuHqcaSfX+SEZEki315aOE74C5XGlCfKiDiCXdr
Jfrfa80GwkBwejdJR8NeYZNtJuYUX0TvqmYO75JAL2Mf+0frDnKhUIPqBNsz
8EdTEPURTZX6SlLyuiNN7BdfVgBxq4EzHb5XKgCcWeLAuw19h86koqaIZRSW
XbAp9WwuuAnEpjXnP/9AwXxusAvfelunT6C3ax87JYY7fInoCFnn9qARdC1m
OAOEx3oL/h1vCDjVz3MiTlsExouQ6/8Aa5Z4pllAPkrS+5q+YaQczuZ6DpFw
IZLCmVI+V+qa5ERohPrb+HWQjlT3w60SESqADdH30Hoto4U3owytTwqWlwNV
UF+lXDqwBoInlIfgurgC0YU6MP4FQuq0M3hEYTJRY/M5rD2sFOuHRQ1gZWir
MGWknVBuL5MYDQC6mbBHo5IZn4XgKiDux+mn9oVT+B7LxegCPCqLS8nzVLee
xM7OhUrWmaEipJEGVO3n3QNQ58fvgreGOjkF5PxAGW7xSEemUMK1rhQ5JArd
VcVf2EQnQAQo3KwWYb9Ub3sXdASpmWjO1BPTQDMa2b6CRXC5It8aaggXh6R8
7l0ycu/EFLX+OIuxbgGLLTaABioi2YsC8pMsGftKmSa/8rJXy0njl2ZrACKH
VZht00T9/xkmPvqjQU70YEcoBsY92b3blwbXGiablTFniyBoMb4l7Ijowxh6
jXe+vFuZ5chQs+FLPy4UsMBYtHyl3OIibGhELaFhNWxn10bmN4Ca/Mmi/cVb
0SbnOnZab8xh2GAyOot4bzTWJPA67p745petqFSA0xBdj68e+SwassWx41OV
qWh6f/vXeWhUIMEP9lrpaLqYZJ1Uw2Ytbtklv3rbfbgAiVIcjvIEecSm6/g7
ACowYAWAmfBdfsZjbVczLpqAQU2tVG6QSKHbghKfIOLU4IaBZTsoiVwy2YNI
5M0QH3s10uBpVLsL52DCexdGrxIO+JRRT6OehvfwOHVmsgjzAi2jMnMcTmjb
JzQArYA4gZYvNqwbS1xw/EmQ9zh6ubDAG54/ODiu0iQ5IMt6cQk4jtHmXxbq
rCx/+VGt1wb4z4rQRX3vki/kn02Uf7/0j4+3fxKlEU8zZ+sct2mvUNE0n8de
iWMiQNObTZLWiyfEAAnvD+3h9ARTRSPQsoDWJZLwBfI/eD+rAdSUWkyQ9Vfl
QJv4j1vJvwuP6Uj5oOYQDo9bonMeY21WJ+J4XPROV5YWZpBEQ+p2FeWF1Stb
gx0mjxE+94pg2aS7be0vE1CLfyW66lX4YNBVa0m8DJgrQS029dv8M1L8PN1C
boGgVMw3eK6A+gMEfnXbL8DEfe34nHlVvdAK7MxZspDXRM4v0IagIB5dR0Ej
Smu1XkTTfPA6iTUYre4/V6XDzaad866+TXtShu2c2bS+VaSpubjpxA/42QBS
/gxlpa81Ft9VhXC1LvesYwwejUvRmgzj6a4utqS/zdCA0a8drjxKSaEmBkAg
Ryhrl86z++BhqmpEvbX8Ceih6ytnU84ajHiFC3JMJkoqZpov5DuMASBqdodg
x7gimpRk67BgN13zKyG39VA7D0Tj/I3byYZFGty/L6RuLBsX28J6InZOrcOS
n7Lj1nSTKoQTCOOVNa2USrkam7FUpeyQTE1gLRYhBa0eVDTGepbMDYE/GeXc
bpxGuqhlvm8dP4EnOIgjZuAgPDo8sjJnX5jnfcTXsA24zMTV9pIK668f9OIT
frANPHvd6ARCbHLFcgMixmQaTL2iQLEXjDVQ9ROIlH8GqEqXqtzcqZQThzYW
aHdDW8yYAdsqYoDuEMuIshoTc3gP6qT+KBqA7pkX8/jd7nMc1h04CODZfgpI
gIByvfe3qdz7lQtWcuhILOzu+KKHV6Di0V68wo7P5RhC61V7mKlhuKzjVChh
mFNdmLM/wQTgiVWAmPkztlpNpGckdqda9OuFVcPgP3DNqUt6QZIwQtglBSQE
5zItajL7s0vUIw8ogfHSKzXfs3VlGOUgLLu+Ri6Q95+uL2ya8GJd/duDYnQL
q4GcsoOEARm7C8uKt2wnzTgecOki/b1bGPfi4mUDlxqyUc48itXb9rQFOjtp
1zpfikwevGj2YzDE0QIW4uhOQqJgrzdQyVuNpIltq6ksxIIGpZpuW3tOa061
sskN/5O7fkDRgXnmvwXAI3bVnqHw1seHgDIX/iKZUtfn7VMzsBVwrscXx/kH
y4aDD3xIYllvh3ANGw02e2WCekqGq0VH4no/FQULuqyawC0nl9w53HzhRNxn
t7R8YQcavbOtGjT4CfhFtAsgh4nWv83IoEDODTSUka4KweM2hTPYnTdEABAO
wqvqSS6n04hVt+dO0EcQriHhvZlamYzpij6i37wJbnOOWliAXapkAuesKehF
Gel0ye67oL24ccOBzCWfBzo6otdxsHRzT+QzCIUshsQBFu28LNQDKCEIcLtw
ugpyVIt/sW+Fx7y7iUBFZOlGe2/BQH9a2ZPxVaiZuNL1rmANMLRrHdN7GLip
2IjgA81m59eyZdKKucE57CIQPof9Xok+X9RKysg8ODL3RGjwFiECwvRfm8P2
wY88JWjyT5wBoIFi+6qLmkCkxVX1VZtD8E6oNh0TKJjZjtwlwBDmY5OcGkPu
6w9bU2fmJLjzticd4ZDzjU4lNC5qiAgNJ1XeXu5DgkGBNRuCTg88KTQTsP1K
ySntALe+G3bIJBjc23GGKlpd8n6FhzCSpIJMD8eyuy179R4pSRvUyBInQitk
Ic5/exp1XlWa9RyERC/NMfFwPVo+0ZAWlPfpGxDyV3cjegaYtaafuRT1D1/+
vmdbn6RD54DqwE6ywIZXbKgS7WpBQ3oKF9+uE/+cs0phetcfLXT+zURQBDQo
23C7BHTKDFMbn9SeSPESb2raIVFfF6Ff1O8odyn8KHj29k3gkrMLVWuq0+zT
ieSQ3JnpSntvGUPyou+qRVQuPh4lirmjSoOGFawxriiC1pxdJ6434jogsUiL
ka7hUPFwggJEQnUlsXQZhAFOfYudANceC99oLeVLvqZI4XTXUy/mpkoxv2M3
f9AbdKqpAeWy72ZeCXJ566L7ieI6uszZKCFlwJ205xVTh5N8kGAVW+Tsba3X
x1GLUM46SDeZdrvpiWRllPj6R/eiQXbxNzTHf99xk1j5NYuyunOjgnqI/H5r
KnXY9G8BnFQe1MwTlaEiJghu+z10DQ4+8Ut4pGMUpWsiFilW7TZ0odxHFvRc
BjjAgxCLpwS+0shJq95sPBzbxVPnyfKtRoznBmCSGv6GY4rHb7xFliCANSDb
LR8CFWqee5qyKZ2GfeyzGwk7yCNIlPicPggbjE/1dILG/6DtWLWWrWTcO7Gw
cp3KAWo3ocvsFHfTYy9o9T4SEXpZRjdFHTay0irdmhUXemGvaa1Vae3QLnDo
/0cFsxRxkOxUJj7h6buwvP72WUiS4ztVZ1IgDTfKl+pv4aCPfUxYa6zJk7Lv
212l17bRJqciBEaWPHLmWtU6fEO0npIYV2gb1FGoptAMLEhqANjdSic1dJ8f
r2Ysvf+7QwWCBzdZzcXXza1PHn3Fu5qV2hJLgvgF7ieXoLEPwyHwe9n8yZOD
EKfvbvYh2ekxAkG4uCSM1skSbsRXnX2yQzfrfJYdd7vOb7XQbIIO38djRL5l
5qm0xoioajiz7EXsdJuNrWP0jkeWR9AYQ9cXHNVA/dcjey621Xb05LG8bXSK
bvWCx/q+3c8z+Cet7D/q4lfqEPiaeAwBo9GUVQ5lFCg+lVU9AhFQgyZ6wMNT
ZtUznV348VdI9RcYApzP0fdKQV84eCMCpp8lEXxx3hxLucCoj7wS7OCwsEOY
9g590eJbrllWXQO/f1UbDniP8gy3Au2DHRdcDCTuctGvNgLZ5Pw7iYAGWK1L
AUni3ZTDrxjqwQ0lBu8Dl4fWQxXKkn9DfPNCnoqG9jSR8nWi/E+tvnPAsRe0
PRBhZ/9Q17xat1/WtMCrOS6E8pkA62vQoN90Wl92OXRwEU9WIAnExOLgwSaW
32+qhKLLd0aipUDj7kC0wGhXf1qoyufTc/4txFc83Y2aWOvgPNwBRYk4euK3
ZQsZ7oJYaAIkOVtdANAV6s5BynWY6sCqrQ4QVTrUiB8XVAT0ros4ATfeRwoa
wDwnOTY/66tp5Qg+dVxTZ91YDKiBCrhunnuzqmekGlc303XX6Bfz/mxvXRBC
iZowUn6M8+XvynZVX6AWnSjoS8eYW5DcZzGk84wDbqnPU+xzV79bKS5Y4h3T
a0GKxe/m1S7kp5wUV6qpVECsXc4/zfou1X57bABJ3IS5smMeXFFK8tjZLdfS
Sx8hKpcKopmadOGWcUfTUlGHNtrjT36nWTNjM/xrWJWOza+/BLopmfIBIJrW
0fpnI1uY3zS3xhPz1B1yH7dz9ib12LfvtqdYita9Wz41K3xI7n4hDkBbepzN
5CpXwVBHkk4wx5f50kGqOz+42fU4l98BbL0mEEJZjqXWmbPY4E3BCVCZkREv
47dvpUGjryZ8dCBSmzR35cJPcA+j5rJYeXfqOZSo/2Xxhe3tyi2IACIyKU8O
DOBGx09Xz0V54tZLclLosdXGy7Bf+8o7UTh4M0olfzoLaVQnUKhhJ+w6BdVN
8UCrRw2HG2I1wabxFqXMQ8bg2+ETTtm+Wlt2iU9PdUkMthN/gHcs3+Ws0X0b
dAyUN5Tc8S1UrFVNAyfMz8n46BzPCEyWdLsyeURcDv+yV1bL+fhaLU0Ldnlh
crrQLR94azqf5vSTxxLR/I4ClkCxPG7l2+gWTq2NVa2kFY7rZ2BbN6BYNckm
7EPXbKSBch7umAIgNicaxtq/a1CB3WAcxCIbOaFb4QQ6DgjXo339k+DTYf6F
srh8SQZXqoVwCP2GQA9tMPEdGd9RG6Mp3ovef4gl44SWpwY7U5zyxKzda79v
z/922bV4OAenumGlXs3ENPGrkPEXW1WH0ym0gOMVghkHf7ZYPgRcXvFid/Nv
hXjKfbnApagrqWWFta0ki/XKoPkG0j4pBn5D/rhjxhRfSe+HVW8TyjPHPUfg
LjUoPl9OYZuqAEy+LrdTFHRyCJM1wUtLtTYu8ZsvTWM9I8O7bCm290SVLaeY
IDb3q+xJd3d1aqcNssnMpdgSHjf3RhP9wzH2PY4cI5/SvV5Zj2CKmVTCOUPm
Qn6+zxUScq0nrkzT+xsIvz7vjrpYYvqjgfj+WIl/5Wj1wQHksrWO6LN7UYDf
xbPO63PUGFbXf579Dwe3iSY3B/jO0e9dYYsKj05qbfjDAba7vXg5SM6kuUUq
zuu0BILBqme6YrsE/pciKojP8k8hvYXwtKBxfGkl8vkjmy44BHkAP0vEPGTS
v4IHIjx1YOeRrFGCdhATRnsbkKWFqTyYhIPq9PewUR2vTEBSZCcNCqjXNcKA
+JebtL+SKOaxgcBWQgIJaE1x5jeDHvgJGRiK7nEurjCaYGVIjAXrvaea78cX
rqq6HHnc5QJMCNvLaManRnhu3CabZrYLm626MEEHyPpgezJIB9L5BJwnSh0H
JE25Xb+ixnj0eH5dNk9Njy1codwrbkLPRoGY84zfYJQJU22C3g2gvwKhiFjp
UAZbyH49by4loO7VbscNZPGj8NVVzNJTQCvbbGapT0gBvAUi7BlT6zMpJqwB
f/TlxQoZQz2EpiXYFVGiwhJJ01KpTwAKuyzLi9OwxAYpgCsBUXq4/u2477VQ
OxH46x2b/XiPrL6R173MbFxmVU4K8284Otn+2SI8ptLe1+4+OD3GX6OzZsa9
5Tzhq0A5fEk5OdqwqpHIQG+s4qN+FZPKi9NZaLB18/TfAkLYJ4KkT2oKnv2l
/CSlLkCBnmXEAtAs7cXR7Lnm5OAVSzOiLAE5bVznUrjY0H+xRnmO8dErHvUE
LCKJh79GmY0QXhJWFt4S3aeqgkeawdP+yVhhn0khQ4Msbw/pqJ/Zyp+nqKOm
Do1napVitZP0Vfm1wVYaLi/QEDtebJgPuj3sA846VpfzXJeeVvBhuSfIrLP8
nlPx3waHQBRTqgsk8o55byGBpBiiTJgiVhZ+6lbd9uG2CFqM0Pep8u+qqPDE
i4iRL6ECSpDZBi3W4qApSLIvjTY596P07f9fT4fJuFdNF2j0nbg3JZneK8yD
QRYoYZemeegDWJhcLmOcwqWjiY8v5c3kKJ4Xhck4JcbAsD8cyHdNA2Rd+OCe
XCwN8MqzEFUac1NaQr9K3JY7uGNN3Xg8F1IG045hH+3GDU/pPgME+rhCH9Es
dqhL/QAXAqqb/1Bl//u/FeZE52Cp3ERQMX2i2vQi9Rhe0BKf6ZR08V7/ZtIb
5dZpVFo4KOxvwkafB0yTPIi50F+Y7MZYaxe+VRjIZlUfbwmUFviqisl2qiZA
MefWqaHPQBXiFRtnlTBQtqyMMNGNHdbOfVFXQIfjjFEWlsRpBjNexqxC9hjh
/kcFPgw4f4V/6oFYYqYU0qO1mcvoygmK90w+vSjXAfcjfCVcAIiaY+20nqTT
d2LapewsFim/lNbnvwpH+i25Bp8/aW6FR4Ba4sv4OXVwQUz6UvSUddfeF8gU
8S5uclsqfyphwLwrceQZKFTpQf6iHsMs6RkBlOSR9ixLEs46Bi0ImZjQDWG+
b1voA2aPRK55N4Ym+HF9pY9lzNj7rUgCBSpffc3vHXTkIXuc/NNfWeytK1pb
20lmj5QVICxrALfQ5aO0XKgwncw5IcDcKXiIgUpvE82Guf05BJKdYxnp3dh3
fKXzivYovmfb4Qsu6XF+kAyK9jWLwswAyPga4+AMwztSJd9Oq5cBVn61/GpK
icPp71I4t+HTtsew+KavnMRCV1pAUZQvfLg11OzobEZ1Fsfss1StV67ZDxwt
dTkudqppwHGqYbRso8ihddTDLOHgRLylR6uV/BR3EU6C6646Aww8F9XdpnDg
ZbduwM/3Rip4xTDxkjW32DsKFEqYsYiL9m1RXZep8I8aaGckzKCMNicaqG8k
s9L9h3X13mtl0TtOKe3wfLHcpyDd0WV8IbSw84GlHgj3xzKaq2Fs9HmnFwHV
BLjka5NbuGwE0j5byppE02FGTmX5vlit37/BBY7gux8662X9w6iqmuimkv/N
xaswamaE0A7a6Wa35km9aDeH+Mvo5mBXWf27y5iGQwGryNGmBZdJAdUywoxi
xe94B84iq2sWfvbpDeJEIUgN8no/H8pjQjQVdY6nMbfUsM7OR93Oy5PA0SfV
A5MylKvvdtV0V8FyI+ZW25oxJskd3g86aiaanHNFuO+5k9HqAUTbj0i5AA90
MBjM06iCC6SiSHpsK7n+Tex1729sg0XzNz1o16sXiX8V3mtDQu9vNtSVKPx0
eZ+kiHyfPXsMSLOF8X44NaA0SmklUOSoYi9p8h2m/UlRQcxSHBhpmSvfReiv
FtXN+zMFKnJVg8ipaiwL0bavayhabncMxQ6MaGExl4QN8fMhinbFyfMQkbZT
6p43ueBUVLI7cuVcygudRM69FdpOG8CZyDmEOmJr0y/Dj2u8xmS1IBtiQw/e
c1t3hIYObOTtyEIbvfoJRXy/RK3BpUEgoWZIS+bIdADV3WWZ7YCT2PLEBJVl
hEpT9QCBcR4xBv1DVPnX/Opr0wsKkBROAaHZtISmxXAbg45SAPndXYw62+st
hh9vMdjHTAsJ44r2YyWwrfj9mjnH2tyqpRjxQ3XOAGkt5XQ/qezQps9OOogX
Qf6IRj4587M1sY1pyhp0HTCt9Y19Y57tPVnRvsKf+MiXolSRkWuTvM1wUcn4
mWQRCMGs68Rp75ljDJaFplFRk60yuZ+Yu5yBtVZVM/wpARoKhz1KujdYkVu7
50mgiZN0FfzyBBMB9X85cgoPAp7dMw1/Mm9jB85uZyIfXGaZY//IIZMNdmHe
5OgdjnnI7ZgMLAKkrwkdV2rzadxbgxqapfkxFiZlHKNy8V/h2wVypedeqJqv
we29N3Bs+q1R8h4Xp7hEuB1fjLskfBjAtifdFp+BS82MyOqKtC/SafcFCkLu
Z3hMTiQ/fzlsQzzdBy398teOo169FH2pEMJOK3x4EGV7WT8QjDuusNsd2pxm
RAitd1jxzUYqP4crgkhADZMSfklBUdt5WIuxA7tJbpm3V4s9CAT2U/7C0aMe
Jphp4W3vgmwUoXMvRLMPvAQEp23OE0q4Z3VZqbve422vMXUtjDnZAhNDqrUJ
vssurcKYWGWbm1D5XdEsY1EuSaqe4wufK5m92PV4F8/10U0K53Ze+NbDoH2Z
dhtY5/5GMaQ8Ur133ZkqEkOHcragroPz1mMAmSkjLNcduB8msTiKLFZYnotz
e9//nxJCIi3jnXqvFH8qtKiTAxbbGCW2Bu2QswQ8cIuEM7Ie/rsocDOCVQvY
ywaOAhumTxRBX8VmtzBLW0dAP2YFMka4dDBDKmQcMMN7+UpY2WnlZnjicb8Y
Ejc1f/kg+uZEiE5Wvjvz/Fjxt6xeLgCGpH4w1/ZGGlXcJxrPs0pR6cDr5OUJ
sPxy1PGkpkyylCqJUoXfC2K5B3ExFqqJWsFh9Z0e21dmh2cxbfHFBX/PaiFm
wEKMBu/SH7A0DKeN0SnZU8/1XkJ3QeMyhGZEO/La9tky67R9GaOkckmnZXuu
cSFMd8kgJoJiJsK9y8zx9iB2LNKUzbWyddt7ENKHzqc6/sFzJ/aQOKz7FlpL
xGy8KOyBomdfRbp/CPpnG3Q1g5VoepprX0AFipXPZ2BjHtk0xm/ueg1onpg5
A360DZJo/zoyCFVrx6Hc2cNneemm3cBXI0XAncFATyI9M+OfgDcJC81ey4l5
S8aa8vuakT4iMPFju+hfgF2L4sfmZsvcefckahNMlV17tGMmVS1UEveNjm8q
hqjj1M8WQ8Wv0qp8PKgP4+FI+rjITkh0dXdpTaWrEivkrWPNpONQZDrH18Dt
X96avYCb31SOI30sZnMODMSF8uJsggid8PbVHU0jQyqQZ0LlYcprHiwZ+goO
Ok1N8T9BIlJCVFhlyHNCiePyb8SGU0WN5gDzJyy2wYcRddcL+kvAxqQHumzP
o1cUgknfqppMxBvckODllxhmeoHJIBQIusx4xbqAcp+fZTIjTEtZXuky+JsU
Katazeq9TqOwpvDmq0EKc7digwjhjsDu+mzO2lKejWdUU7dF6TelFdKkzDi8
6htPZfow9aYzoJI8nlnqn5EwmUAZGMhg1S/QE94t3MiY/8JAU5d/gllzsg56
MV5D42g36RmtpZK4KQ2shkv8dFc027QszHDalIqSuws5pJPu7E1XpK6rTDBv
YSVG5HahLcEM+E+U1m363C2u49umPcKi/6NlJRMB6ONl+xDmR1lRBxMuRfGW
xGva5V5H5sSR80VzJ1G9Sb+uPOSUNd0zAlb3wM8sVMiJjXf7MoZsZuIwFflK
g8+vREpJeiJGGGoquxt1s7LtFuE9SNUg3XdYzLzx/oMUnsCCzVx41F6EkLwc
lrmJl8ch3unguDuF6Vu8BixRKJ5ePY4lJGdw7JKRFnn6kSo6nLSwGiYximBO
QH1pwubuI4xP0eKKMY3UbTMGa+CMDIANARLCfFLP/xSZROorp1ye49EZMZ7c
qqrguJoP6NnFACH0KjTrPRy1DVcFprDhEeTfkeD192FF2+j34kNe3Q09IjAh
Shkq9iO8Gwa8Strh1lDSVqjCAFHEut2xEQopGkvJtlguwmBvFSzC9hCahOeY
udJvWCN4ySm4J//alhclN3qR5OcLtS69jQqIV7VyBIfiTOQaJYHUvW5yvKkJ
IDR7JMQ8xDhLElZXidqAH7A/l0GNB3VJTJRES19LZNw1FrUSJnPelHwBoVwG
qY6f9QxIfI3sRLxxSuwW3AXWB8oD3VDLOnkEqeiWx9jL2MdU/kiwDLlZZpQl
mpQ/THsuuMUFdPkJkt8m4zntRjjM6QbjeQxYnQv4oyMxQSkT0wdzloqHBhaj
rf1tiaKlOa9bX6MjPh9SM9ERa4GHWtssdQ3GaC8nSEMWc+rbhUTrKCJ4n4xa
rjZWAYmtqiuxf2QtyaHGtOEnxtnjJDpa1oqtv8lKLjYg1rIfOBtIQJY7pb/Q
r/RvHYLeF5mSwjrWhOmQ9AVShs/eJcjYdw43BtK7/bnYQFY5L3Xm13XTNEvQ
j6kB09yvnVfNADX0pbFZ3PboOrlt+AtBlFFZpCki1iQVWYrsz9Co9AnXVr9g
3YDVnGJnTWNwNb5yCBf9bpqRMWdIt+hC5QPAeXFSHzf4odVYO6q5MRNCo7aE
CEZdxu5J6T4PE3x3+rH+ve76sJXdIVqlaRqS2fpWPWixSKEKF2t/TLyL5/MR
TxXTsAcgLjPIwQoK/hbVZDUDKFedAki7rJ6WW0AYFsUrFsUuGeKdJOF/GNDT
5vSKXnioAEf7vSnJ3GRI0VlrEt3YWHo/apmr6MnM4hK+zbByGnlcoLDzMF1T
dEBJAi7OYvuFM4o/5w+sFj4Sd6nzYJevpOWz3MhyuyU0Cx7jAeo9AW/8bfcZ
C9oQwCB2bGIkxNxtRtR94KY4eJkmnojiN5NNgyrAOoRVyuoU2bDz7Dj4nTP2
V3poL+RDHtZplTFoDxMh8WD7Fk/aueF4NX+CWG6kryqQiimO/kdWj0y68jRP
Q/zX2aZAxQusmBGzfZWfH4WWX5YIj7KHnAaw/k+ba6QhaPL2e9EZ3+GIkAza
xjay8wC2Wtbq2i3TqD7+BKamp88L6lBC23qvCl0gi7h108D1pWkaBUfHaATo
hF2JIJmJWQ8B2rMGLzChtN17GXrGo+jLdEqHnvYZuMJNTtdBvFQPkddswTgy
MB1SkS7BJRoPH02P9rOFd/4XMTwEDpPjZlTzd+9Wnfu98IR2TEr16EfPFpL2
rzZyglTmtM7VZsmJXpSkdLbSsNfuXB9g5Zs4PLS4sfDcL+AIk0VuK1pH5Gf3
BHco60A4VnM7Ol4xLkdkbWx1B78EcdS7GNMSMQauAkK6tF+w4m61Q3GtvJkt
3lYoeHpGW6d4aofUQ7CeGFa80bW/ztnPupXnpBwSidwQIHl+aczeVGb5gmQM
DiqdIR8AJStfjb7rzaNdVSFgCCe+NDCQBugNm8O4PZB9r4M4I/zxlTrw3JN+
vPQLpIiFjH4rR+OQD56Ww4Nsv2TxaxEBnOYVfpySUmdwDCP1IbcM7LaqrHFG
3aAGFXUj67IISh2YQ7agASJmmU7ubaMY60ZOc2wedF4dcQiX5OlTREAvtGjy
FLh8DTk69mIl7qOvM31/ebFnCZZZmjZMy38STJCWMqXuH1aFYhtL1HXa7R0a
h64SmQhkj73OEjXY60euaTu46MiQBmuJ4zRPxHeJNs9J2LWDbwR8anEtPDrb
R3lkE27KBcclQWa0d0tg/d+/x9rNFzEfOqyj3Q6bUKNiEhMOTZ9rvokhI+ss
n+1fHk35MZpp90LZdGKvfC6NpW0Qt/+tlbW8reaC3R9uUYVNwnsotTQB88Pe
VYWPhVlZ1NDiK9SWntNArEXjrL1SeGaI1Cpn7CnL7cpIvdRGKo1u/mpthmE0
Aw8w+s5GAxVtRrJols/x12QnNQ/hGfL9GTD8NY8nbEMCWwEgfjMPWk1Y78f0
fZXRwWPmVe55bSp8hylwH8RQr8d9kniamYl0cTw4AwWjk2s6EtX6f2Ki2qOE
Ii1qELFxBixlcp6R1qlt9eYZSbhLk+TJusmN1YqeFGC6EcCMhL4sMBxHHbKt
YYKWmXDGIXdfmX5Tjvp8ioDsTSTJOdJiGMUrtn1Rk3gDmwmK4GgiVlI9jzEk
Aco0HHeUqJraefCArfnW+LRFwBUAlPKmSwM5lBSRYDWCnSWmC47n6W5J1aLT
6ouz3Sis1gb6etRlma2+RGGSXzBKWmSfybCezbYQiOgqHU72amzf7sonI7H6
V7rTg1MSjXFkQTrcraUjeRHu8WeT4oQ8eMN/yFDdyuVyYYtv3q5B2kl+04pQ
HqlMqvUx0RrLDt8BoV/UZPfPlguR6ptOmiMG8MgODlSkurIeSNYdzrVaf34S
hT5yWY4lor+D9ocOQ2M//KglRHhw+N0d2elUtfMKsu5DCCyAtfQPS6du7Rbz
9XhRiN5gDj4C1j/Q0kfM5iRyaDhdD9/VyAfe0ozBC+YAsLUo1i+dz2OfeGbv
qOhu0Yq2yaFMO0KE64RwIknX2h12vQPo8SzSktz6RZOhiOEWFCSo+8bwzF1G
rhjDPZEgjG2tFQv6yem8LMrQWJkGnyQLOSqDiP/Au8aooQKCnZIGAa1bsbuA
nttcuK1xlqgwdr8JCNWVotJPDYu/KOSeTxEZdRbhAtymYvuQSrrJonGteolx
MGVdMXuM8jX7+7VIUxf4J7S3E8QnM02wAsarxBy0mHS39ly0tfRt95H2goPO
G+3InRUwp55OTDF6peT/WQFz55EBdINzicehjBrq82Paahugf7jc4UAzbcNP
WacK3jRcVFL59IwOZRxVGK7lL5afkJGMCY5ffQ7E0fQSpYS58RdHgHCarnA7
BLAUALNy0mhV5a6X1GwKiU/d8EjvKV5uxEKFPBmBJNkG0wwCevL0KDKTMPpG
RKDH6gvx1LCFOzyHzBCG5/XK5sHmVYTvUad+27CVAxCXCEc9xiZcJAOlcYjz
YWCOUeJ4QiuvPuDa7x/215L9WSeVJL80kaUH4mzs8/RHXyuAXjHc3tsg5zLk
V28Yw/il3c36Ue1O9v7Pues3xXLCOy9AxBWOemvePBJ73LO6nnAp1uAmCHYn
IGV/hgHa0hlOCIiwfQ/wnWT9iumk2P239aBcT56qU4MWEYMfCuDlIeK3zQyl
haQoszwRYhwu1XBMePhpDuV0W0ES5N1LX9WM9I8ELBcQY8BEh0bQ13n5I+Zy
iWLQ+cyZSBMKZ7UEZD5AvzyTQc0r6f9p+zG/F8UcLqUnZt0dwcdh2YrISbXl
7E+adaKBT6At7dFvcj4QDPiEew0++FnEsvzw7W7BNqTSPOaufjWUTQLDSsMf
ZSCaxeZm4WFi92GOaa9oyTrAliX2eMEtgLTWGq7YSAas6Aaj5n5u1VKV6B2k
0SasuwqNiZ9Y9hnC4bzMHPET7jdnAtbT1D57EDMmYrNeXKP4bZet38I9wZpX
Dm/l0XkeKjj6a8LSO7E2dCYbNDCNwoeGdz/Qb1ax505YQYoqyS83LkdJcFJk
zjY6bClnkHkHg0DcURYciypjASe/l90UxQ4lWArg5xK0+HLvzHE/jf4DHqnc
Jd0z4rX4ClYkGWlvnpVolM4/zRxH6BIX6m2AEH6liGWU4yqAqJvmkTJB65rT
9tOSDZWOmbzLkO53yCvRw3Q2HE/3RtAA22Gs/0B9nrw2H9FVgKORnVS6fOvl
GWmel46yg/caeTA0BMVUo/wPRR58nVsFI51TPWp3QPags9y1wwhLHd5u4SXV
js7p6GGaSvXaMs7ZAt284qoL9Orgeewm0K7EN6bgDeymfFASocv8C2DdaoEf
W4lJTV4VKvjnAAzKwYLmTaJDt3QV9j5kdnUsVRFeiXVuHgU8uwn50QH5VBCb
b3hrOE1sNWDVCWs8eTm+Ji999Ndl6W+Tw3PetnF+SanYWgEcfQS4AN48Lp9g
agPu+aGGXgrnMdm1wLYU7LX6eV1tCP8i2OcZW2OALBqABMGG/EZm4XRSl2kz
X135mM0mIH6ghEa+SHCFwVLBRQMH8MRERzQkqF5ZWaxfpWu9zlvvlBSmXoJv
oeZyJbcW3ZNgaEXBRrHBbNiihHD25dtA6P9+tHtDF1+A4371U8pANplAl8CM
YuuSIsN4IcrHvHue65lxcytN1wbHICMxE+ZGg0l9EXBitzaXuzVwVIuxUAkE
Z8w4leWFRMSe7kA8xu2OK7LH3+iXIqpEn69BpNza6LrmPfDd5c4j73hLQlDZ
OYmkk4UnkyAWAmv74YxEInKDzFvWsa+Jw8F46PjNcfAfoHr9suO/4F1vJ9PB
r9DCtN35WczdREoXd4BIeejr0zArj5bAYwZibnBTXzlJsMJRg2RdHSxy0pzQ
CS0/8UJeZdfmf06Fb4FHTRevkR/kdluKOz0nnq025FgtByK1fIZekoYV1Qcq
sD1XK/X/DifDVne11LLy/04nsFJFZ3Rwsp4RCBOfEyL3LoS8ulyRA0WW/y1Q
2UTyaafIBwRBNQcTlb4GYskUD4LvOs13snSLYsY4Jm4eU45Ws+lwSZ8TsUkH
U2IHzu9vlmzBZN0WG4GLrZtI6VwBHp40oDTqn7yOu4GxRvfFhlTZxZSFPaOh
bneP5YS2Wx4I8CHB9WX20jU/pe7epY90xIYfaa1FFBK8XgTuvrmD2W3APsbr
KHsvTOBkgkmEgfYNqyB+822YPoPfdtBSuTaKWggfpxGZCnBqJkUTsmUp5T4i
omwCZpJrgxK0KfwxI/WVRLazFeq/nZ4FKC5Ah99HspOYvTf5TgF6o5KNvLpb
lYqxuehxL0QlmskQeXQ2uEq+Zwn0niHGCK68ZWMetFohgvungjuHgTTeCV01
vN8pJZpLKNsZ+dLyVQ67uCovOKJC27KWPJ+QDp7EQntJ6RBDBQnrTYoTrcrB
TCo7w7PjQAas/EzPdokkNBWp4pC98YfGrxRzUeoe2dDS2TTIcZNxZZcE2hKp
AvMBnn617E/ig+mpD4LxBjIO8mYON3M+pwhLjHTNR8OZvkzg826H1drQ4IP7
/oH4eAfe9EZrN7NvCvJqMcEZp2489aCpzXrS5k9aMDc7Mi/hSbAMnEPy3WrR
VwAw62AcE756ki0YpGgS+Zusec3eu+sB0Y3Sh76o9463nFypt3am09M9TF4f
WrYjhtdgU0C5Kt4DLYYw+78aFvK9BmSG92HhugYjiDdw8WfpSQ4IMDLmG0uN
IQ6hDs+oXqoqEzJ57fdx1+qy1luP3x6TboE374yJTRVqloYFEF6QU6fuiRbk
SuV4s0fTyxKJDmhbeaGiqgIXrDCDVxZd/ssbKTmltKPec4Ao4LsR434ud638
xMFbQfBuRU1CSWa0bmK57nFTNYWrK8mlaBdIotw6yHWpS/J+b2kdWtRLMehu
I9+UpYDICUuZs2ff5/eU/qkvjpmLU7ZorgvxE3grDhLA647/zUNk7quO+2Hw
F3VqAuNgufn4cXLl6vw8asLkzCvRcHdPDqLR9qbEv7wxxoiFf0w2OU/Kkye/
cDGvRCazsSQh+m63aM8dDnEsMCvtmy/bJy/NRKcPaqIbuTOo8DvEAWjcGn/T
rRg/XcsZEoYCYF2eTF3NGYnIpl4OCyoXgpIX/l1ZIV0Be9ZR1BVteaVtEhdB
8S0e31PmRIGduvn28Qw6tg3W6/jF6zKnIoN8rBSypz923ogh54wdnzisFEA0
3lBx9IcY9M6H5IhwkloTE+9qMfy5dwkdF6hmidTd95cl0XT4M41F6BhBIAij
Ml6ndpVR1X6i3OH/I1mI6PCfPVgd4Sm8o6LZKdH9ddb5Xs3W3J7Dts92clWg
4yljHDX+xNrJ3VfXOi2FV7MLyyu5pEcwICk7rjGztv2zvhMen4bcIhMYK85E
6dp1cow0jguA3DPOLf3Bri+TXbsbafdNRTo12i48E/wh8i+n3rtjM8Yeiatb
C+yt+y8lzagCCChZruKPlwgLe5Ef94eWe5XttbGQax+S+ItjzGavCKs5klD1
fd9XIL22bmswFKIvLx2zP+qOF9ndq2rwZrbtiCUXffvEz/lMewlnMJMNgnoB
BpeOyeGrsvt4nbY+6E0LkY68jrKsT9hVmSF0xJYtspXY0w9JPDZNYfVxUQJ7
H/2HayXzBLe1GXtM4l9bKgQyHwE/C+DyqM3EMSJPa7KmfYyvy4KOMfq0wjeo
7DZUeWzS1XehesWSf9dDaq78vGP8vBlBi+Xh+idykXrMzM58vqdd0VXZHgJQ
W16KMOCcvHVE1zMIdrpg+C/k6PU9hv7Pefy1so/7+jIxvHsr8MjKgM0aPZAC
tnUb5rYDw4yBzV+U1YDCvNQaKyeaa/ADGevy+c1dd+KQz8H2cCR5LodmdEUL
TsoM8E0sOd6+uR9wasRuI2fS1O4QLAPGv8bYpMuZHA8riUmzHJR4SLxyy7AF
N+SZI5yhFGeOUv+TsvXL5FmLbdu+EKRKpbsBH2miEa/sJsEbln3r86o0/h4l
Abh6P/JUVspumh1ULrc8lYAwv/mfV7np2zkOw2gZzHX2F2gHrgEnO19Jz2Av
9ba7SihfXBpOAnXRSvdPz1oqithxBrfkXu2Zwgz4LADCUl1aqeClAgITVzjx
1WLifHOB+j8bzEp1i1aPqAtXV/R8TauhH3GE98UKJDKIbjE+iQNKy3ZahcJ/
4mnw4AG5aNDPDSqYKM2AazdwM7nlmwS7aV5AyH8DOylknDHf/qpIvXy/KM6N
Hiz8TH+cqG84hY2W0OmzFqm/3CAjMJGtk8hNo8eGDm1YQaMA4ZqF7j4saf6t
y8z9CBAfwNbDGkzuujZpxmwJVJ1kXex3qn/+Ce4Ia5pYsUimIjIjzzWv2vWY
ehGzbO8YGFENwm8x7zlZ9z4l+LYAkEcibLuomCVGqVP2u9E+ry/ZkzCQe/lL
Zc2aJMAw88z5JgdgChj5jdJVkYC2b918hKNNBFRv1AflxG1EV4bl3yl0qu0l
3LNcOsbrGWwCK2jA9fcty/9AM6H5QIzEDwYJ+1jgdUcGExn9f67CRAfY+7gz
R/foAwrhg1xuKYNYG6+BPWLbUz4ihFAwIQpwd9IWlqweyGcGfG4pA3M2gqri
dnIptLgZ/I/AmYV7vExeFVsSbH1nouw75pG70OmdsP4Xzi/Pt+9omn6XVtj3
6gZJpZ1m/KNVjOh88beIjm25+QLBWOToQa+2Le8bDuOkDENYs0vNfn2jFfqy
IahgIZd4iCA03yZf7Pvlj9uCzvmaRnpMC7j7FcPhRqvyDQA3rEQrGey4OOTe
n2AQhyty8U+bhnpbXCr3YuaTR9ERSjxFZFmJfwo7MtrKiJOE0c53qC6lBD32
4oIj33ryvKfMadeDpjEmKdJfhvJu2wtmWQpzOxyjqVIyW55/L2Vjim8nM++U
MUZrD/tLCKdEKqTF7xeBU2Um3dxymQlJCndAhjm3j/v7ZOGG/EKaMlP/0v6O
N+CT/v1xBzJJkfExtNHRF7c7yrinBZ/VA+NbzuxVJKc8dQz8jwsuo9SkJAja
08ghz6tzaTyWdWR+nWkbkKqur0emEQqeyF2nVSn6yeRgFNboNyVPCyJDW0qz
mC0hqsSsyD1zxIbz8UPlBEm1smzVBH0ZX8Z78m0mTTFTLor573Ou+ssxD2pb
XzyicvFdZUH3Sk5rJTlZ0a2woauuncRm7UpUrJOEMphDgM/5mXGxoiLzwU46
KWgmWydfHeX+PvEB1Qt0ClNEJcWi4MxP7LMzwLNzM2tIKVoClLcnczHOZHGc
JEnZMUhtRsG1V+8ORAY3r5MjqWHY/rbQfo+ImL2o6mMES3Rj+UpNgXU9c9qs
AMPqLt/Ji7Igm1cYJo59YCNPzgvBhVne/FXzsWGKOv6AKMKpL0RCl7ugIDef
ZHF9+o7wOtSXQtxAMjjTGGtdpz4HbRxANhPr1qy/eJDNbXn97KioFoOvCVBp
fBloeonK6KO9QjQf1tAmvk1SN+RTqPc57FspEfdfZspAVNkI6HdH8h39Y6ra
nhdHflFh77W04FUyn3p8bTp4Fk150C67pgoW083SR81AoQ10AfaD8OToHfXd
3gAqbhB96vVy5sO6skEj36soQb+VdZJjBuPkTxnkvGXDUQXCB19GIwX8Ohac
sug/xnSnQbtRdC7c4Cw1bPvakMeWAyltjRrSLjwMqBrZNb6OqRI4REMH8dU/
5M6JycVusoo8qmbi1thjWK+FAdpSvCWNyGoIh+MFkuioLsL0tuENnjWln1+j
YUx1HjCnBsVE3AB1hDV2NjxMaPokYcXOZpcfiZVc5U+HnmC/Yj0Z4rLQ8BNs
LbSDqRWRpQFElgcrkkGg4/cRgVWr1tyC+4zed/y4d4OQNO8f5plDI9izXuEX
hXP8iSvV+ANZd7y5t+Qg7MKvAmxertD8v1Ye6MChfF1HAHfueqzxhYSya7So
r3TObm+n332B4EcN8aH4c+CQMyJ6MOTzEnVbwHRSdqsNsFrE6wVDzq8GFycZ
QEoaBRndePEPHDvppLH5XSywgz/+kr4UPWSZAwkhKF1+GyWp2gjOX8Ix7NHj
mKsPSNJgkWdaH5bxIj9ivpvirOh57edaQ/kUJv/6P2rTXCDMBxIbYsYtblGA
ZsCN2sV4ZgqU2tPE/2CeVQm8Pu+lK4K9+3Jv+e740WDKIu6leazrglMHftZm
t09R0mAvkg3+Mxnio4N+B1IT/cSEnSsPxY0ro7PIUjYfEjF0qhfG+ev8EpIX
zq73ozKJSJfwh2EIiLr6Tyizvbg9ZDEfCJ9ojpbvPMSqTduFv955YR/YIl7T
sWJnanIkCP1Bs07YNpeXhUq+rxJ643QphZtwU8/dg3OfteSQbizvE2Eq52Ua
EDcaohJJodBo3Y+eM7Ku9KxrbxvSNk2OSkd5RAQfZHv89b/+J3BM+l+U3coH
x/SBMCdkKAHDgibzHk0IvjvWGdx/zS7oLI63tl95Bq7Z5H8pKBc1DqYnE0hk
rY+vt6dhWjWuWQ387om3oSM/pLsBJV6o4gq5dD0PbQYmrruXhyBbzor2v4cO
UhF08W9dLws5RLqYbix/Lh9v1ckr8bTrv3G8nQArZ+zkBNTP5bWqL/ufOMvS
dI+72Vy7f20sXjp0noi2BaJefHkn29nUlO+NGSbWRi4QG0LDDiAY673A+dLm
VLO0YQQ1RudymbNpGeiTZS915aDj+z1/Gw01Wv9pFO9cygkpfP+lyIPak0Hu
mQ5z3yppXkr4JRVvxT18QS0dQi3INc82nBVwRyyRLNqvGInTU3lQq5fbdYtb
IvwMoAFJjEsDH8X/960gIWPK2S1uj6sCQNB4wZwG0gxfPOQGv7i4YrCQOFDH
2bWKjmR1KjANieXusgBHH1SmY00l5Iz4gXGOWoJMaaUDQX5K/IJZsdanvAMR
S3QnY0kOnDcqgQj3a25Io+jahn/MfvqtcLhcXODPmkr9BypNtvjidAjPEjQe
Bn5ahOu7wk70OoCMlIC6zTI5yoZqJFGufFS1MFiz2dFbBp0w1qiAIrIbIKT9
9kZDlvXlUUZWkBRyJi2vC267ne7jLb5MBmj6q6gmiJUYK3GJmsJwEQInSiyJ
hgtamTgK6EgdGFcJ8c84/WANjB1KZUjuPDiVny4GtWIGPszE0QzJDVsPeJun
DiTXLPX5ez+2E7pEheX6SY1fzkaMZlBUPGsAD81mU52ilDGz8Ztm5y2r4TLq
3TtbsAeGwNcXcvnkWwHiOH0/YLiwerZCR4Omzp7OVlFb/YDifYkPGTGAc5+F
j2LOSZtNcfnKAqCQtG3D8eu2ZKEWdjImQVaDzVA/RLwo0so3PA0MNurGRcHj
H3EsC/5ZgNxQ7IlA8/yn/YYuRPyQjs8heuTfRxLH0O4i9pd6cxPE+4cfApn3
81xNCsxeaoiOd6nME+TPRs1DTEXxXQko0ZLOa3rEddIQxHBgMBxLS4KIV9do
wOz+tkceJj8sf9rt1QKwsiYNDvWR+Ih24h/h6mKnNeHRnkt47iTL7+oBQJ3G
CllfCn7cEkPYqB7U5dwCNFUehDQuC1w6nEep93p++De+bNaDnvFJ4pRgmf3m
etsKb2p+/6jP2a8Xw/FTnLjZyxzHDWuee/LzNLD9oeIDlOZKdtksJ/Ut0JgV
Z/aMSvuzRAIMFNVnF7QPqQHCghFyO5PL0HY4SXnJdIj0zpBM/7qruiPW6Jij
0bNIdUlwjNWf8mG5CmO7eYC5te1pkhQ6N0+lPlRzIbHgEcHg0MTp7sr76fXp
0g5Em3j4ZBc6SlqtB3qrWHrMYHAXC8HE0vpYI5fk1KxuT7vSDJ9QCGR8rN6n
4+9Kn/zd/sWxDlJo4hQtVQrlDy9EWDUruEAQP0sxlt5YeMjywt9WQTpi2nWD
yBmZ4TIFhd2rYNRClIYKYYRoaE+z9xVxiOCjZo015h3n+V5guZnm/md5IYcB
6zRQqMCvIEG8fd+27Kq69w3eHrsuS5BZdWvmOfLmMbOXNmzQFFGBwm/Cg5Rg
n2M4OZb+mhFsH7UCj5y/MWD4XKigFxoV2fWPq184cKLEjc8qBXyLH4H3sdt/
S4pQWg4r+D9M27RnnAgmeL2e9bbZbqx3Hn1EWske7XlMLNGVGeuPDmAERRu9
iRGC5QO8qX8ApGlBe+u2e+T0CeIxAb2mnPS0A6hdnNdekiKE89MtEOgLlEEX
IeQoNY2IUtGKL2/d4SY4XRRs4D55+Sms/vyd54vUOxlXYtmzvQWHAYLhMqDG
511jvdJ/dbycE/scUcx2ns2q1Pct5egK1033crxiRrCUA427MAFk4uo0jrSn
D/2lkmEslENVLhbOl+VWjnGxalkboUG08l8Q7h4Q7rphAhtU0PbmQDjt0SAq
EyWGpy/V4qQBwHO0ydoDASriVeq64rR0+devmXGoZkpq/iqIgLceObzs5604
71Vn8NSBuONb7+sIHiDXRsyStanwUZnB+X8gOGv9aXHD7HJHbfLPC4rcfDyK
e0oK8XWfHm3o8dl5/AHSpgDr6WUqf6XJwyIXMUVcjV9O+k3xQV/I/XjGdj5q
MjUYwEatZQ73EQd4qUrU8uYFipCq6KNzy2B6LescB35ydWL/u5E80AoGtwvb
+wL1x+82CMD8iVJEPoc+CZ7GL+C4qw61hKJuphnyQ+spjJK/a8dtu8N/UoKc
bhY5THlG2F7Zoy4UJoFbkKOWQfw0O8WpRY0ac5XpeEFScGkP8vMpJ98NyRd+
zACGaH7HOV2znK07QVVJEUwcJuK6R6yI23j9tOv5OLjo3lXnT/RiNoMD87j2
QdffetHn+PmVx3VTYhIB3wKl23x0FoK6PdY7bESm8OgNNmkxP2R2VWAOvS2E
eWflutxN6mBq5+O5LjyFdl4mC789hVD+C5tgnvKTgL8P/Da45fBTxMxL+MiV
ZrqUuTQIkTzAnps8UuT2ulCYogypbk/NCXMMmN0LoC1rbn0wIL+AIXmVbW6+
tj/9NA7wT1tPkF2JIVznDwX1RHUAtBBy41eJlzCN6TccTfBQAz6EYhzJVLrG
+3LYObexsHlPMJaSP5DZ0y+W+SfAs7hbRa7IxT8Sx6Xsj07NV+RSxA9mmEcW
rC9Thfan+zCBiaLTzhkmkuqeUbS/FRgZI16z+qDMWwf7iI3VKmnRNHfkfmSC
bxK38w8c5DxDx587THia2tsuFdgsLIAgghxzSGIMnwI/Fj+T8tKHlM6HaufO
9RJZ8ePtnbfJKNz4fgsnxiIkiSY5RgC1sZkHBCGsy7xvFv8BRF/kVR1sLKj/
QBr2L0gyREbtGfzjmiAEZkbNmJ2CimApRUG7diQQhb4N/JKwMm7VDSLmlAlY
T40cJa5+ByJgEvbr9hGcL9cPsMT+OCWIyx95FtLuBrmif9xSO9Fyg/2p5MUu
gQZTa+9wVImSozixXZLo/RPqsaUtBq06LLimNfoysFb6BpmY5l4Qpjv90n9V
tY/A1D5FPOURWNh1dYxDILW9kJAJIyCuJRC2EVJbPOjdqO+X+lS6NXMFe6ER
AZJ/3j+s7ofrJNx61U58IZJBUJqTcJdWyaq5YUuSa8mWcz/XiejneEdAoLAb
/W3pm+JLSTFyd1cH64Krsk5jG6h2L+vfIiBnJ0faLKjt4clxZjAEQ/QTbTk5
8FXHrhLMpMI8+oepyWcu8pawo0BDW3zn75T1FZEwB20BRQAM0edfjMWaaxdn
ZcVPKR69C2Fa/FFgf+Q71HmqfnKzH0bE9/dwjCTiNMKi00a9hUk2yOG/81DU
kU3ZrBfFd+tNg5z1aw5QKuYqjB1dTV5ViJxy+6ITvQP9BGiOwql0uLvWow4w
SdifmN8LHsUijuq2UYST7l0LWCL+Dgl1lh+DNyvlsIP9uOuJ9QGBYKKOvawZ
Fdo/uQl5RFY9h3SgGZUkHY0mLbWQZZomGdGyYK/Nm2HAMkFoobksrzRd8ENl
YyquQmlzZCQ+gUJEKtLHwO8mbhoyJFOmXA891S4hLfEIxUzN93Z/rNRzFVf8
yHzBBjoP4B76fujwzsIJrMET3+YXps467jtpqhij/v1mqU66XDrVyB5kihIQ
lQivx5ctFBmQQQedwbhVLxh3jbtmc9EKPj3HA9Iv8yJuDhZw0+8elgwSQC6U
D4CQK2JcJMOcxhYf0zp80EQCHsbZSaLOyhK8diLuZvdABGoiopdbxPb5n1is
y6zWiYPOGAmd5X3bz8IACHgZIK0BolpQTQm/V8pafZXg48TIe3AQgnh+3EW0
2z7hCtyeVLP/YwKv7HSeYvhjKUZIdHHTgjLDx51yuCymsfSoTJ0amVYM/3+N
lI9w8p42XRJr8sfoQ2XuGWGl0MKdAAH+5iZbkvWrNHpaK1ys/SRSM4x3ZzFg
gCSqWQxzXixTdCVZ6ICi+z28vDHANT+D8tstUu6tOjxZ5wzIZ+cNDFLhH+zr
pRf2L9ukGGvnFsHmLkeF7pRp91VYq4YUDSTpNhMK9xFWy4oBVc6GMnJrVof1
jtSQhyEw6ib708YYl6nhT5MW4DzrJbkXl32h6Z/2OtpCyPO4CLZ/SkhMXcTg
70CxqHVGXvL+m7fIsFSkJwD1pjH179JVdb70WN/ulsd5iPkMbId2Ugew4A8b
Gq01LAbe6/u5F1EWOHq5sTVztWdLXSEj0Pqh3KL1mBxXEZR95KKFKgYv7IE8
D1VCvUX/s7hUZlBs5wH+pEZPQpvgOkWBzaQgiGrViTxxxDY9hlRN05C/g1v4
/m7mxsBFs6ZBEZVEwR8sUDRAflFgjZYs+ivbr4gLir2Up0PajmGQZNm4YGg8
X2w7dILPVKSKOf0rzX7jeaLvWqXqSXvEmNH9ogYw/IzHms/X8stvYP/xILdy
ybRF6Vebu+RsLhYYpQSy6c2GAyxbB0+ocesovuDq+X/7TL/B0xaMuKZAhn4F
Ers3aDaQsrweRvFwoihK3/jywQLk8oRgz2UfSL9GcIwvBNtx9SXYUXxBJ3tZ
pXUoAI2Dn/8aJkdeG72/ZiutcfOtLuZZUSHxCe9/bStbbqv7JXgH8JnNZRTR
QilTIP/2ZASbFYV+LoPK4tsdqOic+f31wMSrDeXnULWuDo3A3wWx6hACkr6A
5jlsIzWJTWk4YM2NaFs7tHe5xc3a0l7tfJqK8drBFdO17dnCzFm11jkSYBAy
UhmWsutoksp2QEufr7hWpfjirubHyMdt0hx2/v1Mw23Ad4yJDYRlSYf4Sjfj
enZVx8hSkxvdvD2Jqh4QBecKxBWUevZCn4HDXfTCAuM3+WKNjbFBbhnEtSbU
zogM3D6MAOZfmhZNxyZ4ObeIXxJAW5mw8yeds3oFVCD++jsDTtROw/Tqh1Dc
CQ28ayDzyxzGT1wnqlNNrRpIc3R29OiovKQ6osbKDRXqt+yagF8HeyKEux/6
zK8DoioyA0N0fA24DA5xpb7//gCpa6X6jALUXu0Zlb2F6Rs9Oo+vefa+3oXH
h+Z6I6bsOYiWuxeEcNdAO2Dgc+LsV38f9gULcXFeVhZGdmvAzd/1cngO22R2
cB7sQPGB4Xx/gVDYKG3m8Eh7C99AdKFHCBj6uaH+Nl7mAGZvTLz1TRhTNeL0
9rdFO3ps6WARIcFVHpHqYaAGaVp8p6CEWWJqnNA59Jds3hoXibTSQzHpphqV
QvIdhZc+g9KYSSSFoOTyY6uLIw5d0oAco+KrNjiM9zwiDV/uzLZuG3HQ3DSB
Pi4DcC8+QdrNLvNZjwXlqPyiJFiZa4tZyofrQsCUIbfSwIG6wF8VzbRfmugY
1BlFtMQBh/qnYXowlVne9dJw+AP0djIpcdoHUemvjA+isjjPi5DP5PxNBkcU
7uS10rJD8mnhLbq50GEoLkwgn33rJ5QeG2FREb21yaGZ4duQslwPPaoU8mZT
50sI7aRP4fCCwYBBU83aJDBE5881r1ZWPCDAMEHkQpen96SypbEG3wPSJfHA
6HnwZd6mFUwNFV+LLhJuCcqX2zJjE3Oj6Jws+BJjIfcwNSCLjrFi6WECCGBc
57FxhX/goVPWLAGWFNETAJgryqvSGBxWrM9kzv2ECvBByso9TvaIGdyRixsQ
RapPjXIuOnUXnT0CGPQUS+rn29apoaX2iVe8STynI56OfJ6nvp73tk7A2L17
KLM5phhUAr5klMQt8FbZF6WBnrf8ungJ4tjbXVkwZW1JMN+VPK3aphU+37GS
AwaizFJ0S9F9JjFMkXmQcQjbkAMEa7nfA1BTtGQwLoLIX+qrkWq/CW0r1KEP
cwRMP5pe0sFzpUexla4diK0WY6jfZmGMaJf0DFit6CwW5iKiFqS85bhadQAO
GBhMcL2o3PfqdEXL2yM87pOaq5aP0nZSY93WIR9kjYbJI2Sbdc765vrWEmFZ
WztBPrQzBPAYeEJh2UNCL3qjFQiqOOV3xlPK8+xBM5+n/edYxmjgB2ApnX+f
gHZLK1RQv4dZqaE0bbf8tx+ueej8D7LmJbC2AYuKYXQWB2igobOgSItbrtIT
tb+2tTT30HC39KvYXx4Dyzf++x3GcYUwSP1OuZMRgbpewTUKCaVE4PGaTR7g
AOieESx38hLP1nhQ4RdACNnmyi3lFBf6ylkKzj2igFc0TH+WOMs3V/Cz6Ehi
qDLD7CPVU66QIKUDxRC0PqBjw0aOer6o17XbvVZnjFqanB0mtRXDIinEUOxD
vaRsLDIM0a/KVxz98J6nhwpbHICD2SagMkkXzkNCXAPzUagvKNAYMbFY56qB
AIA+EA8D1G2eKdY+3TxyJRE3qOsNgw0UikOEtfsf2zpHNyaG1UwS52PpaMq5
KAxyQBPoJ9QdyUq5xU/somE37PV1wBtA30pZWzv91efU1No5/HSp08KhuTyU
To+uLHK4wgbKqeArtGFV8LP4S+Sx72Ms1Y3nmBo9dqOgccbBLyPptBsddzLE
6fYGBDCSHFsk7MZGJR0SGVXMS8gQfeieTjdE2cjJl1Pyau8nvRqUNrWKI/uj
1m9DFG72rMBleIo91LaJNFo8CC3JB2YxW8NbdLs9s+XFQQ2muQy1G7lT1+Ch
IRBNZ8NlgmcWJgSPFDehpnuTG4nr42iMEP+KpOAK3hANlqtP2b75g92UewFr
tcbyOOfoIC1SLszgT5kbS1BZ7WosGJr1wqvt1IEmM255Q2VWs46O7VgvWvWg
YxIHZQWWY5KdpV3zF9EtM1rHS7By3maufPEh89G+hCvxnFdI1MnMgFxYyRBB
jMEF78+RgxovmsGYqyE1wc3cBV44POMMmI71j8lGafw+6wRToesg1dNDGBHG
iC8GEzqK32IFhbYClVP1t06t3vX9KIy8S0ELU2khcMbTV37KebpWTDW8DrEP
7ssS9Uu67nNx6QmcHashjar60/tTgMQME0nWMOEqbYnX07Db+QIgc6v+po9q
epV3dng4qfgFYE4uuyHKFN4h+fVR24US5dk7m9r2C+r3w8aI3efYxa6Cj902
rDMy0ljOwCSjvIAsdcobeI/+aiN+b+nLpnroBKYfWWuEXLhRu68HMMm59Juj
QaiQzHXFu3TmL4pw916wDJkHwzfRSFbasWDPOPcJ00j27gnz2XxYoyXlF2aS
5StBUWA6ZH/UGxhj+C7M6PYwJyAZwR2h8zGab+PeaW4MXcDUw467+L0THmwW
uOgVQc5eZHkYLlj8NPJ5M7OzlOjdimMAxbCfUMP1Cps7PZhb5oqC0vQ9VcPE
CxjXa4fFsROeW2ZkeQsG6udNlVDP2h9SELRNybdP3PnUT1yeVOOrWffjS/J1
pzBdYjgnpmuGXDmarrqErXOA4VxKUHc69o+jh1oCx2RvRvVsG+c2oI3fWVaU
UcZPgfN9TFDIunfZMplYdTS4zndDhqFBNznQw2drtNwFP9OHkhW1BwyAxYgV
afOkk8yPMr9eGTALxDEWU9bElZs9GQ5LttR8mvTZ5Vja4dh3dLIdIwxpTUEm
8wO8gXV2LSGjATFRhOJt5oSmcRbtwCJGAFk4DOOFwb4/pAxIuhtNZN+D8TC/
vA8KaGLp5WdMs3z2k3d4uPSwRqM+fQVfHUz+LoUFNZhMCIob28nZRHTJnhNd
ax7lxDBS/QNJ0uBL/4RlSbusAgZZapKsF42wZVSh0ENxQH3z7dpPAHMaXL0f
L3DRz3PuUBrWOC73wcSalDN8mTEHm8B62+aVWsdrXrjyJQQHyveIBIYBKe8O
+BZaVoqXs4yG6IE01hMDCP5+lGAzbZC4+iTlmkRTHR2Rk25Duj6fyLIjexuv
JHBlDc8A4w1JGawqJ9vI9B5mCUfmmo2ZvsQxpJ0UuX+fV0RR3hSbKFMTgQFi
7ltz7Q9mqirnMMteM0RFXejspgw5NQQma4KdG6ccdm+qUZDo5yAMk9a3OPil
i7l7TGodKOV8TtICGhlk2qPlpnQJANjE7Fg/yuywQ22tUSwI9tpja3Pa2qNy
rliUNUtM10+tMPAkpBKTLs2k6L5lKLJWwRa40zDliFwwlxiXgsZ0D/fGsFo5
fWVu111ivrpKvBzdEjwkaouGRkQpUrnFd6jhtQT6UarGXQb2Cn1wAGHXEw4Y
cMtaTaIKfluTn/xOxarzk3vMtoNpVI/fokx0qdqiC4ziL6+421HkyIrktFBu
FUglNVDc6PzgxRTffFtvyiHOPz5c0ibY7yTGbojwZVYybZw8CCzCqMTBinPM
3Wdng71DLemKNemzYsiLABB469bQoFM41hMA9+xKYGY+FczdHbWo66fzvHeW
ZWIGrzIxeUTDPv3rjnmx2keqXArE97CUwQ8dHWDce91g2CFR4aNvQemG5P/5
opd92Z3k2Y5FoVxCwtO4vTyF0lzaLD5WttyafglsLl+0Ta4MqamO9JkOPhW8
CTVXgCUiIoMCEg7dBiYzJRxZAvR2qFAYH7kQPhNk9gyfA1jofVscindfntL+
Epye6jUmvlIFQL9Nnct6Wx8WCeDFHHH2bwtkp17TZdo/Xyd3nzUZtcGDCv36
fOEUdwU9dYgcGmf0aALCkrEerfXY5qLjnzwWROciAER6c05KBe35prZb9vug
7aJcQZNQL1kT+jgRripqqttNgW4jtbNgYGMNf2Kib9hTIoNgzhS871tvNxz1
bJhiPkUA3/PhGrLQd59oNASHT5dPnWMLJSqQTWf0/Mwdtnaut9QowVDrVzCW
i8K5qO7bk4Lg35tLn1YsaKJUIAjdl8OAkFFm9I36B91Oz0gcioUyx3Ut7HkM
Ki2gJnrWmwA+2TESZMfwGVj+HHDd/AELBr/CWv/B0mrGc7tCdwO4PLsgIAtp
QYsucRLHbKz3+6rRfPY07bOohObY1clx8+IWxk3xojuN5bvX4Cwu2+yisrem
Hy4rrb06Gw5tuH17+c2oZvbuAUBpHedAXLMmqGVEfLZcaVpLET9gL2t4ml9j
HQAXVHKh2actafIcrJQ1KfOLcvYSJudymv3QMzqDKZ0kM+qbVr5bGFe+n6q+
NWMllHRBQDE/us0saddfHrjKuZJehv2TEedI43x5765zzmJS9KZWshK6nC04
C75lpCHHXPnHcigzgcwwhlhDjilouUyXPoBCIUxgUOPOSsVFbl2Nv+rPdl7n
CeaE9xPh2YCBPTemyeAeEDNSM2k7ROy4bSwgrhqvXgywK31rmtxvp20rsFc3
VkI2hYTLyICHJz3x8QXlomS8irItGUedddNRFdS/6TEFd+a77AsAkB4b7Opw
UjB/85seQQWee02Otpdy7qcuuIo+WR0dNYn5d5LRASAJw2BRb6YktBSQEkXk
AZ5mJTTf7+zUlF1CijdJZ0qFBrTv9X3Xi6yodP2SOAmlam/grSMMhfV3Odgt
3YOfmD6V9irvj1SErAG7gKaVhfFzKBLhuDNnH00zqlHYz8YdaqmWUav89jPD
I4FVOdmWsBfKe1TUexJzaHeVu1vWNjHOyRRDy8kohs8QpCeqHuJ1z0n616Wb
kts3JsWMxnDm5A8W1AFG+NBn8KhaAw9RsERv39QOJQck/0nk3iByLC9n0ZnR
9dOjZUzgRPhtM9qM5rUqTdbZl6uTNkARg8wk37QFV4V2ljnZg7afl1A32AAU
AGQvjlbu6Kmw5osKhEU6e/Ll664CsmPtmlEH3m+qncc+jwDlDu0ogmO/WWcI
kaocZfbPALFdaSPZ6Ul+zd5cuwnkRj9rFG+pUMZKJgld0UBU9qgq3KJa6kyA
DS+z27DczsygQXozYXhp6KG0RZWhS5QhK7puoAsT6pqbaZD4xkcI1Gcdab28
d9TPiqnPi7RWQoyxuZCDTJM36vmAa8KZzsgD0IUAxW+QnfPFk6GxbZOvzv7S
Gw1kLrfoGeoKXevXONZjs2V54X82EQMMBQHcMmzmClnDjvbrjq1xd5lvqlCR
IAiecckzvP2TckbqVeDho9VhsUTPJIJaMefnQy244cTivMsyijFmc5wSg2Kt
55I2nj45wIFMj8FJlMRI8ZcHIcM9LRfViG0z9sNyObH67/mH44QqVUbaBWfc
C8TZqjKWDjCVAsUUHGK7e9dFd+9FBpt0GlJye6MI0HXlsC774fMrrax/ZLDJ
k3xpoffKcJKlAtbQr+7iD4TvpsQR4FrDg5fewQ9r29S0oIGP+IqzlujEkQ0t
s2ofV+lLAYhR1EzOcrESwwS1QxIhZ47Bqf+uMWp6nU8SwpEroyaz1Aowrdvi
gz/NL0HEdWFvtzPaT3ZpKdYQFxqqE9QaCF00t9/Ur1uq/nCBBJkC9nN1YCw+
4GZdce6rT1CEmf1IHNAl6aDFuC1YlLPNtfWNF69AC0Pk5tD/IbSfiyMNtP2s
NTFiwD9lFo71IBV0VV4I9M/KVs0Kky3Q28uL5Otz8zQ2pTiBo/xKElbmvqss
kIQFv85WueOtoCcs2r25TIN6WsLh3/2hRR3eLHXUzVZdRp0IQTPY2g0AR2yX
sgJoZIMjHXR2xabibLa1/MxW3XcR9hRb/JLNZP8pLgTd8ZgthaTNSxCLEttW
csx70KR1HH6vL4fEm9JkIyE1h0ZF4x2l8PvrqulExmL8AxxINlSdlUOJk9o3
ivWr53OjlsWyDWtBWXAVlF/IvBkPhqvyoE72sYyNegshGSCLBg2pCXlg0u56
SXLHLytNOSy7PFO6ZXJUcrcvO9uOx7kVPYo8URWApqSyitexP1Z9Otkyn09a
T5b24o28KObkUIEbxuSlkTlODZcEaecMmXS4aLVQhGofD5fFAzRMilLKSynE
YDRmxhHkjCnSZKQwyyXhAJEuRjebywTGx992v5s0J1V6W8rTjM4DGneaa/Y8
SJ25aUIJuLBmehphirIkwqizR5pXlXYX+cn7Hj0l8O+Tb0O7ubUHf0itkZFB
p5Gl2OlSlU8RI3f+8lAJxQS4hx5splhIatNv3wplYevuUdJv7z5Tf2XL1ndg
BTwrVXT54N6f7VkWsOMLa+XDUwSdfU84XD4Gt5k5n49Mwv/kFFH/fPjoUGvw
fXe4FpHM8bCsHfYUS53niISIMBrjJVtiwK1MkrVh5Vo3iKHh0GQZJFZR8/Ud
yylJW8SRK8o3aY+98L/bU0e5ak+lvHVSFatTs+5f+lQfMS4LLv39lPiA0Pt9
FoyHX677lsUCOhQg/48W7dG/TsFcp9eS+dB07T+G+hfNMfKRr2PPHCyrHhPI
OaJT0qSWir1jL4ukm7xkNYgLUJ1tDCvdj5Lnw/f0wiGDPz6yRdjrYdy1ClVJ
9GYF1mhBiOn3Ysxxliwzis4WRCzmlBuW/heceYSE6z/xC+yRS2jshtRpH5/Q
Z8Q0xjtug3OsncEsdvd6+7x8k+TwMJqIaUjksFu7zWl+PedzWqe59A2odvJ1
+PmlhjU9gcXr+lc/77//v5Th7AdsVgJBfe6pX/oNCVBfAAGdXB3tM5cnSJhX
yMC2K9UcjLxwkt0o15tF9SduRoviDLTbsv6m0iTwoXf50jD9HK+FlyCmQj5r
MM6DNZlw09U6xZat/YH9VRbH2ptW3zq6n3a1SCtPBkWUWZPOh1/TuPm9Jhou
3lV0q2Baq5l/NyrU/uH/M2/JNvvbKsqAp+V4ZyogOMgUj87ffmEU6mbvh17M
h5rbGYOWnlpJde+IntD24uOmFHRo+kRf39la/tAVFnNFjOjrYBb2ZnNwoxQX
aZJLT0l8jTH2Kwss1UdQ2hlxmO0FPjJuaYPfqYUkdMpVnHwG5Qxg9G+6aiNO
Ml5GHgLIFhYrLf40SJW7l0u47xuvfOcqfNDgB5aO+P6qYs/EjZzrwqLUQ1WX
SJdW7bMCEaCi2LYJq++tUT8Mxo8mX78uBMiYyPU/gcydBKsSqwpH3sv4HlnJ
QwZRhqArHiwcjRBkaKk0asPvTkXx7zDwlRGlqhPSvlsHpcfnEIY9nmAXbspz
m/BPqcFHe+fsKmfV0obAzFlzhCasM63pVs2e32hDcRvSkoSeXX2EDh1zusf/
adwCMEBD2oETGM2wT+cmZbNmjnUfdXIf5I7V8ocVbUd87hURTXhZ7xPui1qK
42I82DAFOGRQ565vEcBEG+FicUsfHoOrgeCG44VCdJXeODeqaEQ/dqLFpM29
FRo7NrhDSx8TrOPOWArV62TE/EUiveG02oKw+5vPSl5Gil6BZifPHL4m8G8u
kC0bVVrnhecMazdfKUm1irHkZLeOVK9c7BQ9fYv2P4nlRt0Au07lPz/iQzco
42fWvUa6OkerQsb+xxm0j6JwcHuyycu8gxYDyr6EMsqldnGK27RSMqNKMZO7
4HQhNN70hX08p52tNhrm1xYXZV4tECXhWmQWY/huK/1eO3SZYugf+GUH0ZC+
jMl8Zv4iqez/bSBIXvZ/iBm9gN/HX7Oyf698OIhfOfq22eVvPtW0szJ5yd1Q
hQ+OgrkeShMJoTUxhh+Aqom2kMuKGrVpYD+rOq2HiD0U7n8w5Z7cfslor0Wp
W9Oo8klBWA+FyJuOktmJ9Z3i+9e6PSnpCXmBfxOC6RfblN4Ih0d21qmNWmkL
8tM/KJESGNqXt6pFxTDN4t2Agy8WZUlDI6/c7FQ7YyLbDUHyG2kHuZIZ4Q9H
w/nfNhB3/+KlHmhiFrAA9j5M79Aenw7u6g8p88qO9cXq86maOtHYgNqq4S9e
rCotoyebI5soyz2djh483GI5lUt6qoVmSRATJ1cOk29VBmVa5rWZ0fzjeSir
gHZEi6VmcbxrEDIW9fOvzbQXEPQ4L/ciK7Q6dv8lu/GeadJVBcey+KVRYmDI
w0dL3mnig30BQ83df7H7tXjuHNfU5i2jRxoqVw0Zh7Q7j9iyhImZ8YbklDKs
9Z3CbRnAByMoy4t6/4ct2m7vjZ2EvWq5GLLifUTAGcI2/brJ9iTW1rjiX092
XnbWP+YZOgS0gBmyJzsQSKfvsC3CqFwD4aObgnQtrzFXf4GgQhNuqngGlwSc
UJvP+KNsvWDxt9Cjm2EQDDXhyU0LlyWIgCStzfofVgVA+2EYgRSgLEIYv0dP
0E2m7Ljw0PF1OqXtuvFQkvZNhm5FvBr5rxqOnj4mvj3iq6/++N+FrWzpO03e
dHthUDdfy4w7pbSVHTOOnFFRz3CFai5bHXH0hvRIu7EEpWQs36EEJ/jP/R+j
wGJzh0CUTSHnSmJbfOLIRJmAEoScnAbIncwbeAZAtz6uzWspTIMENzwnSCWN
QFeBEfNu5w1vzYOCgj3SRzl8cN7/pTsUeYsvkQuQM/3XLqnzVX80tjE8xlru
X5WexoGxgHTmFI0p49TtzreGnIPybXsW71vFyfml1PJwOVG6ua+lGTViedXN
mzAmNXfB2kv+lCMC1EyU14OEc1VxbFf4zBNB9jHT2XGinMxBkHxzekwlvDgF
Pk3jb3nEGal7l27TUhTh5i434kjUbZz8/WZIAS9ShUY2obNvHywzFjBn4+X6
nvIEWAIlg8ZrJu9Ruc8w1ZDMHsZ0lOtsxtQfqUo8X/RPxTYqc7Oq8Ut7kgD3
4WXxHC+WJP4EHIVyGn/6+A0U4cQr/0sBFuSQIJ4UiFY2LpYv9Y/PuAD4+YRU
mnyYsKLuj1/YKXAzpu9D7v2Q1Adjpkv3P/a2pV/MtFUosualcyLGvSiydhvF
TMYltGdO+z9aqR/IHkHlvrgmkNkAfIPWjXimpCa3Exh+RptnTemD1FiTUjk7
ALXgI626xPaw1mbcIgce2yWur3ZPROI9Wwnrq8R1WdYQ+kJyDv5SQ7oy22Zy
8OIKmpoSMe3fgbYDYZEcpKNbKLslPfKPMi0IFtWR3xVyAGOQtZNSh8f5qic3
GhrFaolWzOjvJ80J3OwIx6vtJxfclYBvmF6ZGpDFXa1Mhvzdte/XyGePjrL3
xCtprr7hf7MkNq3Vffd/lCRGlncxOnDVREbzVg/r4x2IfD/7oF7RNd4tfHP0
kNU9rGfeaL34H/zbyCK0ng5JJUtDuNsnWWKEI/ASjdIGqkzuw7ER4tW294vX
sDorA+e+BralEWKMStZ6kgYuw0fBdF5K4oZDC0V7BvyU6IiVxGoq9iMWNV2K
d+UnWSk+FqGrIdeZAa8WNI9KNuhYKAT4K4gUEajI3UVOAcv2Kzb0SA4+5tAN
eDllDb96FQx1xdkjLgPcmcZZK/ytTc3myyTT8s7H24DPi2CGEDB7B04FKFhu
MtpNgQBqSgSnHxAAuLSfhO8Ntro8CVQ6JPhIDefSu81ZMht8/3RSJBNBLMGX
ikwRmeaq9hUQOQAOH1FJMx22aY1SXUw099MfUmq6kzW2M1gJkdN63cUEn1kb
sBEkFCWpY7dlVnSrREHefJw/2FT6ZyEXw/7ZmMnY3CYnsYflAfAXzOkEyTrO
A2bYIu3vgC2oz7hn2NokQRXwVYqZ87n10Y8SWwvdwrzGLjvIY8oooDLLk8TO
OWTi077tiudLJMoQLnOHCFdzSpQqcyWrHGueSF0UlBbgHtYWhUMTea9L8EP2
Uh5Z0Z1d6/da3NnY+0r1WD9IbBHo8RpHRGaUFCIEoxSFJ7pqSnURWtfUrv1g
sLaknCh8cSfajAqlb2qrMXDr5plDlFB9/JebF0P53zbyNF0I0L/YTYTwCEkJ
DZEHN+BvZi3YEh/iDRMVWeVlWAwz0PTJDNBxNltYw+1YINZ/2LocmHWzCBlS
KlAdwQECqYeO6em/d1OCTMl0R6j46o5n4uEvcUGgFwL0JvPWIgoogD2V7gJc
vjMSC6axV3BTVFl5aAffKsOdFU7BslQURIZEf9MfMQp2J6SphvmlU1jIyAIQ
Tl1SLhJE5qDV0NW9FuH00nStk/hJCQpDUOCJ/Gef9utyx3xtTKHPQcE7R6wN
x1BEhk6qj1EXR39ZTGXidN1OJFu0X2K18cpbOBNpnjnslpYlTWrwtfD4CaUA
YZwD37/Q9nmvWpN/qKooxZMDSjJMcke5LbybRTIwYj0XeHbEeXtgmGIPj1KD
oufAjDYUq29vSZ5myB5ZXA/mfeOnv/NbYgQIMJwFJ9Vlqtwgl0wiY9AAQqtD
U57VHWZDlIz358K+dDk2q+H/gPE0H/PRD4r4I9q1lxQbO0GXRv0eWmVFzBa/
PbDAQ97k4L22nstIShTSwpeZvj7F6AmX7fHnn4kWUVEhGgS5MOh7BnIyWr7x
XMf0rswubYdt/080nBUXbjZTpk0KgzyMJdBbWJ5tOQWkwct0PXyiST5m7Uwo
9rnPwJOGmwuF6JUi06J2+kB7bUtgrryipujmhWj4vNzcKbSOdvjSsSTDnsjj
WgH7Mk6wQU/7COpJTYCc4/qrjn9AsrKblVtULInDrqNVyQ1ixgfxX+cYsq5a
IpobmudtvaKw/p5kdO8THIGfOVua6UNIqjPZU9kkWZy/3FrjRuY606fT7a2n
ik9UEUJci/FxVvUeHv/oLq7u638yeneWwTnSLAibP8nUtn1djczoqlmz8nMZ
qXyB7BSJVQu08cASdLF6tD9Iee+/pKPt+DlhL5NxZ/x64Af1awvoYrx5jyB8
564lqf3t2t/RJBnofsSa4Fpdv+d6EnPDgNjSHP45RQ6TQY8UtRmoABVaDnNJ
yqQfK0ZzuoFvRhcH1hi11HZR2U5xELZEq9Qoe8e5ri2L6jHqyAwEMQJqx+US
kIRAo1/d8r4vYPjKYgbudqTC6FliUwGYDGC3G3FSF4ti1yNYKHW15VKHGaKo
u/rZzXxTrVP/y4jzCznzPoXR0poMJHuVilMxj9EcBcoELFr0jntiZsBwNR1u
G/Yp3+HP5bB3zeKl0Gcagtf0cwn4ByCYxEdm31s5lK0tDJTArSCP6IVKEh3J
2B77X8AdyzfPv3LUMT83XXxEo0GotGY3pv9a1ttJb6IeyZheF04HSrAj7d14
xmhmjYDSCD7x2KLnyr71e6KW+lV0NXqINdXtG0xpPe7SwBPYuJed99dg7ePT
hiBXdk69rgB2nnUwD/2BoUvDn1l8qWSVA4uVDpxSamCKBHzy19oKgxpPKNdN
Kav2qguehfq6h9tzMxXTO2tOsKOn0sxvf7ZzeP0+PuA1XQ6eZKUp750uILGo
iT9D9cPwGp299IQbCjmu6e0oh0+hlf4B/WmuQJt6hUGt6bAg/KImWPr01p1Z
REId/JwB5VNrYMvkMvMfnVV4IGMOh8h0S2/CSODpNqDVrH7tHjDYFgvDqMBf
4KF6SyFIwJT3Igjd0N3utr9KS+7aaxjlZ6wRLA0b0v4WqpVV1XBtmBxyuEa2
yzxqEX/E2Gnm2u2oCuOBB7d4GKxB2Xis3HLWDbHR3BhQASLA/abVoUKuxc8+
iFNi/17zq2RwqSjeRrNYKDcpIolSusNFcliwZhgVZnPykjfuzmgT/0S9bNmx
mm+2Z02BYVxS5GYTpgXfJiZQ3XRqHlZplf5OId6aFQ21dIqK82gRevRdw/ha
CzYf0xcFyAhrs3yVCKRZOiKO5kf/ay02uJpTcgF4qHu2tsKDW0p4vexhStrm
S2pMlFrjO57vT7TxZdqKBy3/jLX9oyNjw8ITTYW7QU00DcoxbwY1E844avdQ
NHN+Ffij3wS/pyEtNk5IsHbPWJy4/y+CbyPqGWxkxHrROffI20cxuvkPOIE2
upMKuo+ZxN23yOD2F/jQYsStVujPxl4l+xIwSMGykFDpWOkmmKlAdqRijbui
MhiY1l9ZkiJl3iIBFaLZ+FHlIRQk1Kr40vxdvT3WzUy4nOa6tO1mZk33h4L5
+BzfInS9/03XpY3ERMB3/Br1NX1Hyn0NST0qFK1OyECBVe7ABxgAzFwmjFIr
n3E+Lm6XEgnUwTnMbPyYnFBtLj4Bfig55e5PVsGr7yrHG52ydR9xSrMrvmQY
erFFGNWNEJTkHxW+8EEGaw4qR2dj+j2DwVmW3B/hYjAmDXh5nRjsSb8HtSWh
nUxHm4+ou0LmT4J54JlVLHnQPT1+oiqTTWjshVedRsZLiRXfGZjYSG3suxTC
qlJ9amufeiX4fxDfJVWeLLHjpfp0UMDQzEFj09mOdLdZiKBbgHLmrsXz0NLM
gHBRNz4kwjTTHV0JU7QO9/8XUOMd0PBvPz4MQmKxrglXVgHYWBCFEge/3Fz5
/mRtQmm7r33mfn9iFSGy6Vc7FDqTgmAqxxbaAH4lMWBi6/dFzWq1dllfSSc8
ht+LnRubdFCOmKTi7kTaTU0iOd9jw0/tWtxdKASTOaVuJOY70shKvWmsLAOE
Z5u3iYHJTAvn/z/o5cLJl1NTQsNAgtiVy5/+RmGXPFI33IIY/MLftqD+7ZU6
osaAk4LdR81aGexYzPWIFrkXFk0oNn/Xn47ArlyuYn8UrmiyXCPWniBqr3z8
/wSr0aoMfp0FyEOpWDUDylwuOHzpPrZGOxXaQEBJfnsbeD6G/GV1FEGfx7f5
k5tZGVIG5faWA8da98zyeKYcCvuUOsrbEWN9WQritptEI7mPNS6TfLxeq+LG
pHn+xtopfNk/3RdAz4e0gZUB0z7ulvIKgnTz8Krxl7ASQ4AX7jKk8ienV5g1
/6nIsWA3ubwQoqrCxVkHKd2RjgPKclsxroHaplYb1RHsSoEe2vQjpHPeR4gS
2WvafYxazxRSz6S37sjHyWR/YQG4VMANWt6kvFK/KfraL2+8/31g8tcbYuMD
Gs1UaWkRHxbWq/qKkl3QA/KN1bX0yJqJZE3iF+KzdVPiv6tIHckOj3KKmbV8
sirloA9ZoUeZ//5M0sDwwnuh3OMyC1w/7fZ3UXrXnDBY+RRQuM2vxWwbqbgI
EOvlcRtmB4scUSL/gXLR9ID410yRfXYfRyyr5KbW6URliUClGGV150WDd/6d
pxTJqMbK91UUFYzi5Zb+1fETrSLqQTNIaPyN4LVvQDyzhkR9/MmjFc5wpQnR
1SC8ArHD8+4L/p7+AbMUHwh+X4F2Qrwc0blC0YFo+XGCluqDlyYHwc+4jqLd
kio556YySqwmpac8S9XtLdyUBaclGbONHECc97dpi0FdByGbEJLlmn+ypn0R
jc3pba2iTM5k9JUL1wsZmZL4OWRLzSuywnS05vXhL5dDk9wTE9K9nD89E6Uz
D9t/gaKUglFQbQiW6sIKEJFV0d3uXKNcSK9WIBu+06L7FFTVnKqZPimFfHkA
FHgy2H2h3qjfVBWy6O36DS4tAojwXImt6R09qoRAk2xU7kiRxJVPK/vs3WW2
WxhwSrYNrwN2j9h4B80qciVGHNyv+WHUtI20fD+sP1O2Flz1Rzhgw6d6981Q
qCWostLU1OKQc5RzfHigpDMD+lp/Vp/+VUYhER/b2xHdV7nRYcMhw1ghiLyW
wpFhpcRG9rKPpTk0juaxYz8x1PRNM9F9wjLUJO4AMB+GgQix/FgPypP5isZV
iuh8EOELXvfDxxddOklmmXRYwJGsCAabWFjlUXU+3W/DPoXM8QdPPb8apy/B
0Y6dVxML43ENmOegm5jMACayYNEn74jqefjwN9pOWR+0enJn1hmSna9UdC+e
LBMNrJ+M86VwX5PPXgj593bwHaMvvasJudL4ofNv03l9G+TMdzLUABnNnqAS
abafRRU8VIsFm/Y6fS019+0eP3k+haeY5hCo3Zvtw4xkbdamb141o0nTd5/y
RJJXl60+aUr3ospTp0JxclQ2FNSCKkV5sDcnw5s6a0bFajFkySHiC9uv61UL
0/GPICiXDJ2G0ENhvYTMQpa+8tsubDXPLOH0sgRLdk+NWvjt0moynzYAtBin
xJVQRdFbmsPwul3OPaUPK4BliXBLmB9IAEISbvAMqbeN9Q4Z/dI5fsK6gU//
zlDSrIyNMfqvmPsi/XjE5kVlcf8U+dyRJ/ebgThNf+8pVu3qqUcN+/JdBbMW
0csPEgZZD9mUxW95SnazaBkUQLjvnCfN/3SwtD33BJP4akmeQnZgy+V5YT5y
WToZLkN1ZnZ9Uasvrz7JXodBpPXbFq4IpZQ9jbq47bUeztiO7aqlAzOrTqqo
sLU7bLJTFT3lHs27jv4VXOr1PyJD74HPN2S9TdmMXGLQcb5QiGGTKYXu/KCF
cdb1PCuAq9E3xLQHDCLS7jxx7Nkq9aP9zXHuFqjbq9//cZBf8hndv+foa9Xz
Y0AzbVz3CS7l9emezsEzhu+r6PIjVg0AYxkqmcSRTlgPVOKH+K6ecMZ6rHFT
BkZj3guzRXNnirlgi7BdAVagSkiTmr5K1w3CmePmiABu35+YuOItoOlJPL79
9wiIW4fonzN3qzeYFD0hNJKx2A32CclaVUyete2PQEcKQkFQjbqa8T3tst+0
1ii0u2hX1cyBpO79o7+kWC53b4BePXyMaWQK3WjgSDYNxWjg1qv7/jKjAMEi
rB4RRyYBgv1hhYkciDly7740pwIO7O3aMaMw0NfkNvGOO1bKKa0kaK37wNI4
H8jRt7cC6xvegmc9Kr7J9v+Hc5Z/x+Mfp/YnbNJCK0I2GfKoztUJVIsuFwPz
oTJgAqgv3y99eLsEcwDqlkTY4mXZOGUe51llrWkxZRXRL9JFUjqhFl5ywgGh
gCKnSY2FZI9AcL+P3FS3ivm5TiqTF+v6scKnPcStG33J+nH86cVFR/vp6Jj/
C+ijyA1IkPd8APDpCeBJQdSnMr6JGmF7h9Y4XipjoQcVraUjmk/EwR+ob8pZ
g2CWiegra1j2s+S8XesHuFybZtWy4Shf/Nc78ru2r58jWPKcTDJfPlENnsHu
5T20PzSkX03j9Q4EitNqrXNfO61LXvCz4KXHupqv+W0uhBSl7cgkFimaSgDO
Owm16n6aBfdKErAvvAr8ET0nq2+K3PoQQn+pTvFcQSIxQrYukLRD2sfdet6P
1fgCkohFYx/TDljjmTs/XKLiaoS/001McQZShROQcCQl2bdmlvDVQuzrOCPr
rRaXBJRDrCG7kigab1aQ1XSlQpkG1XOGGZArTfK57LVkDdMKvsYrqO5Vj1l0
TbQrRL3VyLd9p2h/xe29IBPTJHWEm99cI317M8Y9sSGF+LLx+dUsZ90AyoO9
zxlHXUC31bZ7GUUZTLrztl1j+OOWxkcEF3oDUbncQG6Y5fq3ddfbB+VoYXjL
vBUff7BoJIl40pDE/mFb6z9qJ2DSjhAkQbh5QwsKqMH5EyuzV4zLjxlMSTC8
gUc+taegcCn47cnmEMwsEwRsZ/lp/+NYv2CR1l/6jcQ8Sz6mzAvysKWNYUg1
SRb4PA7JijTmxU9QHLuCJKpFVSYYQMnci0Cc9kOQjWnEdjECaZM51vKf09by
OiXLFIQ5V6AR3v3YU+5uXtGCYT4OfA6qsN461eS09dffrt4HSiXObMM9okdQ
amKJzwykOmAbL34c5S86renX4/uVUcO8ejyM9kiT4AWma6TttVcVq05H/hbF
PFZGqs9pi4aB0GVdfmqvRlgB7z/fzTR17G1GJ+krPg8IDkyPMS3agML/J4O1
Ck9uagy0gtrjwKOiz+u86yIFlVeimlchQsc0HjDlYg9LixWbDpuSdW2J1pT7
rCZjhMSi8xMZEz4bMb4EuL/0XSdeoqoynLw70Pggr+raTli0/Ffs2unK2kw4
C1IoThL9bzpgwo+Tu84TajE8QJq/d3+OhJeN6DCj86NMz61hDagYpXtTPTM9
pBDSKNDsRAD0JplqmqVZ0nQeDZ/8DIj59eJ9Q/fIQZtNbhGDK4x9CwTDlBa4
Z8fchbl1nI91sIJ95MYPTvW+pMwaAVBewR1JjDrJcOFpqQWqwTRqgRpmp9d2
DNkUqQhdJH+QTFwGL6MEMfIsB/jVFso5JHemqbGfreOpaScgYFTJLJL4aPlw
kD0eYd8Zrg0+aj/KOFKpnlnLC8PTqlX7hRWFg/AXu0fKiFIFCTXlTz347pfo
otOifJ6ChyofM4Sd6X3XDryHYIuEeMaz9ZyV0r5LiNcz5gW7gvj815uBLKoS
FNDR3yM19+L3jElnpCkqxksNbKZlwKkYj0P9kVZ8BPqBJc6w7mSIa65HnQyc
YE9rD7AdQd1sSQ+BJcMnwbX9+lreyOhax/UU6OQvPPdTECCjHNY/bk0b5Hn4
ISMtgwXQS5+L72+JgIRl6zFNocCghvF8E4Hp8/qGXXvxxJuvo8i1WiMFEW3N
23QQLKe6JMehmU9IWhwF/eLgZdeezYSjByW2FWKEis76GH5nToMkuenWGPrZ
sfTlJ/nJat6JvZgcU4gxSq0GhI91xiALTVAbmzjzKta4RJijX4vnRYE1yone
Y/XIstoWusysItkHorNwmXxeMpCEAixp+KFtD/KrtQ7jIjoh7xYghXFYNUH5
2mFFfB49d3Xome6lS6PN+8G2e0x1fnBeRY5DaMtMW0bJGln0Am348R9mzIFF
9XJpoJUWk/Unij45iIodpHYR0rtEjUoh4j2qlo4oVZjq8IWb/5tp3743N3Hq
nQHPzqzfuUoH7OIp/jfX313l9IT3NrPyIPulkf/LZHxW6UyaL66Rk/9EssbG
BJpmNQW0sjn1h7AsWHSCngfK9K4v03ju8Tsm7IwhBG8GnRqZK6erTHlgge5y
zUBC0rUWgY2313ZZOIfKIluJgc6cRGb+LMslmWmZ1Ml8Tjj1dIOwxrCYBIGK
LeMB0+k4ZJsZv5seid8PlClYmxk67LAg0WZeu0spevfVS42mOG0pCfXTCRUB
IeuC55tMJUUiJ5Qvt0wJT8roKSW5MGYqy78tBHgmjbU1YoDBzU9Frc8DaPoO
vx0Lft4guvkcY0UBd/Y01idZIj5l9IhpBX7qJToYKmnJ+bfcjdwvb2Tc/aB5
W44MrV5mDOwkNIZOaIXQqiLIzPCVxOtQmLzCBfapXA606fy6wluPuYHNR+rk
hy7WxMJpDITZ2mRfgjfk+efFcPGQOcOoQq5zvAd1WqQxWmEaBnCTP5dl2O2p
3I69CPjQa6CYwIvo9n0UkF7l07URNg/mm/4XtCuGULXGRIrZ3CcdKyJyZbAP
iZtuESY3WJZ6FcRJEsW+cSxhT0EWrzckgdPlz3eC1rrkuVT4ImyHOLeAN+tQ
L8BJnWOPChnl7zNYgpJieY0sQPJgID6CNh+j+dujmcjRQ8sm0LfeIHNQWtQ4
2S4zrClbCPXCJM82b95h9QCdbiRGg0V2JVnzIch+Y3+aYqhFfu55Iqt6EC7M
8o08xM2hxO1TlQkfmHi/SJIgRYXqVIgdMSEYOZph/lQYkR0qI/rrtR/ltpir
4yzQeLlrBhWF5XmyPduQeGT1E3+iGIocPjdoG4IIWRh/hM/hnfG2Vd+8annQ
DFiELXnHbk/oEC2kfW7UvNXZJI5rb0a6XYDKDLkH97tRVFjXUtBIgquZSL31
9St+oSRHOc5aa5UwQQsMOhwfs3MBG7xOyoGFpdYQu6q9pvD3hK9J4vGXlKVg
5AFhEABwrJa+ksEy9zC8a0zspV499uBUiGgtUQ+691q4/3CABjCwLFxoq1AU
yX34asEaVF9sfCo6LhcyPWJYFRKGQNOzYs5Dkl/Ud4BdArPZwstDnAntvvPn
NtX3jFdFMCbukcM3ND2EqeHmJ+M5LSVwuze8UwAjCsoSjgyXyt22mjvfEHRu
kSFE8b57oAKUimA4F0JUbMCUw89b4kCtW1f/vvDdTvIJj3ZB02QS7/cbz8j4
8+2kgDgMntKOEvb+pWSUXYEg0DKXnAVol+Rcq/DULmvrFHpWpzgasiSpZolY
xH+iRlETDoXGxEtW+AmBZr/VBHz3c9C9jYsenlGCV7Tm+Y5YGT70iGw7oPBV
5JvIEKbsMeJjzJ4igaaloPLEMCYavMwhXItYlA9Df+QhnJl7f/abL8pHCTjx
YA+FuK4Vhe1JjZHIZqFyQfFdwjb4x2dBmMoePR8524le/+NbUYI0TufIuqrD
DdenD+1WmOTzTMROOSbL6AaLWhSBMRzVtEs209EE1pp825kp0Lb5x/Cw3cQZ
Y/kmvpR/fRfGvBVGiB82vEWTapBiwJCmMZ6GBA/ZYqMOGYjutVTHHhw7eV0z
JxpzicpobH9/bo+XGsaoLqnCfRa0P+NMEXY21m7g78JG3V5+FXzMy2uAwmIF
MiwdM8Qoa4gDADbpWqqAy2PS+DOs3Pn6iPEk/zZuNIKVwB5/GP4fujiB/V0+
i++22g/9PjfiKXfo9djtGBLdDX0dZNAraJGAcxoHj0815mk+2QywO9vG/+5n
QlSOrLBv+bki74Pnv2kh6qREswNvWkQQEWVFZ0FU4mvbB8PYLJWlHU8331Ov
0reRxnq0a2oFLlyD6FUYOfCjXbA5o6Jc8wjzFTWf0/1Cxl5askZSkPUxLiVQ
dzDxqjfjNcoNKF7VslSVh6N6jcOl51+LUdwthLgMmBAvCNqGTN7FQaBbyQLk
w9yeWFlp+xjyz7lGFReYiCYeKXIJIoES2rDsJUGgMzXa1aqfs55g7aoM0rgj
Aez0ECo1LedTekLdLQWu9qJ77ebGBszfZUbuGKKGJJI5K1U9jELuDpciGjA5
bn4/XKxjBtc9sW58e2yF8uCCjrXRpb2dmkzgSOOrioAtpY3I8+CjVF4SteK6
FRPTF+XvYoG0YfcJ7tn1GoyOyMYCI8BiDnJ74W227A6OQP7OM5Qp5Q4chx6F
bhYmzvaNrhcjV5uoRM3QGQz9TQYqQRf5GkIk7WPeg7rZCxvupDfiAPA0UfXA
nr9AGUjUurGoiBLfJzWUgjXAHAovX6zf1T9swM0IZgX9RCrEMmxk3+XyjFdQ
GOGnkiEAp9UAyu+R7Tcz2RjWMYZZrTznLBndjB47v+AJpC/yv96ENab4rLI8
P27HG3RJpoKDCR+mKBk4FVWZM5XapmoG9fCUxGIWy0suH7P8M677LvEiUY8X
ue0+n3Yz+sZ7LV9+lZndcgZiyfv/UNwBzz1r27fRZsruzVX0LKrUxFiwtSeq
hmRKdRucGy/56iqsi1+7pFSEEAzoU9yRqWoV0Uk3Oe9Q6bPU//4DUxdz+1QI
vZnGmIxTzcfZU+n5IS3UQMsmZaK/VQWXNRJ4KGhBVsbIb0mmaY3VXcHWF3cC
YquFVGR7+OhKF9WKTHT3uwse413Nq5zA9UHOTct0DWl9adxf+JYoljZWIHK/
kjArj63YL4F+Hv1fOIiTJJ/T1IkJm0eNNt6dFFl6mqpy8UBwXo78B1F+PNeS
IrIduBWOY3Zl+tHD8BLJad+iVIyH2KinEhQ8jf+O5X1v+24mr7K1zeHilMmp
dYpap8oJ/WMqaMWX7qG3YwTrti1ws/XWb9IYUeV0vj6QyzyHj3AgzItWJfeG
K0ckQ7s/27Y/3Rua7JJKzGcHQc6ky34fauZgyov29m+vfYlqzoWJgu33psdl
fKNwNc270WwNCFN9Fx1nPMWw+E+LCuQrLXtcLnU6F/5EHLsCoGvK25n/QYfi
a3JeSISz9RDzIKLU/l3aOST07p46Q11oeMAvrKityYpFnWX4Zx/C8G25Fj6o
e+qQDjul9dAXNLi4U/fzlyQCFnJKlpTvut4DYzl2Ll3POqrfGxXCJrAw6VGS
7I0hwBpw67HxOpjphPiRBfWg2NedFPHtSpkExjB31g/J/DCZIdvkaoBdnLZf
r3dD6H3v6vuvJYK4zQe2bhvZUAAEW3WoTEZ4R2KrkYxtT1G//B+aPpN0F5lD
LelRWXQwy/z8jRlZqtFTql8Hr7VtuCTjjD/CaTgq+OL6aNQPhIx/t4FXZB+A
d8O/InAxDx8lW1FcWj2RivjjbXRATXzwhjXJomY6xbpLKCciqWaXuen5OUGT
Pl2DyS/eM/NltH/JWyYYpeAeYL7felDEWyDDEAKGpNWxf/ImBaXO41vQ31qz
te2aAxFpwqwd5nK4hnG3892ZZfxk9Qu3eHfLlcbepZbOHK9udbGUCzcgnVrd
d6Pq0i81a57JHfVqfaoB8+7Dw8VZy+Ceh+bDwbzSDRccCmjVzmFWpQz4jyKI
BLWqg5+AqWyZHLvP47M1ovbl8zdr5Rc/a6wnj7prDOZwlvui5T5HB2tldGAG
4iYMAGqV96dkAe/5Tyn+5hmv8A5qBk0G6LyMdBokA9dt8RLf1KWljSx4WddN
ReZvGPQx+kEPwZA+siYG/8XY14VNhmtr9r/W8GfvIUOi7VDbBghxPbEcSkEa
yTPLu0oKMtQzw3uBCZ5xlbpeArUQyrp3DZK6YJktzG1H8O+6nip/cvYsSzIV
LSUjpN3T6Z1jX2q8nfX0vcZ03E//CEQnw2b7RtRG6+KCD8w00HvhGQT0PO/D
tHU6L8zXv9hC4x2/VKiTAD3/8xlsDxG5zt7Qeg6C0EAOSt1bV5bDxnC8zZDL
m/yK/pTZ88AsMip7/p9StCYDVv8jf8geeqZzrrAqDa0UrEe0Q6y2KqvqWjAP
+sqVtl97HwP6jTUgxCuyv0yOd00pC5T8KLtLZgNBp0etEzk2yGKZuFytf8K8
qgZGZjJNraMR+Jz0qwIBTjodNpj0/WQjKg/XQZscgcX2IdHHo0MURhhtbuf7
zAnRMzz56pt9LFv6DwhNAyTs/I0l6AWsxvMoqQR+rTR52lmVyOhdkyqD5pOr
vx9gHRfFXW6H4Bd2CI8/qUoj2ljejeNj06cblSpmyJTfvMv3xH7LLKW5bzE3
0d6Z/Z6kEE50ks4k0izYslFuLVguxmlfzAdWRTUXKuOwuAOlhtwlwDzyg72D
NXCkT66KZPh1aE5egl+rZteHX+ifojvdw4lUliAeTsh3CmFIC8DECsPjUIkg
G/IZU4XMsaP0ukfoZxynrmfW5oogCBxr9mIs4KG3Tq5akWxLBb6SJngBAQXy
7az2fJIZqZxGMXxYO8x/svGxb9nTmjyxUV0XK+oxcs1euEyPYSrNYQ6lt9UU
7aPT5VIJ8wUvBJGRLYHmWbGdBcmq6g6I2I/gwA1e6nAPOXxyBUrXEbRscoii
I+4MyslMWWVYu114ydufLmt6RJ0qr6zzcbsQBZKrwoz1KDg4toN1npV8zEDi
GUOLnbnCOfB1H6HV173x90V5OQtFoFxNIyk0457KtqZ4X8f3jqvLVzl1lqQ+
Ed2nG7iAXjLqp4SLDsYj46BtFCS5DbcVHnY4lVAxETyMxd7hPPtRPLAC38T5
P6ijRPfXYkFSYVRp5Pjg6oNCgRJz02d27umBcc8nHDmK8XtRiTvAOMvlq8gc
Z5eLk+mpve9/mSG9b6jUWkUhyPZZto/6oyn4KSd6yVLirPEqOjNJbQ/k0i4K
nBFLSXgwqTlZMlx+JDRlF3b9b+zOemEDdmJ4sNXcojcGk3Z2omgq5P/P3PJR
YroKnmggjwTAsW+PA0fTcsJFcyok/JJjdnP9YTEB4LmJ0Aapjgaq6Ejao/q/
9XKDeWHUYz2KhSlqKD/L/OpRVr4sAC6OXsTyV9C9tsFiXgNaww/ffTncTQwS
Gov+Mq0lEcq+Icwy64MWEJXjHqZedhhOeN1sQobNzEG9VPM2ScPaPbMWTGC7
viX1deCkWk8YFGDlksZy+zq74OcYOeHOf7OGxSeBnq+6IR6y78weIuC0DaM0
hKz3dpe8pD44pcLavJTEiOeRJFcre3aRfyeJfkfsQhkLjnpzGuZ7aV678G/5
uNjqiSqo+/UNTI3dq43JyzxRX+64YfjpgfSXo6TPavzmE8woTmPoauQThJxS
HlZix2+75sQlokKbKNHvEbrlMzR1AS2chkM/lu1l91azbmQ8sCtCYo8ItuZT
3mXhno9Er8/wpRbvfjoHMKZdUhLxgL1PDB7uN7/XofyMUGHcjMwFVgHUpxM5
4uLQLBoCtWp+ST/hon+gep8nB6c99jiptW/l3UBC8WcEOEb1oSKdRTv8xL9t
oYjk6KGtfY0DNwwbQ/LAV7pm9JwP4W1nEfQgK0ioWnpPctU6HJ5lBqxKUQ8V
VX+GdyMN8lePLw+9McRPiEaSD2ZH1tjRLZxZy+V07VR5It587NxtdIhb6LKH
p7qsNe5jSpEM4XhAsO1Uvrvr1Y37R/zB6Jf92/79nQwAc02aT7dQmFfW/JvZ
byQ7gzwzRZtP4mYTXeWqX/p17Fg3D1nck302OOJlrZW+QGZvULIyd8h3ywr+
AlZL7VT7PcbZEm6pAT7PLcN+S2Ti99qA6OqsbxEhMli1pZD+mVY5N4MWuPYA
RbQtJiuGLjVWucbYDCrmlft8jU0BlsbrKwsZavzpLgIq8cLWe/LCHn2wfrgs
JpgiQrcH8DnM7VKWleJBq4Cic1n87JhyCT1MNvaf+n8ARVR0FG5Q9SzAf5z6
IZ4EyNJ5Kh+2YyFRgzikggKrquj+8yhqQ8As6pbJT+sQtSZ5JJyYlhAniOiw
0/xR6FvKCXFlKDkEUdrdAWdbNiWi2m82ahFxHIYZtxAdw0Lg/V+4CiDHZM3C
SVrpeTVg9fxGVyFSPpoUuuJW0bwbo0Y+M6fZh95kHVY8w8Qgdl56YfPdFDV0
EHBEhnz+W9DuTc3fEOcpECRRLlfRj3nwvuGOrkypcjpTqhCRH18+2jI9+A2V
4Gxiqqa17jMc5AF8K2jmNmnZ/oloq7bXnLhmtoiz5BotmuZSQKpU/Awl64YQ
hOw9h8fkN7Vu3nwl9rPC1FZfEedppMft77cNCz2mxQHgB32qOvraJzBSO6My
Z4igZ6Bv3uEjZtQ/qj4W+vMMRFvJqgbDW7lzBi8rFS2IwllTN7OCXVLMwjdk
8TmX3moTNBlftgaO3+U0xCw+BAcJ0D97S2ix8lK8aWqQ6KPoUw1CRYZ7lSK0
m/Q21My6TVRWcyjRdV7n9DKEtLpTsQxyxlkhV9rFENESzEqEdpDwIuWb6V/w
3jYCRlm0UsJY3ddlzNis4oHv28mH3reE96x2rUOeGgdhm3qAYKwR1zXIDiTD
6cHcwAHTAsywWE9JyQeuRuHusZoWC4w/BTHGZWjgrxZWB2Jyzw8hGYdQBaey
EBYQV5yrPAmkE6t+yRYyyqcXXOSfLKxoyydwkHTWAz+Eg6hYY4mlO6Jx1t5g
LoILao/D4ZSMHkF8wtfvhaovIUnG5wIj5v2t1ZG0f/PVPQ7iIK9WoLggfAX8
QA585m5db/XcL3tSFXl5jCqPFuj+qR4ydZWdMPWn1er2FCBJtrrxzxGEwcb1
akT5+ib861vtBLh3+BMVCSDSfIl7q01Wd94Slh8VP5nWhHc3cDJlfOnmPQ3B
ebnHHhgLZZvrYDiYA+2Nfp+aOF/5Umt0p+Y0WXrPVNbDiSJKQm0Ug0FwaWqD
NmLIoXtCxwF76Yte8MiMCn2V3JqX5UP8wTgWOOL5tlVDAHRtkC6P+GVYULnc
PhcCm+BvAZeMxJhRkepno7uDXnYjzLD2yvHKIEw0Ru5JqyR3kPqPW3vOYfWV
JtQtWGRzR0fOMgyGLhP2/p2ByjXisFWPFR0CpAf+Z1ZMrmiE4rlppzOo9pPf
YeWpJJGEDbx7+fRvmVxs3NFVYOsOXBGwaawMowY38hMnS4PPLlO1noG8Y51g
yIoBA8UBfkB2u1IRa8zfPMsnZhkHmRtxy/xAApjJG33aHSmDCPdrwetjIWfi
zgqOTDE+7OE6qrEL4HfDeipwG5DdNFxBmK84aLfuSzi+Jc+dT1HpU+qotf2E
hZMnkJQmhNEbS5msS/Z5LZijzY+OcPaaQUiFBseqpgO9/Cg8WTmeVu7v7AA0
mW7N13xtw8cDSneXlGzJoSUqlg7RluNFsm5o/f0Px6LHeUrfUufsyCBbDlqA
rdXTZdg2GLdulDPHpk0k+60MNR6QkQtYFItx/96oEJ/BgW4uBj6sleEb5mz0
k9zlMKtZRzAeFdAQrTVClLmbK+FAL/lSCzlntk24U5JtDY+z5HcyEkjh2ukv
sdUdnWGnPJhLo3w5tNjcgfsWXXBAbhSvyAg99+P0uiV12GXCfzcLwBlj5CY3
C4yPiixa3uehyXZXzzJEVisa4T0eSqyqN2GmcZsiTIsu3GXzay3d4R7lkb5k
O4G5+Ef/JLMHfzPyySUHi6ISFY9lafkpcrYONPxR27/V5oSH1e82qkxvxlft
0f33ChlUgtkYdQbg6HhSFoxjCBHxVXMVwZfQfQx9HnBaQiV3olR71PI4Tu5d
Jx8XZsBLxGmudQGcCunXE60E4XTH+oJcesfmGNMNrP1eRBJIIsnKaR0McOZp
g/+TgnkOuTuKvdIGVNf7sDNircb5Ks52ifep//3gocc6C645NgRY5+mmf1c0
MLeG3SYbmbXB5VnDH+4H69PreWd+uSKEki2GwjAEFlS4w3RME+fdeYgR9HkH
mHwp4JcqSKNUAE+hjuC7uS8aBf0f+vZYvd6vjDzDtosmheJ8ffBoI8z8ypg6
bJe4iSxUatFkHYhOtNzWBJRl7UsLaWiYA6VDWw/Jiih6jxBuEaTkBnZlWS6N
EScjT99gFA0yOXp4neQUfQ5n5toLzotiYbXLIyhDPyxy0tmeCQJkNRukTzd4
R1d6osfN6n1y0zfra+IHLVFy2e/O4nYtvElXYfM6K6pnxmJ3j1F7bezDkqbp
JQfQsJ+EzmDSbYttsym+6Lf4AHoFN5RGhSNjp1Xss5kNX7gC74nKyGOi2UqM
pdA48BYWLMg+Exa7rl+5GLLd2TBObjxiUDoEv2nhGdatLwb73u/nwHWB0PMN
SlXr2yQ2B96cAiICNJO5JvFU6GIxa8JucdIr85V/IGZA+7vIdF+Ten87Hiov
6g4i1tCMtPNO9J3gnA8kc7VHmnd+dKZUG6VZCZg2y3FKbK1iw+jgz2GacEHm
gaof9la9H5WoMTTBLj1mjVeWw3i+1g3PbRFPZW8w1kE7HFkAuF5aGNDlkQ7k
pzpKDxIt0F2BQNfAkfe2tNdM/OAbzb1O+70fcm9wldaVj9KrTtkndfeMDp9h
Gm1u/lcjBspFQ5WfDQmK6t197CpTxUSIOWDqW+caRlxWvEWQJKHgNZamQ6lh
YNFkGrLuCDHGoMBh7N87hqPowIt6Slils2Za7E2pZp95FOjl9dKB1fCjwLSY
X7CyNVmPRbwwI/zI7q5fIJ2nyNW9Rz9VrsQZd9QtwALU8Rb/Jk6OcZPe4ZeB
HxsMFeZi4WIECJfzniGBhbS7QLj6umyDlUwYsNhm8CuMLoqNYg6Cb74SWaKU
z4Z7iSIwDQh6ygEW2uO54/owpLOH86M4hdD/6JZx+Oa6Wxs8oL38KM5c7rh4
NCbS6J5PAgdaCZ8gSF1BVkzgRE3v0qpjdu2aUU8mS1neRi9vqDYAWnYzURYI
bpnjntf5RBV62q1hjACDWoHIDN1mtk2+h1VLwevh90mP0/AnLLPZgjfgZmRe
cyvHKhVytrOlv82EtvJYUmYqyIdLKKd9pvjaGvVNaiKGlQNELvTomN9jLHRB
qJteXtv9Tg9FzaMq/JU6SfBZAvpthpqAiT72wVsmijOO5pRR3YLKDmaXdN1J
JXAyINk9V3eUINGZVr+hYVAWDbsDkVUrgAbnAlfk977BING9B4HkBINTSlap
fe07YAG0SEk8hjZ+WOacqN90p+qghyflvBUoc1VjXZR43Q/bgDOPAdVtKlIK
0IGKPOMfcMbhg++I+LbhaW/q2iO+IU+XezyjmgvITQBTkLaAhD77PdL72l7b
9U3kdrdYjK1ubLnJ2x4QQxHpRlvPjO0SuKYRyGXgIo9fD7rNAa8yghGNt6M3
pdzLEe3q9Cn7K7/t+4Fdxgh2d5ZJSrGOlsING4BlxqHz3ZGABXm3Xg+Uy5vI
YtNfU1YZ8Tt118QN8YAmphglmt+/rDlm54e5IR22dsrWmMav8m6XaJp9hxs5
mbdWReZWJQzb/xugBIv7lHBgEoROFjDkz6yPaYgZRdqnkwMTPKC3WlF8cUsR
n3CKLlMMI+vGq9USsLVOY1dRzz4x7bCWlJ+ctCzK1odWAADIsEseI6uG11qb
ziB5o00OL5ZUTxQcauFaQFfe2ES2bzdTigb5FTUOYxdnFDOIP2oqzaP3C61r
fFfIZmzocS2QC5goGoV5WF/PlvkKCRavyuI7qummle/d5pUijg2CQVEUaoRF
0al80UZl275BUdLYNYytWjLKM8gdlfi2WkbX1CcGpIUWghftIiMTa+4hSa/l
Oa/dkS0KLPzNE+pHY3cqm6/zNDh25ocqvpXmmLjRuRqMNotlbThVOvkW7NhY
8yeGE8Y2PfyAuNLaQUZN5gbiWlvbVbZE879ZvoXM/1wRBopSu/OmMLuDKZik
mtueUp+aosBJtgPVLCABQK/YdpLWlOr0q7mBsuk2XVRaDOS1vbWqpvcsJaYc
yYD2VomjTrVFeCVjB2ktgB4JaXtFxWUpdSNHei+8HtdVMRC5qHF8skKYSJBX
u5Uf1A8IR6gRoTnNSDmDaOf5DRsIQ5Z9D920ego/XWiNQtLcEa64+zcUn6NV
kOp6NvDhcn1HBT/RnYLZnpkgjyH9I0ac2pVT0IHTXTvT+WcfWdqZbczorgLS
jJnre3svldExwNMeMmlcSXjEvcWX/E0bNG4a7nXnkplbCAN6O1QopSzS5QOM
R9fNoaSpQ+snd6dGw+8FsDVmPJMA0msSnp80NEp/fkeg0YPI7jVpib7rzaiV
ULN4BNEAnr/6EfRgXuLTxdj32z67DKTdJje3PVB4Bqc53Omf1eWd8b8fG/mt
VxFvda0wSZv71tb2uaSe61NqaeqQsRlgz7bnmXkt3mONstNxbzf8jPeWwxPZ
KOTnVxzQg4vleUTGeV2Jo8dT4pkptnLF9pXh8Zu4BiujRGnkKTBEbGI0Nkf+
i90Ue3FE4uuCUtgBGgpPH5cVRgIbDdTZt0kBX/y+6hM2MpyptnX5A8LXUMHT
fz+L0HPfa2Fsk9t0q3zEwqI92Sxu20e4OESIzaQIJseF/+iCife9BfWjGHN5
6VMlcbjW/bJwamaIAcSOmiN8wlXt8CeKVp6vPawqiwkjRXJg5Nqb/FtSFDpc
mPfFkiDHtM8jaqRtjCacLftFA90blIOvHKLwSwEjfHFQMfhy+wPcucs1T3vJ
Z3bjZZHyu6kedd3bsNi3f1OpL9ZfKHcpgq2PaNkg7HMuXvikWat28kAjhuGm
bYBTXMWGzVQS4az0B+8T7CjiKc5VUG9W/HwHiT1vYH8xHmjMajNzdhcUmDsB
8e7+EoVkpzuVTIbutql1YCGqu9usa9LTyvlyYHuHZHIDMTqKoQRzb+yAYK0H
ulH47N6ANonDL3SnA8/WKLFQFm0gFkzrbamX7SGvEesiTEoA7eVqOohV/r45
4uX2H0A3zepj2BIxdWPdu7ZJCmUdZniOgrhW/ZYa3455XjvOzN7lPeFa/jgX
nTCdGYyyvptwTVpxUGpq7oFXbrexuqORahf5jUqQM6WGgda9GCbuO/DNqJlM
KFAEJt2EalyJnAOIGp9O00lrbr8tDUcCYemX6Wj4pJS/zWwi6w3Pku9mQ5eJ
SrTBTnb+0+N1wwefCUft8rdVpZNYL3nIxhPAgI7FPd7cnRmL9LaFBjAUrtww
cDXBqf+/RZU//GwuCbTn8rqt0SOLbXAq6jlYnmKktB0PLBC4lnifJPrwiGXJ
cYDUjQHKDm2xm0Zua7sibG0pfo9blp+qlDqr0IvKAOFB1OQtMTCQaKkDOh28
WnLwuAoklr2+7xw+czTT4OHNUDbO4DcX8d91B+3AKOxszydUaSVjo9RSU8T9
qhyM8JWO+KhGrjLuVSVdkmB0YNjv4KNvEbwxmWjIZMF1oQ6VfcmiFVz4TlFb
I2eG3b79cSr0t46CQNDXPh/nImhOgUfphv2v8PmjhkIt3UwXaeBzymwWZjGL
q3SJuyb/I8P8IHLligLlJrIF0WkfcCWUYfh4fkjVmXMfynE61nJDPUyUe2D5
6HwRRa+cgsYx9Rr1RZ4eaYUCQRJH45+LSShPHj/Zo3GidBub7mUfxrxSUKKX
9lG1PEp1So5mNlTSbfbEPU8wsDiJGb1vcoABvy+CVRMI0m5e/xmtkeC8lbnN
XoauRI4euI6Q/kE/Ixj3E+93By8fEYzP37Eq5TPgddnNSUNTb16+vnQL1tQe
LfTC0w5EgZo3JZb1mhaWM06NPL6l97Sk3Z0L4rrED95+YoiakZSImtYZhxMJ
eg/AneSZSoK2ZCi5brM+3RkdBz8/SJdKVi39ykyAQw/F/9ZATGz/6pDfoUy7
HuyDwU8Q8sQGUTZ0S1bvuoE3dHxyuvsxuh4733uC0bGaVK6SYXfvW2a3huTG
DIDTKhHbvwy7CD8AXG7kshtSRimZ5WuUdDRLeExgoecZua+vUIiaEP/BhJjY
eeR//NEPc5fh1RtY2jfXog/tsiBxVEbl1KHDbAV/IV8LC6EHW/YSO6rWWJEM
qKWAu/axHfKqc4AMH+LRpKcxuKA0obILXzm1L5Qn/ljk+75euok8/gVOJpGV
jdK2yW4vQ2pMHOG+cKm8tYXc9yR/qE2UMw/Jyy7WvvoZuBknrAAoqH2Mla1l
DnufjrVzalH14y3QTjwNwEruAZSUYLjY9dsU1tUPu+XwrGJDgkbIelAGX9t7
/QEZaBx3m3CV5ORcLorUgE4Dg7Je21V7fX80nLg6ZdjjdKErlBOOfn6lGpmn
0PhgJb+TKLmFjCJCh79KHp6yQhHh5JbRrscNxWIyDKQ7+huiGaXgzg6eMRyv
grLi+g8Xv72CaEShISaQtN0rsEc1SSI0IyRG7CxcFoOTBPsbq85rhalCYuoT
xkJiPCkRhuwlsz+ZywBHKwtvQ3+2LgPf4pgiNHU0U1BUH1Pf50kqFqKbthfv
zMsGkCDs50u1VVGyBMxoUJuj3LTZIuaotMHBe5HF+bkYoKhWrNJbgkhTyzb5
UE+6CR4miHMc9bGUmA+kgNgTD3gTtkZt0bzchnV8KiTtTCdT4QMKai/3WEF4
cO+Nh9Zex5Y5MwrPpu//PiI05Z65kkLaaUgkKZMIXU+R7hCm78G6ejfsB7Of
ZQYmI5bHpc3/a4ZIpx+ZKQOVpHQs/a/8f2e9Dx3lq7jTxEcnzDD8VsbmfPSm
u6+BhGYyfzhvHtEu3OclNgM6cGih0cLeDW/WDMeor4GFFz/2p7/Yvwf876v/
nHA9BF1jo16FIQ/quHVuiCoxsj2A0l2GQcJ3wKr52o75+6LQb+sQsowdPD+n
29oTfZCo+sed7wJBNBAMy4enVPY88lo2OHLxb6a+hc77QjpOcJOb+tOUKGVZ
nqrtNupN+ibk11mW6R/ejqwkU84BRQDDDB80qRP/AUG6eT3V4FOpJLdq7PNs
bMzBHEM8CUdZL+UjnjbFgN3mjeHpzybHQaPdSY955tVYjPxveoWBEQbc+LT2
yp9K/T/n31vxEVCNxFCau4gkOX1tctyl7Csby9t9fmmG8ALp6ObATK8pYMNI
vH3cHRa71TcFQsqu7BuQkxrXSf9gnYJMYOXBL+lXWc+VgzyU0vzVzmEy+ygS
XAeeYJIDnFZdRnGTFFV5oqjXds9tOuRJ8t+bg/5k3GCJsWxFZetDxmzEYFEA
VAqJigB45Ob1Ejg+t8fUdbKG2FkUWm4ExrAPErekzq2DlNH05K9/oJCzp/Wo
yC58z6CT2mLcsXJLuCqKsAlrKibS8p9LoQqsFGBwMlAxqmWEzO4WXTEdlRej
z5/6ArMACEvPbmFWSOj65nFqE3G0f451HgLX6RB5tiw+ORURFr/a9RiMHp68
uPdMHqazz6MuA5hQLtOcX7i6t581qPKTW7gtPncgtmeacc7OGNSHVk7XZT2c
Fc0KNiI4zmEQTDZGVqrK0Ey8VzTwt//kZCNdjPpDZJfQE9eAlmkyLKM3Xq9v
DyK+pfe09U7nvFClOqMGt4cOP0cIrftz398R7iPpiZs8H8s4LyWPHB97csea
k86Tj8EUiBxjfuha2f3jhoKF59R1KfD08cmp6gwES00uCYdTpxOgkIwda2F6
JoCAn8bQxWzubd80Q5Z8rXIAWboT/eut244WFRUJMVzD15cB63MGtbad7lEe
1Lwmpeq+vFk0TqHuv5oUCfTROnfoLJuKL0qDCw8hNwxg+Pd1VYbFNMQzqbF3
sVOHPkrx06mtlhg5pclscyl3owJxs5QumgTWLGackPR/U/4ceis2yrDifeyy
UF1ghKaIdqmdwjgWYcPNbQ5432r8UzdZO9z7NhqeJ9kbXKbFIycNJC7iwifh
MQKgTtgxMlpy/+7s1wvO0vPJCmDgBK4ZttqlcSwy53nbOPgP0WyZPSNvUrR6
AP1blGx9VdBOAz+Cvz/UXTZZ4dqdWOWzABYsy0AdLsKu44gHyPghmtKqiwQc
sJa/Op4sxqh5tC4rboHWno9Kfr1OmTtNknv0WLIR3EvMl0Ak5UadRbp8NRMK
vLlbKf7ZkbXl09ooGyA7Vwiv2ciSN4bLv+VIyn+BlorNDc7xW8nXczI7pfsc
+sQIsmKpeA5OjXA6ocTjAq2rtB/cFPuGt8dQbSdxjMd52OStZXra6RmZLBmz
8pZUWookjEUhVohTAoqgPysfPw0Yd8/X8Fhjdg60v3v8A/O5ZMrLiW9EHNWt
fWU4dqeYA7/u1XiB1XqWapjnYRpDyIrVdSnAL6l3nAxO7I+XSnFiatFLDkzA
wbMzsmt8PEVSOGJFf3ZEL4xx9TKwr1h8RB39rlDBYmEcIMgybv5cCECeQn6h
p2Z+38FzBHaB7Hsb0iFceiscAAOmEdHfqOCN5uw9APlhv4utyYAKUxwEkF/v
QVxZNCeI08NAyQB+19otrYMNnyKKjL6zR9DCBIQnK4wNJ1tXG3cUpAUgKzQR
l40HmJD26gwuHc4m8wzg3fYbVmfEXEcuGUpSl/CCLZqpkwcM5L7/2ZPWKb/b
1U3bBkRpHvZkVa4EOMGWPxuRq2Hp7q2x2JMqQXKj6UFs1ZMnp5SLowUl1M5X
tTbBMzAh61tcV4TySI7bxmbNgVJbQMHHZ6eUxbPrbvgPDyjxD7qhPetZkYgX
HLYS/wO+86349ZAOejjzgp+UyucpicnevJWlugOehDIjX76cfBoioAmWsB/S
DZvl7Oqu4fbMXb+9iwGuKU75792a2e0q80286cjdObA0ugJQ4I68g/FdbvnQ
zV53enzodXUPWH6caQbgxqzEnHyQUsocjKki8Wjf9id70LO7AiRnbGiyxt0i
6UZHIIjYeUBy/YzI+zbxpUATIddt4RAoTv7/NA7dcmVBB2O/b0IPEZyehZ+z
Mj//gI7j60k8d78IAe1syktZP0Xsh9LroGMr2mBhQiEdpKGjx8IlkWXvDMZ7
eC9z9bDOYpQgcOULK8Zt5fyEM2fhKkXs5vSROQ1P4i5bmo9G4REwI3jO0m0b
4h6gF20QkLfev+3IH1B7IOpYXUdRzeK5ynNV0dpirAJZckZXjN0sSAq4q4qA
BTzX+1DMkx+ceocMt1bSAdd1/GCZt+PuZ7G4Ykj6LphZpW60WgnJqKl1IiHQ
qRYCCaWfQuDx6+63uU43dTKmWIGM6i+WG+k5DuFcvszqKkm/fPG8uDAkkk0u
T5TnDwrMLAJBbEYhZP3yuL3KzMkV82qh5MPBEzxlex6c/5NYvp605r9+PdqE
o5aIgloj8/Loit842UNWe9xG3FZXOWExr0lpZNm00TeCWrM1aags5d1N+kiD
BFEJucOEQGWCmWVaWJ36IpFqAVvN1dSTmfdzScMqwId3bmsQNvZ3VJXRNn06
AYdZOe1WrIl+AwDAWZKPuAjeC7wHEMRWky2njB5cHsxsIaNJ9r68/krp+ZM1
V9f3NyoP40oJxRZf+uvfcE3+SzuhFrlGJfkOX0e2wXoRWeaJj/WBiyDTNZzB
9Dhi3J5J9xmeBzUxK4hLqvkTjeB7RSNpJKIUQEV+B7Ji6tEIe58AEI+rT2IS
sDX9AnVHAYLOPw1NrMDgzhk0/I4gUuxbBjZl3gPF0mpS1yqnxn5Lwwn3AW1t
W/n3veaI3DvOsuMAhZwdon5S2mZEmQtE673RdM6u/ndF04Fg9ylZTgV4WbfR
/XYFYiCFsXivDY47b4zjSTr2Z6ZierSE61FGYGYfdHpvqHUnosf4CIs0Dwp3
62+6vTMWJ3nd0IVsyvTRgcPK1XBzP3DhzbH6akkF4TOR5y4RoX+PFcYI2/S/
mkRTEspkfzahy0TNH530U94hGbGxuI3d+Ym7+68/1aT2URsMwyFg1LAUrFVX
NFrTBWzhPpILYULEBmQu7eMSMxXdV+xk5zFL29xOarazH7/2fA03ubK8FOU1
zCRdxCRGY/9QY3yWnbV5K7xWZmdr+Z9m74Li2CFjVF3PeF7UbGa6nVOkE0TT
2U3y/Mv3yLlraFQimIOBFPIXiDTjk/9ziwc1qDX/Yb4x0bskxw0gZFbCyHYr
MUcX18lHOPetN1U3/QTibJQzKwp6kXsN7mPZdjmWe6WIpmTUw9gM23zz1n2z
RLke62nLCAy3OtCljPJs7xY+ddhet+Ya3OGjBPSpM1s5vRVrZS2vg1E7qgme
eSjkY+nwA1slUzQkszmBRjC4k4+ShZ5f6TKIV8eKB37PQYR5IqxA8Vrj3E7k
e4M8PDU0CKqwyGR2w8/ffp7APRljm4aNC7dDFlTIc1kKYWm1uS6r6Nnbf0d3
I/WRTcGQk2jTz5MLQ5VMT+Edf5sPdf4UWkabf4EtSw5V/ikxMS0ekwPLXd+q
LLpVKf+K0TS9yZLJ5hnqfmKRR1nnDVtzJ7ZkdE8bpmCtnVmFp9gEDqXv49vs
WO1oYmICac8WfSe7Wea+8vNaiRXzAUk/0GDw80AxAbvvrJpRF693ez5S+Lkb
D3YpRWak1/La8bYLWsGuCjQrWqOeIAN1FUItIFkTu22DekAFyi92/Xz+Ud/P
xIKURDFXUvyO6Hed+kglxzQglqnwGIyYOYiI9FiTWL9AuaUMtfvv33M7KSOM
64uScilC7RXwu1HJkdk6L4JZqqv4xPFiYUZbkM0jyP1CZWeWG/gEsQ6Z/lwa
3292/fGkuvMDUSxvQixcN/CnMng0lgAX2qG19c4VLlqNwybFtzDqKc2RjiVT
+8XYt50B9O4B8tSNYDlmw3TB9f0kVFpZaFmo5nko/wVWU553ktu/U4AAZmpI
NQ/qQQiR0jeITmTls30eHRcvDsTUkofe1QQJ/1i0Xl+uVgVTuPb6SZL0FVT4
GYYdxMV+I6H+0+lfk0hy3c0B8D4vLiqlqM5H+bt9OmMlB6sUGCgw3HskKmIo
oEBwg/f3QF8LuiINX7MRYLonCU8rL3fPBeXdFKaXk0tWz9HkWrdaTYo2vC/k
QRs+EUcJec7L07XSRRk1V42i67nkDMx/JhoEHU3sJC9jQhPJQcZNRwyyyi35
4NyxvaHk2hh6EtMzYShqnmYIgw6U8bpN77IT4NVLabGzBkZE7m/TbVDqo/oG
3mWRmzx7SFKE35Podvba2VCaNcsvbuvkpITP2Yp/rPaCo/yTsk/x8DnCOz0P
Anx0KPWFtZMl3pa5E8T4edL5z9ORBZlA3W/6gXC89+bNS1T5JZot4S6WYF+d
Nyjla4Madq3mye+DO4tRjU88jJxlp/OyP8wmsQXhOUdf9QAmBBtU8qT/+CPZ
VUgUlM5fg16D+y1qxbSM07l3UmA/HIK9CrOt/kB2nKquWwub1vlUxVrM8//c
M528d4UPJ5Taofo/2SmJMGVfYRSUfgDVcLvSXtYSVjAtwKu/IJeabOzJTDo5
0gWCVWquDKBwN4Q2slW9FJOJreZ1tywbnBBe6h2e/Dls/Ap/0yO08tziScns
k5KXBfD7kZDJTv7Hw6FbGJ3YpRmK1AMOnRx0E4gkZGbyPMDVND/eY2RxT6bO
BJGyfEJeJtefOO2zYOrjg5X/d3L6eNETaMuCMf0yQO9B6aXq+UiiuEVyVxhV
bs6l95q1ag0l1QIQCam1ljy0aAjvE1Lj3LTsrdnkH9O7VIiNACYShwxZhwDY
0iqG+6XfGa12sqiTJI+03Z0ojwB3A1TEbzioxVY3RxbC2n+g2iEzlcy+DODN
g9zmjyMqDAOo/+a8+K1fliG+Tkt85tYWKIAkTxOxKjipJDeG+siVluPw5hOK
foqjkwH7IRRVfdnc+Ml0EtiVL9ndz01z6L/l7O140ys3tq5Kpe5yy4xxWghY
fEXHLyVamBOD3NZQNL1hW6CRGjRBh5CkKDOMrb3m2Q8ozpfGmuhJlZsBWUqR
JbcnPjm/xkhIkWlA6MkM9yL8iv8Qh7k7MJgTknSnGGvHxndUOca3+cp+J6i+
ud7kTt+mII7nUw/VUs6lGEFcRZlB4zNLlOMa+V6vN2fRPD7hzzxuc+odW4OE
FG5Emp9ycSjhbRiodhfZaHNA1RjRj14wlGFLtrhwZcXEyU0f8mEN+7HCnts3
WlDxSRzf8Z/uvO8GxehfEx3Kfnb4yC1rzGavV7icjjAhaE6WG3NeJaFysxfA
xTp88JkJ/Xs1LzQo8eZQZNkX4QFz9SN4bnJDXUl8S0k5f3IhUeYeQRsKLb0u
bNBPaxaRbNeJ934FefSsS/uIM13H4bceanB4x5M5KXKlr38HgN8rGS+UQG1Z
i6ry5XMGXNYlbNn6U/H09C/i01QAPOROE7zZvbdLnp/s4jmnngZ8i+xrCt8i
JExVrdTa9QLrrhhzLcRXjP3hrhhBye0wLQL0blDayHVmOZz+LqfhQDb0U2tG
QbH98u5hwbrod9q6u0sp7gaaaJfHuCd9GOcmPgNPRI9XWIgW5gIqj05QCm56
NnnV/Ws/XA68z+vmM680X9UrGotodZ8OoQWgkhZ3swrfMpBgUMemoYaa+roX
LoOh1PgjNNhgv4CovVjrAwBfBnLW8nWnRZSsq9/C1itzpwtE8v7CwaCVKdU3
P9WE57cl/sVCeO02reVuOHpqXr64sxgKW8yRS5tKOIb8atrMd4p/l+2fERIx
sVYVKBSbnUW/iu6c3za+5gmVb7hhcH0EYjl0MacjnFPYnypqiHiI7eexytWS
gzZYNYMBCwnPCc5itd0zhU9U+Y5x5MFXmsn4VaACElI5li9vc8MGgQmrrerC
IMvHR9VVDFZwyqD1cNM43cFUnZuwbdidyXcme0Gyq+ecOU4uEOFjY4oBmN0t
TmMjsAuQ6o1PCjTTyCBWR6icTQhCChewXDGfL1rTHbPkHVM0GfFmCKF4sVxZ
kDsJjHNKG7Zf9Wfh8KfJeSV7/losq1WDCv+fdIBe6csCCmBC6uWxwl8y2B6P
yvV2JPRDnQKUXGapRBV7U8qC0s5D5AGNxY6p5M1l0LZ68yUwMcjNyGdFKYJL
HtWyMQvjbUT/rpIS2baQCW3yRLzPNV7erBnqNVQd66vG1EZRV0/cJBtaNxQx
6FZgByRDNUfLmCztsY4dvtFuxNHkV3B6Gl+HQ/5IUpVm4axw+oOM0TXJ9gd8
a187dsMOhKSzAxwX6x9N2jgriW80qnV9teqHTfsm6hi5XnWJl4NiLCaWaoeB
t9zhYFr5iWVGn0MEsh2sCopc6j05vYI6LMNUdQGZ0buiU/FKRKqyFnLhPDz/
sZXOvAlSWKqm0TMg2NscH/bYSXNWrH9dcO36FAQyytZRH3zDR82XwZmSXXCp
Q4NV3tEJgECPdRHr4qEvaCokRAALgwPbDNZyggEZyWN6xk2HtwCuS59C/LpF
W2TK5iTZkHeh/tlZHxcooeV/PhUxc/FTkpGHfONUxTm5OOIbMDTbiQtUrm8w
H5dSuPRuVRVETqZLybfSNQu5Ak460G8DCj7X4Q6EZ8EeVqZ5sZIOt4VWOfDf
D/hUudoPcRG/8jxueXoZrdWTeT3gihDKsMlAYiOKWQ8qdCry6uEm8avKzTDA
62wsY7xdzz8OnNwDYo+YO6vgtbf18V+u/yspz8QRRhhQ8ktgUF/y58X0DPY+
T0Dkc/h5EWKz1r260z6Rgj3MO1mqPpYEBGsgLAu53q/FWDmQSgtv8aVrvsrW
XX2C85IQpXr4HcJ5OOtxknsZlY6x79pnRRcwDX9M9RO3JUVjqf4crq1VX34m
u47gC2pEwzNHKTchdeiWqV1YqwZ287YKBhxd7Fq9AGDXndKDyxTySqaleonO
jMd/+pXAmzsA2QPpSdlk/goW78hUqto+UM8/6dJSQ+MSLoZgyEJ9XClWQF38
upuyJhGL/rK9beXvXU9m0mg+eF8uNxml28VS6aRoMkzLUyzHR8hvXlnJbSCZ
X6uaH2Y3lSIt/pRoMWFjMn6bY3l89nkGmRUuoOFVeAVTXOl7SiJGPJPS+nPN
z2nOxMtpUK98P7Fd/Sx+/RfQYAmqT9Pcm4yIyPaL/8La1wVkm6pduLgtbPOs
qNWmw8NYLmTq0IKdbrcxv++FmWo8LU8hNdTxj/ArDakT/EWMdTixz8bKPul0
CMGt/p5CCCkeK32AmedAH0kiePEjvy94Oo0HTpwkSRHth9abu2/a7Yovc8QU
8RPx3nGOfzxGqowUsk579WPq09tKBlL5bFLF/TUMhyevPi3fJluuBTjAuaUB
jHhUvrA64aCWoeCIvJpYGng5hXadCqy477hy6ykDZWzS9YlHCoQCDU+XsHR1
KC9jnfT1jtBbYAOYpIu/DYKl7JI+Es9f1kMAK4w09A0L5dpvxEh7YBn6HKok
6ZTkzWnsPYBhjE9JeQr86Db6ABtvezp96NxAVjnP5WcYWqlG22YlcXFRjWlY
c+qS7j4UXgcJxf6um5WMtP+hi9Dfu8yyxonkUxOv9hjbyaQnxpq1BW6EkJzh
Yj/Vi5rRSCPZ+Vudh+KVekdJfXWLGjXcIiCQY8kC8VwM/HDN2x/xdpxQhyeS
mx6fR02KXVRIYEZasiAH4/cIQdimoAapNaZs6bpQL41bt/Mbbl8GSqHQKQbS
WrQJ3t6RlKTLu4VUnByP9OHl+0aXM3/aIMGyBNLX3HZiN2K6LEbRtbpC8yKC
GxIwnVPF3xNHFWI7tkd1RRCnHZ3dmGfrFM1DgInusXo2OT0nBq5FE4teLYNU
kGUll3LxeKaRL8BgPpKMtj4jWZUDLeVNzpTwmL9OT3PINcFzdtRbr6eULydM
yL5MuVDQG+sbr2m4zltZwK0iKloLcdT/Al/oCuKoJnCAti/Y96vX216930Tb
Y7WYnTQeW/qKHf9KInABF+lepGxHtoHIOITCT2y5spW6jMTUKz3h8g8Twpc3
vB74ZvKPlocZniYIhJVzJfncHUKnzIZbiX60ICHI+1V3cnNDmxdryIiYvt+w
DVbEdy/h1UZNhA7T1G//mDXHi0GrbyNbKl5U4VC1Hdjveugs3eH0v9WrbrJg
5t51bJmzgaWDblBlpeNrp19WoAf5hk+j5yHSfeXeXc/wsN/R7upNacSuTJvN
2hmpAmZimDBO511lJY1d+mWfFbbKgAT6giCGB0byvqXdUiGNGFOxVCQn8zTv
WinfZM8ini/wWQ5lEEU3YsDoVAiH2fk8RoUiNGTR41bUgWtuKqQYb7LTvJXG
phE8/HLxATf2YubDXTHH7SPb6UHBt7c45/9V6wYu3Rk3JOLIe2mvlxlb8twL
jN32GslWbgIGOarmnBZJPYgGP5VwtNKQywaMxXcIZQMFLhN7WlNIuhGa5mSj
9qqx9zDAoTgTiL9K1vtAVjA8wlzwDQmS0O4Bd1CZGjsfHcEjQ1xDd7/APojf
3Fwe+G4NS+gwVHj+dIEQ64ExWQo6p1vKM6DPulDyii5UZcrT2ZxjroM4p8iJ
ch7d/A9l58dDQuwkgTzzy+MlwYBLlL3EjMd60Xr8VHR6rn2BKvXva7wNI3as
Cjfr2UrIAfFgv9QL01nL4LzdanwR1BN1YvMQ9AbmkmxzG2ubdOIjvFQpFg0Z
p1nCwwfr3NiEhSAXUtQ+w7nUYspgWs+feeDpP0Im4MZC7wWwe/npb5sArTbq
wEmbuScLKLjshHgMwlZ5ncfFqvmfYiINRFB5loW+Es3OL6u6DSyTuXMoNCW9
PoVFGsOvjSFcQTBH+V9j60G3pK85TnkzHiHGed2N0FF4TFbXQWI1blDX03tX
ZKXwhcjzc/LCQjecAAHv6tCVF19WOMSaxuBL0ZUzHDTsn1jrSRotmr0H6bFj
VMhhx4JK0o8xsT37IBdOr6kP2nXAYjs8dgnUxk5cCAVfbhmUI4/ypWKmglcu
mNapso33fC/c9yyW0MFGYtNXVn9POa2ribNgKCRv2jkggwWacbOibofY7I/2
AGXwHDBzPb8dzsWaQUvjmTLDdpJMtg06fk2yEw3HYZ+mHKhut4tZusZtcl39
JZO7EvGkG4xhO5+Hu5cNfQyqb+4arktSR5X0WPHu6FMOJvqvnWvAHXbPTvbs
okVHZXV7GFp+KjTifg+gYJWIea99BCn7Qq0nGzDofWODVnzbxoQohAq1t7r/
4ZPLA/Fqe6q/O8Yky4mwMGlwJYzdXH9Mzn+/PmBX1inOfLNSaisJ9Ijvoy0w
ba1esprs6tdjf23KsC6xpv4/4dNx8gPYfh1sDQPgegiUfyP19NGbGraDV2W3
knzTdy/ZpHuSbI73CVcHkPqHiBeZdDKA8zKrJDMNo0pwBm6eL4A+tfzMgIDT
kOxlnx2GJ98iO6nPu9MrusFgDAA2WaMcIUDMzDuFDjk3i113nRrKjPCyDIEF
0DeG7HU1UhdmgRpBtetVjm+1jnooTgzXNHVx5Im69JpNyCpC567Rgy3k4rCK
jyfeqRbBBaKncpf1lLU6Prfz/pQWUSM1cgNFRO+JkCH3AIA09xVYN7SwA/VU
4nhXgtvUGVd4t+ZxjAGSwlc6uy0ZQnT7lJap1lsVq9OErbvteq5KXp2DyU7D
9ODtqsN02YDNP9BiD+aHCSvQyYCda37G2Ed+etLPXPytU/Fuf/Tj3/mOMT4S
X/eYLw6dhKPI098y1C/SoLhkFipiWRtp5Tm6QXtb9nPPklMP0h1x0t5FH733
sO7YlY1kqp6J5KWICyQCIkv1Fwbl9p0x8SkKRgtYOGOY/ykkfyPbgdaXV2sM
JG/fgXbk0sg5pvlWvHnR9PTJEZ7lz/v314/RWfI7RxsXwqvoOr7hOZF8IwGF
R9YXz5ciOm1kpjMJDWxz9rDu5b1+VhqNfLWmOHwxkAY/BdFtEkfLjFQ354GN
4uQxNZMXjpOChkDlidI2/SDvuXnk+PLuyMK3cdEhNh75fZk0tBGhNvDlF+DF
Wjf7DjAD1FUiQuU4wjg8HgxczlCyRE5lJhIhw+D9QkIEUUbWf3QWVObVc+YI
WlgjHO9MV8i/qXJod8cuguuzhe9YXP/d5Ff2wxdjN/C+SNifrA/N8HQcafb9
RRR0wDwCr11jg0JdF3aNfo1f/NR2JTKhHrd2ViPae50mULo9k77/KeVJkuHD
3xZ8W7P1+TI4xGJimKsAujEe6GoGDy7D7cVC1DUcrz6Dl+xKQJSeBdg7oTm9
SBCgk45ctifIImztmMCwvI/HB9IIBxATxBGP1zRbCKjsbIptQHdJmwyf9Kyn
vGkuNqueV37vWVlZefBMKBwSqM4Cx/yzzlRXUlcu/vhoVPNNWlp15hkGzHzY
uQCKO4ZR+REc5Pg8HH5qJ2XmL9CkSTEKqbGhklkHJGxTCswNHwBWWxmsJGVS
hSPW85k4/2skdxFaAE+tSkga099EQWXC31DDYhRENoMhYa6lxyMlJBHIUmkH
RcvvT02EJJ2KIywiVVEupKw1pHWrhPMqu9wKFXn75CMv9mw/3D1qhv+JX4ZS
A3Dl4CmfeF5RoiWTOE+wF88fVXeQy3PvWZ55NZad8bPg2cltFos8slvlUpUX
iFSqkL1kVdeR/JZ+0Aj/rJL5eFDn6dfPuCGhUjaMmAZobz1eFZt4ARZSdSCL
RktOMhQpIJ5S637gL68aiRsqqDdeq1v9fqv3Yfxwt7UiHpTT/DhuY1IBsS/m
qQYO3toc5S73WmLOCBJHCAz7VgGyTZmNlbzKR8ad8CM/I3qNJ9Jo18JMY+iI
n9nDtulAaFPWC+hEkXhOeiVzXzbQiwDauHDn4bbf8NKuKmVwHBCYGqGH/7Be
fbwJB3qCD6pQ0yFGRRp5c9iJA3d9oTKHiRJJefWRit046MjQrr0MCfpqlE0Z
x6jKYtR24EfGQINsjvRzl4mlGBgazA6FxQUNnHKShOxQ0FB46YTCVp/FnFSd
KCqJRI7bJYAb3vKk+5L7eDtsS7Azid28hEjcPJuPkUQj/QaI0H/K/ic7NEUr
57DXChRTh8orqVdASFwJB6xYoqqYxwmrfvlgLUEOHfmgG3chZVd/D/OUdnVS
TFLXTtHsvYNCdgS84KjDN7mmozf1tetYmnJFN+TiCzGoacIvCfKHwSh3mS83
uyjHr/NlJJZpa1GYAT3jWFRRcWTuYiALt75QhL4DrIlZrSkEwjXgJF8SI+NC
FHaubBypn/rhGTwlmeczMo4npOH2g66GWEz3vizEcna2YVaVa/gqAGFfJsn6
ninPRLmpx+zlu+nVhgi71RHx+M6vaABVPgfgRnlsYqshOc9wfVVJsekl9oNE
BndDN1dXrJ/kkFWICD/SsfsNIf7Qx0OrSYUnpbHxGiKOaSujaa4ys4ZpqPik
gRigZVKfct8O1vkaiehp/iMxXrLhNTMz56FrCuJRWyv8RW8DNpLyrWlz3lGc
e640JGbbUHan9/KAOo3zGdE4P0E4rjiDr3fT3zWnJ0MMqkL7epPtNkJeCPVi
YlIBKuVf9affRpUunf7cbMz8tUzB6U8kB4GlF4wY7QDXdICvlqAn23/HnjzV
tFasMhRN1cXpUChJ5MMhdYr62Cz7fX7F8sFkdRn5WOv5DCRVPiQmOFjfMefV
xq0oZRWGSz6Xfyp/YRGPusDwfkwytwQrT7kc727EC1z1lWgKHAuG1ddsQzDb
4XnhA1uqxmPB/RE6

`pragma protect end_protected
