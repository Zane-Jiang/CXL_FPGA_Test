// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O8kV0XH5rrxHWw8fFNHYvMpgGkPJta5jTbtGTU9xK56jVtmrwEwbrWzdCXRD
0zJitpyy4hSaM4r45CaYB7M3QgJSj8Bw5RsUpxZhVq56OgPS2GCpYeyDutxs
r87+LTFXl3EerBqBoCF8+rnpWkQPde4/jUUdefR9bYEECpt5I/6bOJq8maSt
o7JjdZ84Z3R5aavygXUoxdP4jW/5r7xZHaYXclzLlIE0ska58cn0dS05TswF
0Vf8Zl5b6Vg9wW8lYrjCFeHCWDJITaR3EhVVq8BFHSOwZy6UYUA3SZ7AXSfK
EtwNCXOZuEn/l16+SF6O/D8ZDod11VZtPN7LttCrHw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jBBQEnZzANqlyE3rYR32t25IAKvLmu9DzMq/Hk1LeawDfAHB401iHUbGk0IQ
lEhm93sXHuJolwB2dbpaLm6bl3BkoxBpdNWgdhQ3DBXjLiRJceer/r3HqsAF
DIq4nJlE2uhqQktVpTO4Z4e3qh4TzoODc4f7bXARWTmWmHdxaMzU8R8PKjrw
HQ9WwaVj1zEI/VOK19LRheYuJAqiAYPYOaEnBcgAWkrVPptizK3nsx34emB7
XHnmsLW42d9ttEebJjVL1iwur9WH1bozDO7TiwZxsPaXDEuEPt/xQ8ikZBYw
iYy5gw7yHmo1g+hnAAkRvNFFKHeu5CATSQQYnJmKiQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eTlBV0istBvkUubniYoSjTVRUG78uL/Jmm8V+bB2iDQrp7hdpcf6F6Vw+iDU
VBa5zc5MsMiqksd7edRWqkgCUXXKZ/INbo9dYZan0OxQ5kW57sKO1Q095ecJ
F6X/cvwL6mM6R71S6N3v+wv+LOum+NueotEUNoPRXkwtIcX6mwtOe20xxD3N
+r3YTpasN0sflDCCN9UWTCRA4hm7m1U8Gwmap7hMnPl+Y77YtiD/lSTpOilt
SyhEJV/pBeDp6iODB/AEMbQ3OtNgXjvKJV6LhsBeKR9jYGEtUJYk2ARLLNtP
HDu0d/oHwjT7QrwyVMluVUENj9LSSqHagbuXnsMKmQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L0lF0N+L1adMzLhjOoJaqfJQEaHVyUvXTxB8K9XoQ6TuPX1hN/VIyFOrYIQZ
R2IqfcjP2hra/BtPqZWuIknRLN7hGJtlIRJ9OhyLqbGhokdUGIL0Z7x6AK19
el4DQ9ZgWmKQFLLq0fOv+2Lc8+NKcollZR21y0PeH/Tm0RWk+p4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cB451V73byyQBpxPmov0vQqiN+uKB5CM7ImHfVzkmc7gt7Nh4+sqPVpTpJ7w
bVlFgwqkC0ETjqb+m3PkpzsP3+ZwEp2NppiaynryGfgh134GCmcPUrHomy0/
5tmdab0mcyCqdc/8OnFthwykmr+YEJpPz80TYqZfErL/Hw3ipoH6DWBKDaDq
CSmR8sKT/V2NkjnGS7Ze+MHAxawCarDdMzZl86Hr6OAxTW4Y2CmT/dcCLpbv
uoNBp2OppjYz7cJG3OfIxcVhB6fRTjXVtUSDlHYPn/TODwyC0Uwm434KMBcH
AW0EbEZ6Q84gxObvZbKHAUiUzS+cz7g/CrLFi/CL9Vv5dzfbP51VwtdNbELB
2AUTc8o67J+Zrvodmxt/JyqG/UV5zbFnqq8DtuFQELPVg1IvnJ3Wc9gPlu82
LRoar1rTu/brN7JRZ6e+wsL8ld40fJiSBHFtHqsLdZE5fgctWQLsjbDTx5xL
99KSHRP/8otLKqvfBKcMdeNxki0WRWFY


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Didbd0Ce1ZReKDMcmY3r64+yHqmXkLiyfsmmpuMiLfxOWl+1bOsDjgkgg3Mb
Ifk+kMI035jOq0Hb+2eZjroxV6P8w7KkEGJOuAPRCvnLvC5x8WW2QxV6LK81
W+2XBsognAs0u4v0WFQ48CNqjUvaPte/GBh/kmQ3JBaLWafYJyQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ps6eZmeb/fY1PLUpHxyxseEzpUs9KjdVgQn7UYzkdPfrnkC2xqDltAVd8ELs
YZALgB9dMORzxce7L0DCTVCC2OTJs61AX4JXu6zuPmpUiLIA/Nby1K2BovLY
UMy5u5wvr3bnnYQSWppbYM3qrEp8OfdvU+WWdXhdnPAtxN6OBqM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2112)
`pragma protect data_block
zRGra34Km7VSmPO1Tx35aed+YBPDcjWPitdhOZPzaaE7YgBQfcZoEj5hNW41
6DMmQ3SKQ44X8jQD6MvA+vcncBEsPMMdk3tW6kPiZ8jCwxFVB9i/Yeuyb8Yk
luk5wSEAZmxjGDt0hoqTAxlBZP0VZqD4QbHZCX47rtv3a+yZqLH+kPmIaffc
ZbSVTRy3pk21fgldv/C/n2ok4CYMxQjvPeNy79vjs1x2EL5srRare+HXIkwA
5QVhuF2ja7GbNA/NR+AAzQKSvd5YUI4v/OQI9oSDtJzi98gnF4+5wm/9uj8T
tryyxlNKOSVXnGNIDugpRjhnu2o8DoIDtmAmlC0YFmtCyCl65Wtm6gg4MMAl
+T/G36+U8n9EMaf2IIC6zViwCZYGkoizJMVLekkYZeo2ea8ewyyl1o4vTnuY
morOEI2xJdL/Yinxrh9LLfrWzeeW+/03bxhqKfg7lMrfGB701taCHmaKZBay
muhs53hRUmjZyXdVMOWwvE+mpNVk/v4qp3kJClTLE5eX36LZM7P5mRsBiZZS
Vmq4aG/9fFHpTDhu6cUN+o5NXsaSTzx03tarl+AGANxTMnkd7Q2L43st0JrA
r9VRcv/567Q9Vdq04nw/MxyIb0TiDmdqUQmphgX5bqLJM3zwjoJOfmd8Z1wy
d65kiAC+DcsSO3t2fuZGWPFMyI+xoJMwr61B3h+dIDlCpVGPlullP7r/XKML
NPwfIRDGIE0p4kdYI5omiB9HAJvMzME0A7NFhewTB/g7UXYe1fqte4FhjsjL
vm3J4vowira5NwkrTcO6LcCTey/sTU6M1apQT7Q//u0nlSxhWwgulJLAG4zv
n9trAvmPkGdNesL0RHos+c+O2e06mb2TKSPDkLG7cPulwfmZvozeZ8rkR9rG
AFwjysP2r/E8YjqjJi+9eoB92GUy5D46/K7pU6DuKMtXBh9XXhdl+oWT9ATS
NyL3umg+g3V+SiemuI/LYdrMZt6h16WtxSrKCPW6K8MDSZLu8PWoUe6KDz+H
JNPm7A2YVwRJGkjypStbz3MQ02rmsuu+cvzmN1xlWP/JXCrhejI1J66jkK+k
pLWi+qm4l0mudVW15cdT4oUWM88SJyJPPYmp7n7Tr3DG5CZ8/xS2Gzy+fx/1
HqvwRV9Wss4ZJe3+17RxJSdeWvIQ4Uw4Dc/mueew+vVg644rgwW6C1ibX8IJ
ywVYphsbmRx4+UsQNzDO4cOfnxw5kIe3xf/MZgssDLw/XVAnsXXGBZtumnPp
a6G/HAIkIEnouI1ytXQsB43eUToW9Z5+goar5VFRHIgCppaV9YVnAmfrawe7
EdjQPslt7qIO3CVgbpgmnKhbsbqiT3rTXQn0VPloB2CXTJzeeMFAfuhPgnV7
P8ZXT/jj+J9SfaHKeUNb6jSrj66ri5lo5P2/Fgb4c8fpJcH0jAc8bbFkAnnh
MKWAnCiz/NPpnK0nA3n5Wvpzcr1vjJ50SUsGZECj+E0pNuP316hdOhes7A/v
72ZfP5OLkin0kDF1f9BUJPJ4iDhkDsOeAG2YJFf4qeG3luUhFh8E3aydMkG9
C+1L+Racketvtx08vaVvQPLYPRzbn9ND6qRJpZcrVdmUHrI4wHiojNWjzK2Y
As1Ja7UJt4ZCh0RBQl3c6TXhQ1xQeid6Lw3381PNuabw1oxK9xwuigqt5AgA
yuRl40pwUnEl5arPvnOko3CXQLwkKoBzZ1QHbSpwIfw1vm6jiA9veh00Q8OA
dEGUNl4SC6kXSFnHMVcvxsDMtnti8khpKm5CBIKD3RvizLjKKuzuT0OYR157
vCE+OU2hBfGye1Q1b2T8K1HM9jG6n2PaLISpRCCuCX02++d50Q3gtWGQ0v9s
/WV7OAK+oapfwTMrjmmR5Qm6HUpDYClFqCR9sKi1CuOnlbR3GTxX5MVPBp6V
1rt8xnz5bdq12K1NSU9wwWBmWVlS27Mqrve1V2LqzcV8A9g9fy2RyP2vjBLc
v24Hj84PYmxrokpBH3QEV6unUBzq4YeRGlQ7lkYDrqH40azeKkwRz8Uzo59P
8q5kjjkDOlgvra+HCHltpp8VmSAF7jJTEvkgGE8ecsMfZwhv6rmOKUR5OnFA
c6PnBdiXj1meQojnG2P7qoMZt+urChP/3a9Mpy1TCsJhJFbR6izS6JMe643U
fcKBHHToDCiNQQrjxnLgIsmWJVT+urPQ9NdFUCXibEnxh+LmfD1MNP8TV8Pe
ncYtA6Y7Mpqhv6Ek7zJKZKG2raYcCfvD+DcaFfcLBegUB+nClOGSWGD5QJVx
zf+Y5dmZ6OxmYRyPDuuq637IaTkH3p+DstJJ2VmDZRDyQ4TtTlX6j7HRTPx9
PrKJgfNy33ZTHHz3qccfINLmFmB3E9nT/tlVO6btbXDSXARoxjbTLE35Dn04
iTB+xpIuYX4cOr3NbOrqjYbk8R5ATL3MJ3UhSYa94OtGVfoPAMUTkMnD2MfH
UoXEy4jzU6wD3/Iolvx0VYLNB+v36XnYb3PQvSiLqLDnFF74x1jHcJg0MsNs
WHdZ7N9/rRE2mTKwQNVtt8gU8EULhmyeWeIU/RH8hSXMcAkK+1hdCfK9hkKX
0keRTMFeDB5LNoENpO2JiOU8e13Pphd9pNTsrZLm1rfVyO9XBPo65Dbah81e
yXyxhDoTAwSpvZN+Pu41dZnSkKWaLj3SlHYx+UZbsS5fi1fEj9vTG44KKDeG
gjYg+KuvssWq9R9lWMfYma0TEpyMYyO+Zt2huKxcjCkhoqHLRsQSIWIfE6KS
Ng/74RYw5H8ENYgTPVGmch3cRtXZnQLxX/OZWlfMgWHn1VUbcxzS+cWG

`pragma protect end_protected
