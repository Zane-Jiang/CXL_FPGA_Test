// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1VXNCeBHYkCV8kU7OrRP+EUzKuqFWS9iYpVsLKdY36JIVh0Aj7p4OcDtUFaCE9NC
ma0jyvLgZRKQh0CN/bSFYj7NEOa/DqAvYtLsPI7mzQDlbnZQYihVGfEHnA0THuei
c/KAN2/DryL7bP5YPlRAvJOtMC2ksSfiynWDyAglz+Q=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6144 )
`pragma protect data_block
FX6RO+roVSUf9ny18nmmDuA6MrtzlFsVlkrbbC4yGZjmdUwCHOBC1NMT3zOPUP4H
puLS1lL6nGrztY6lDxAwGkxXbvWCK5EF6ZeXKbuRkeaDmki3OY+rfXs8tDY8pCol
+mgoxDmd6EKdfvqiTUUbmuYEmE+qOsmOcyvbR4Uiql+l0u3xF+mhdCq3P+AexS5l
jRYfNp9fp0haar9cVemtTH6p49DQ6dGNUThbMDSX3DXjkTjO0lJ5poJGlKDLVyTR
1aPHmTe3r9Uh0P74BedAt52jgi4IDtC5iFI8M9kejajOrg6cVveVGdmS9jLnR/80
n+NKupyPXseOSdUYqAqyhUu8A457WNK6rKAWkIPfxWFJkcY8gzMPUXcDCW0k0WP/
UqoBOO5pIa/b2xum7Qvvl0a+fs19hZ+BpDjhLw7Pu2bgOPXwIIGBHRLGF5Fz+6aX
OCBMCvXohNt/SRqeE2LVozE1Uqtjkcgj0oOq05UNWt3eky8xdYiWvQp7HAfurTMH
ibMJEeupHIphQtWEgsY4okPYphjdZW/gaveDmboP4coxJwFXEbaq69uoxR0+UqrN
S0d/p4j3sLe5se6XPBmctas56ez96+m5wwLuW2nZ765j7KLmXNkohyZeDMDtJeiX
kN6ICUj6X+rjnIJh3EgJPaxga/ksf8JSGu/+1M6JgJGlB1o/0pdJhjTubUV7sn+g
UsEBohdcLihO/5myWeq2uO04J84edV8Xm542ALDIHOGfgGkf54b2lGGOknbMqNL8
fBQdv4HeRolB2zgQZkPZYtk5NB8TEZumhYaY6jC6YZ4Vsd8JZtV4sHY7HMKNkvxe
jUgs8YNp7tTD+PzfgsdZ6emZdbONcUFCy63QbS2Vb52tCO/TgwEqWUKez5ZbulKT
ox/V5XSB2JmXyXVcVkXo0yVfQM+KWR7Tq7ZJTy3SZbRrJQHhUi4QeGWC7AbxBKLY
wHsftEWTLpV6RsSB/J8D7MmaEL4gqS7O9Y0PxV6P82LPIdMU6OIwKVL5AM/3DeSA
bFWwG7QdIQH+XyGt+5FPjOmY6WAL4vIdpAtIBDaCeAGB8jOyJVDUXb1YFrmom47w
3VqAkurimTH2JGmWgnm+VKJ+DnTfoLW9fLZOBrBcr/0TVvfuvpgo2Ux6XLGJuzCx
EbcOpocpGi/cWTxDLX4qOPFMyQJbjwGWGXbQ8zdngCQcA8w5OJ1wy2+tiasGI7qG
ZzdxJfZzRUH75SrMPgnsmpT/SdjRrlT/JSYL5In90sscv63tau50585qgwHsVZn5
kS/TEFYaoKigq35r6HeP3w3oXIGc9K52EBdD13hGFM0qhyQSgUKahBo8SDtkHSKK
5N5lfmeIO5iqSe/OKXYW9rmY0pqdOcdzfnKYrOA3POBmvERuHuSY++z/tbAoEGmc
ItPG/Um6MwHWBNGZi0vmN9TQWb4b1m2b1tvZR3xEPtcRxvlRIxO25UXwe4LUOCvO
lx5XxZKLFuT+eB7lyoyOmTiCOWC48YPehNyh9QyhfRIS52x5YN0TFc5J0b3riwA0
CAzRJm7a+1kFmaUzJno3f97ySHQ1Uo+dOUBM96JQZ6t6zDKBWethQDAR9CcVgR97
r+FQAyYMOtAM7SnPAOKIzdrLW65iHBnXUOeTHgGMr1beWLHQ3TcHWhoRrOcpE+dK
USkWviw+hRVhSzoRaPa24eV+x5x0oZzY32MxVwWtUPs2sxrcnbQ/GtR7+uIGbRhw
1km0kJocuymxlZryzr/eELJ5jLagbuNulJGZD6ELgnEu0DZAZRTL/jhg+JZFcJlX
+2sTt27bb/AhMFrAYcmfXjEaN7XZsi4Vh0JIYAkYr0qd1C/FhGw7ecCDnkGAPHAt
G2Pwwq3MSAUkBCXJZ7qKyoEB2IPvEJ+1KKMWvqkLO6jCnK269Bv0pEkjvaVARk4w
wBxpCYvxgObbd+Zlgj/V9kQTjtSh1Yiv9NfSRFkPOaVVx4wAAJ2pAXoTBMgy1tSA
cKif1QQZinv42acYMg5M9Nj9mYPnyOceLpIzi79Z66wmetgl+lLWCULA4d196suq
yapHxgAczgga1pUe7f3/p8qu0JFG1gus9slwnt/PZrCFTIsn/P57OWs731XexNWC
ADro71AxYqC8pekBfVKJHtF7Jo5wn+AKv5Wrogl3laNimXJSZW7P6qV6rTwvOUK5
bpixhW0ceLfC2UWcDB5mj+rYiSC41QWCf9wgF19t29r1/mRhOTkWyLa6c9TJLCuc
dzs84eD39451mG2CZIdLsaxnHi4YmxkRGJTL8cE6njtxRz+NlVw+qsFC0Ah6hwya
XnbsjaX0/N3jVz1aW8pPHsGxFMqWMJdmCwHL/ZH6XPxgzaTVojoKiNmytuOIzXJI
f3tEUAjvbI4zdLw7iZyoSAovAA9uqKzym8hffUiSkEeEQrF4+z3swokpcSzJh757
Ev9t9NpBChdqFLHJ1NTUexwCXC+DJQlCRT0rMP+wp4CzYbI5i+QKG8QSijIcOVlt
rQRmE3Meg/ku5vABKBRqg98qGS2x4FMviY4oxklIDFO51HL9fDlyp/FCbzrke6tJ
SkTRcbFMAwRtta0wlVGPZAIor7Tnr2Fa0kceq+HH5/jsatFIgyE67AbUx9B4qaC5
b3o2iWYPjCZbh13x/LEpsyQxvXifhAWx9h+Pt+d0eT+v6M4s7jSvjy2ZPKVKl+qw
rUKWHw8UENNN/DdeHQtQblP4SFWlDvdJEnCmQmups4QuYE20n08GnwDt0k5N4jB7
e0fM03AN7r2ZtqIa9udISvGTW7uhy7AGpB+VdlF8trg0J4WIVh+KiVQk1D0Ynu6W
Y67weQRkd3CNYU59I6HSMxIhmIiFihlThKLMFc+mOquTBHcCcwcIS6Jv7bDPly6/
8rSQwBaPYlIKpX7X4BBy8e14mF3EcS/CUGEEtLiJI81JZ7P5bYtUcu+HKND5CVd3
jr9e6LNVTjsGv5MkdjO3kWSBjQoBi9KDtVanopwCotR4JGsF9wHNUBfr23rKamzq
mUCm86QSMsD0fqG0rg8Udp2fmxoRzqpWEni5MiBgpQvdsm5cNL39VV65wRg3Bs7M
xi8yFQgxZwor7AIB+3RNFxb4QgNoDZuSZXZ9Sau8IhwuCQrhScRm5r+VSB+gi/Iy
LVEHGD+oJLPrdFoy6qFBVz5wzs3NJQaPBSyPm1xWlBBRsnSuCFxzZyuxdXPlO83s
Sr/v+OeXJ42tjzYGCWEG6jjXOiSA38Gd7mw7vTS/WSKiPXtkejtKoYLTus4/BE9C
J4LQuJAJfpIRvh2IlU7CDcSh55OYh6YKq8qrhS9ZvuPblRdSiiIGc2f/qs5mgvAv
cYQTwpJVlVXBqAgiMWA1HhE9y/FU7aNMO6CbY0mmOLD8SAOeKlrBsYbbSWn9uWUH
Hvx8lvu58MNAuk7aYfsnB1LhZDwoWFnU2RY7PZhTjht8mnl6vaEUU3p7x5NfqDXy
EfGk/WgUVH42Lgxlm8ibPDu1sxF3d79POMlgJitVEQdzNTrQoVMbJteh1mr3hDb4
xSpj+4E0xXlYi0Tofl+IqTKIWymllmKIfbOkPELdSt7yuNs5fKe3uWKBBUMUSc++
X6a+1zrk5fq00363AHfV24beogF/GQ7Xs/JX7qCqLcQyje7gXOo5m5z67RkmiOMZ
6rxVNbxQvmWkbGc4q4ovnKWkkIRLTFZaG7hU9Rwo47x2s6wT9xKyQNvs0xLQFtKn
ypZthlYAKTt4SZoISUaXvdCBjXZw/6lHO8IOw9gwe7qWkDBZFGYOYN2c4eDJ3Yj8
NuzwKy51gZnbcIlyXG3xllbmz+MAzfWzUxQrP7aGe0ZNdGUj9aPeF/9WfdYu82rB
xnCYeAfSsv1sCvbVkS08XyDPb3ZaYUA2Jz5hHZujAqMcArq5PO3g+eQxXkdYu+gl
nKq9LgglyEwl/JiJtvUdaVQcrbWcy/v3OUUbNy94N86MPKjxX0vJNBmVjoecxoo3
NzG/1+E5GRR8qck69RDfUC4nO9uEnlR+D710QGj3XKOmkJ2g9htniFgziznzCRcQ
cFEKcoy3jQqlXzNjDeFLaeMpkv6wA2ByQejg8dGLdxKjzLA40hsgwTHeHonyYEjh
qSfVkVHv0YdkqL82vlAo95l4Hf9QpUjrQOZf7Q12hclJdQBbvRyRgah3st6Hmf1M
UQi2hJG+JPYMgRRbWwsvvUeszbPGY4Qam1gsXSEImVothlGihlOirQqL1+vFFLEf
lOw34DoXKUq7o4i2BycqH4/Y5Qk2yYuUSOFSThdOTdtRufRtPmyR0iiNPlfVStkK
VCQJS7nI37C4fpNKFwA8NoB1oyK95VgHLD7C8oLzf8Sh7NLSBcAp8wjAtahxC9Mc
R3RF08fGZyUvaniGlwPCqZOMVdOatvdJylFjrPvuZiphyPQt3VGipsQebY4CLMvP
/6oAdzxB3bUf5w97A4tcJNZxTiAN1cODm/uJ2LChYQzY/QtZPE39wKsWKFXvxHq3
ud0dULovAhy5F06qP9RQp4J1lXfyhw4lcmrq/uDI4Sl62TJgwS9STPTjsFUmX/IG
cGvFMA/512pSJ9xjk0nWp/2ojM93fitRGFdodmY/yJUoIFS9CnWnUicYOYq+9HEw
c7I2B5MtuthJAcY9M6DbQPoHAsnDpSVG/LUDBxmYKMOrRky7pNExw7MQMnxAHRb8
FfB49AOQ+Ckl++tnVvuBzuL+/kdG0BqhTn8MRZ+jNtXeiSe4nneSexIMJHR8yH96
e4PAYrOewpzwA8CbyzRGB6sw/W3iM7bzjAxzocnaAfP8TF+HmqCzUZEIHvOsc0Ft
VgI6bJAtpyhXey2aMUZCEftElB0Lid8aEDz9VId/9BDLudxEgAEgNeB7FSt3le+J
qIUFuP4lc+V72G2uhCnA5bLU72MSqx/hVHrBDK3/bMCLvVV7mWmjQ4xFgBGcDVYx
MWFaNNY/zbRUMMZSs9jLF7OqPU/t2qx2/ayDvP5HlFtPtC4pMEw0Mwj59Cva7E/u
vrEV4nhllKRZyI87+o6BnMENP9YL3kiZE/ATwUiKyum/sxcKnOdgxO4Da7CyDsjB
eq3tt0e7yUXO+r6G4RdMLZne9MqZig+qoyEdlecY4De3bq+2jWs72/jc0xuN64QA
JzTkX1DJ9MvWniwWvBLqrR3wpagOTEdQjsXtixDBAaHEGb7RgswnPWD2FdFcTI76
7VPCLdn77ZmVPg0Br3WO5wYdQZrgiuAdbuCrfnr1cSzSkTjEytoNz8cbGE6iEoDm
aygrxBGDwHlD1OdHxMzu2hpCcxavLS31QFMM6ukbssFY5GODduszxhIXkjb5fwGz
hnDh0SIkB6u4qZfdRiAZpqxcZ/mB9n++hb1xIkNIOqPjIPvQZ7jS6Rz+mU0FlCjb
a9TGPx6WgMHUC/moowe2CXgHI99MQnUtyRRu/Y+z5ngRUfbuMHqrfeKe9E54LqeP
HB2GRhDoI1O+RdyHh4D3RwMgwHttZT2rxSJDMWMgR/+n4IMsjx7ySD6ESGqTBjPm
ZdyXK14Bml4Cgc4mMm3z9voKTzGGqaFwJcsN2BU3MfzcrKY0ashVs+ID5Co/M0Sz
XCjzvlzo6JnAL1TkAfn6qcywMdM+nOTa4WNDfmpgjOg/D66PT1BrV/NaFaDb2fSj
7hl8sZ1f4Gtu3+MY1LkODUCjXhDnVpSX7pw2nSia7ngBUAvLt6EcHVWhXA8rE0Gs
EA0wJnLJARzSHIsj2lVkbtgrIG5kUVMGdSZmVzDqUcDbroaiEw9NEI6VsXYTvkHx
QHJFpt9PXt9Gp+jjsxuE++YAWWs/mVeBoUzJ9t6fGe0hys6TrsZZSixlC82PByGu
4bSjwXIa5ADRpeSkqZLBF0YtQeM/Fr892hy1eI/qquUbmkMF5AspsNVB6UcI99Dx
FgoqIaO+waBH0fFRwDbXp/cATrTQzHbpRBFQSAWG0S9YJ1qAsU+yDxZaLs5qJAxi
/RW7Wctm+idbfny8MZI5GDkTHkds1cHMrKCykbyM7RSjnkyCA4kWBmyEtAMa43Zt
6cD1WCcwmuVuuu06zVxo69St2CKw9IYx4kT0ea5AZxYCc1ZE6GFAwgIxGuSg2d8f
ZcgN8/a8N4qmL9hzzHlmzYpYn7RjPo9GK6XJb9niZ4qiNOWzD8pfSRWc3BBTBnD/
ksESQBuwTU1FSP6phgPFi06YQZ0/lvzjWbA1EamcbmttnL3xQSLB+I3NkNZCuUzu
aI0sMjQmZnj6KnKdkZTFgkJC8rEn4WGbkLEJpOPw19n9Kb0vhUZUmM5KdH8qePJz
i90+ptWxa16pjqsBUezYYtUfybBPEWneY3UBK0P1/4fJjWzuhMFnKAMmHmN2/7Q8
xMawfyRA+hpaW9PHMy+UM5pMDhC4XW4nOGMTCjPxGxUxUzql1daTC+dWd+I2TK6b
PE2fdhn1ZIekgPUelaRfFPJQDrRfiFFGCOc7sRr//Ds8AtGNsG9e3axDlVNk5p4M
G2S2EUEuBFO4RPs4OMPbG1LHMsn4v1Fw1qXG1QV1F4MwQUf/ve//SxqaSxJZYRfw
uPi3F1oh+EhCQjoUAXYtBAivxiT9jlBA+6wGtnbeGvQex/mClfROKsJYGcdsmTNk
BK83NYFm9+4yBVa+mDpRVYQozoMNrcYZ16F1pag5engkYJRm7mY8HB/XGKUuoFSR
sJFT6MIDuGfIel7zxrjZz6E/CeyjkMMjPCAVT7ElXSgcnLI5X8D5k4gPvI8Vxles
ZYJsLOB8mxdw7ugqqfEJvfy6+kKYSxEPjDrT8pobvBZBRKJ8rGOPG9NBsOG3K8DR
FKQlG3JXOlWLJCnr92IHtW5ZmnCO+i3Td9Fhq4uMv2gv0KIPg+Bc6o778t1JVXn5
XX3Wou37gZskHBP2DVnsjIev3ZCvwW+2xFAqOxulCMyezluQCOuDBLnZyIH5RP44
gT58TI/SmJWAa2i/GLMXjLcebyRejzLLKM6QF/XOkh2XoNCCTQi7bWi+RM1xzLLw
4f+BBCLJoKvISXq+FHCWE/e0s2tU8KzD1+DrLlMjRbkljxU70yPNSv6+aKY2McVK
h3KbF7NyUjB2BVM9r6Ax/xy3En7y0OT+tnIHtBmskJO6T2PNFCFmaz8/8p7fsW6I
m/i6Udq/tfGMCyLVtCF8G6v3JHjRtG/0G1AWQCSA4jcRbtz/56MQfI7p6u7ApyA1
d5xPwXJMsjyErZmKMEyGdc37qpl/J4yjHFGTerTSCvtT6/LhsYdfYn24HuUip6eb
fvTRG9df7LWvLCR/4uhlTP3z2B1zGMMFEH3XFw7j2t1eXCXwugKX1fUfMIZCuya/
VXXkDTbciIIlTzTCaSjr1vQhYiyRvkyQNKisri9EppmAi/614QS5rg/fvfp2a0Pc
E47JywKHi594xZcHXlTeu5mu7L7RDGAluBz9kulUNYYTMsbikFrIagBfnzQvWAJX
zRk03tyYUx2aBKTn4lrbuKhQ/eMwvPnsjYgj2QMiZp0Q2cX2HPEurLA60If2/m+1
+xbW+VpkWXX59RGQnigbpU6vSa634XqRSg9It8j7tiUFnxHqyMJk1/W26u64y0KF
KQiL3VB8SRr8dDF3lcIUTmWK5eGQF+yXhrmOqoAc1topqvzpoC6roid37LbWGNfy
8X+1O/9tLvUFqHr7PUX8QCDuss4C3dIJKQvyRzFCVaSc09Proucpb8V528yx/LZe
vBl7quoVIbNRZ/SZ7JgqVKzrN8PXsKTJk5rozioyoiVX09qCey/sQwE3shteUyW9
vFn42XhAue4ms4VROF4mmvJtGD3F1uJdGFB7Mpm0u9a15dwaStu0x2iddRLPG7uM
ELq+KfWFhSSQBoDZrs42nAldQlDVVWHeoiPxHKVAnwE8BpOBedg53/5reOCTsQQU
g3ELBzwXF4kB5pnOjrmnhC6PzeOBFjKt5/sU2DKoQslI8YEeFC4Ww4QLObgxLIhB
g2HJ0ZqCJVeJv6YTcNl+BrgsfAtjickdt5olMVnjHtJyYUH4WHLb6bCoyBJzM62x
8SSs8zAL5UxsZb3YMzeePSjkXzghGp/wbIKQ3Bh/dam7hjEBbFvEb1hlVD18/dIG
OpHlvjtxSie+oKSf7Sz1/4ee7StLYvl18uvAXwnDOwAFmgLSTAlaU1dfWF9Wkjy8
xhjNOKKfX9PrTeeXYRBmsIXfPdQZhhadW66C1VbFMnioDQ3RwJ3XwGj1rJRaS4ch

`pragma protect end_protected
