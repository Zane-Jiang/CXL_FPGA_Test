// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hjppEFZsAaie43mM61UtsdQKphyNLHTQu1LrFXRGHhvEYSsbPo6i1b8/1rHn
mV6gG7waHMr0s8biyleHGVP8P7dPJ909g0OEhfm2yxExLhQec4DHzhAcPLP7
CL8OXxwV0+SMO13N6CMrihutJC2YzzmMMGns4u4xMkb2IMng1894rwD+0dDe
r0KHfl+pcSl2LmPqv2LKh4aYEqFmRbiP5XbMHZkKJnNf6cJh5k6Df4wbh2Z8
L41DRf8RviJP0f1xXHadBxyX2+dBUMxT9YbKf0W3fW3yzL1j5EzSsK24gbl5
O0Vu94aflAgDkTB9PISy0IZtXK08PvHrBwHCcBvpNQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bOWWeGYpMSNHk+FuW0DLm0rQmf8Fr4J9Xxbpau0wMfYpJoysLIidwB9MhBXO
TTJWMMC42SIm4mi1j0zTZGJO9coFTY81DHa6EIEaTWUbn1gyhi0cXHmcsbhK
HZ8BWKB37v/10GUeNH2PzGswcwy9vXdC3pMqPeQq4uUOmgXLX579f2V9PzXn
Y3tL+/3SCwTY2XHZt+oCpkBRA5gMoi8JCUgzjoexLihs3eTiDPcL9sY58j05
kIuv8wBw8Bx4pDLTJzQ9Cic9nSY8QikpKi20O6VN/3UgKjdg8gUoRhvLA7/O
WRW6vQrG1RqYsFAmJMjMidoZPrXA2Prwmd/3eSyNdA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iZ7fPUfz1R874tuG4BfwOA0fJA8RD0+2LtZ3fXEWzDefIKy96JRP0sxlnLPS
J+F0fZDwSDJ/LkJylaolrO81Up3VxYcKU6xujb4apzSYWKOgmkqd0Q5p6VKM
4IOwyxEiLfLDPJQhpXjxB8/IG86LY8fSob0iM5Lsu1zLtLcUnDmFRazdKcVl
o1ZChNTk94/NuVxKAAD3VpyXm5/Xe7wjXt2Pi6hjLuY6jzpVxaGmDgAasFW7
8r03H0Jyw4YIVhtHcerkKJVO02cD40cQrN+WZKrD0qvslU/GvGKH+Iaxs2D/
22e7lcKK1XNAnIXakA7H+L96qwo6r94kUp8iP1/lHw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
caJSvdbuNVBrTmCL+Cvr9mgPV6Y3wuVfMnqagR4qa4HuGcb3m8Gr2OEcfZsn
IvM6NKPuNbSDYjWXrUGlJPqCKCm4tKOsAvYxyr6j9Y+D6jBKogCjBaVeRZaP
JNSOagzcWXpyxS8IuLdmH+61VDQ3Q2tYF5rl40YFFCK8AuEBT5A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kTt2cw+178XJ6RpPvo5mV0gmPAU0Gyr3nX4+L4nGcwn3yZ/++6rweSkRWl1D
6oFWLp6aYhqqYZr87PGFu9gtltPxpYuaI3cBPX+F8lV2n48Y2hndzPQ1Bf8b
Qt4Dtzxl7I+CHUM8cywaHDd8KAWIcBdzt1R/oixyAPTjO0JZ1jc0/rN7mOEk
7Ifshv98orDQ63iYJi0VAQ4C+hdP/NNSyPyCKokvOEtz7+4SHX57IOIylKEP
R0hxOxw8tPUR2DJBpCGf7dYIugY46vqqY9kuHHRKyHeqwOi5ISxbGmj5p765
Ku88VO2HidmUFFHTB8LWCZ+vQCve8M+qjG0TjZYSNcSfJPxOCt4WqEg7BPDd
0kbjraNHAQSuQpKTngn9I0DtmwtD7bhg2yf29ujkVIOajZB7PC1lJ4USgVka
cttaQxXGk+zufkj5hVvgaBwYKYuNjRgZPZU/dqH4pfXnvV7xZgm5fPUyHiUT
MsxGvFhUIty2pPdUWqeG5IgTajxHAeK9


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DGZ0/HEcYzgMyxXl9k8IN6IuEjI5SB0V9M6e7CVW3ZV+FGbnsdmD+/tAuZQi
chjn021vXMjoxveHvG3TuzFDCvVfB5Zf4rGc+kWmt9+y6dbf76CT5E5qCb/6
/7p5TOGCfNOHpyBhLDuQoBRnYfYT9EIanN/QGe/oGcpZl0Az8Rg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G90nHNYosnNYNdsNCSj3f7m+tK7SKXMErJORqOF6MKqoRVvOI1RvxuyZy8zw
ZVrID8J/hjiPVuKkLzGieuTk9ji7hE6Ik5h08i8lgGrIB4qlx0C2RwJWyiQj
2+jKSK6rflhulweKSfuXcqb1TcZUP9SsXvWnJORBV810zXhgMBg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1424)
`pragma protect data_block
cvxcjpsjHb5/UZp8z/MWDwYU5QioTqSd47P+ipZxVXEUr1bbgIChHfsMWO/H
73Yq1AYD0XVVN8RKGZKYMUNB7gfwnHdgxIWMfI1lyEELYa8lLXBlust8LdFu
K3zFVlbfN+08BTL5kAqhsmscdfVcK69UNDU6zv3QRslrlxggPoECMMAWlIO8
HBDQ+NGpF3wHQg14zMuNYhzh/OtWyjYN2W3pD8bK+hl//ZOpIWwYyndPZQP0
WI6UUCxNSwXGJpdfxx+OIoo1RLtnLpdhaYI65vCgt7sQYOjKCLHjDzlZ93TU
lDHYXDEpMKIot64/XYyPpW33MWgZlZ17Ex1Ma0P9shSMqIwAbOnXFCZrJhlL
9o0TESTFW10ixQeZjqd1DC/fzLq6sYQ+J1GqH4AkvkO8H/kpa8MdPPFiVs9o
owvgFldLtcbAVIhQN/EKJ854JOxeZ2Pju5V9+cAQN5bhyuApHg5XkbqzpjfS
E0DGrXEsYTffm7mIsuxtZP44tr4NtmIqL7VthCddhE9tG6R9aoOYOxwfSWDu
Tc83ai/sn62R2x7AdLvmuOGxTw2CpkEjqdjHaGRiNNAWs96jx7FWCX4OvyxO
6N7DGt08XhmPmrO9M1l2nBF93f7Q1BiJypsBjlUt7jUsQWywfg5Ta3gG0W1f
6euRsHJA/1h41gP4OqsBVdtEUs1IZjfrWsKoahb6yRtE9q6zdWqnhPfZ45pq
vEqmApkz7FeuK18UMvVowAxfv7bao6q/Y9ziWHhVLdUTOh3aPj4lXP0ONsLX
zyGtEiDfgttIzYAW/gpIQQ/iD+vazFGIa2Mrh0l5zebzolGyKWRU7JdrWWoP
veGl6jBEJZAWBGKDVg54awnhxZ9W0s/OM6kLNta8lC00z2OWEywrgLcAwBhH
k60Xholmefrhn6PoChgxxF5zpWSCK3+niR5tb5zD41PghOwyiqPtY4F9DDBv
VzULwRLmuwRJCUoycGkRG46MPEtaVtMvufX5ojteDVmN5x6F7dqu7ilDHPAv
NlIFh7znJj9flEn3wgMS9yogQEO80GR52WnrCAr4h75WUQYHagG5eHc4FQ/T
3DyQY9SVVWJP4W3CXM4REjz8hFAnZ4nig2SIDrY65/8LIP3e3Vqd4ES7cVrV
gmJKqSPPFL03e3AYK2C5cfRgQdUytX5OGiDzSW/rzOlxEHgz2IryB4nJU2Sn
ksVUWvdtP+t6glkl8529fbq5z5ek+i8MDu8JXABeaCdY/9yUbTX+0euhdkEZ
1sK1cIBaTU4WLvno5CnQoOCnHpqZiosPs0mc2mB0DILZodLFH2SltAcfEIHV
QFEmE4tfKoTwD1ZHgtOPTi4ytmWMXyZ38ILvRkndA+9lw519AdBaXJ6S/qPt
w8JABiN28Obk4patXlZdSJxQutUVwBeMV4UBy8pbbQLXah3SIBDDQGWv/6KW
zHd7K6MbuxQQto/kfxwpcaprwpiucvrte892C2LMQdKuJyFU8qWsDR2cZDQK
b2M0Eqlsc7GjAXRUQ6Nx52jolhIiCEF1lp1L+qqDLMritUm82DzefsCSJYXt
bJ5M0YJ0foGLvloXBHPQhz8ca45ghqqEoih6ZCr+cPyHhTDCDhxE5QgbCKwJ
PrS5R8jXyC4zOCqMvA+tJyxqNp5etPDo2FJcvK4ai8QjEtjPuHm32MEBwZRH
In/oLGy1eKcW78tHH+Dm4nSLhS+q+cEWax8hXVz3O82yDnKk3Bqu8Wc7+f+O
klXsqf2GL9NlALf0cuyGuIsMWDGG8AO8Ijg4+/aIc0TO0SoDoejjBI8xOI5h
5Na+Yb3OVOsGJ/n79+2Bqx4IKJQFzSHoYOcmTbx04DmQvNdH2Lp59ENDYK7H
qqLDTWjpoXOKWsIXQUEQMQPF1DTIFDX0/Xq4lCQ=

`pragma protect end_protected
