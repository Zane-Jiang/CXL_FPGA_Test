// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
kK5T2XZ/GHXf6z7KuNuspxQBHzVrroZUZw086V3HDV6dGQ8vzhVqoFdzTchQnqRO
bT4OetXJhkOZp0du83zn5xlmCZDECnzK9MiaMo78iy+2+m8GYUyqCGyxnZwJ9C9w
yeYpssDCKNjKH46MARCeU5tktC41nlxKbYXRmfIotvM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 31408 )
`pragma protect data_block
Cy5VkUM7u5tXWsiemKM7xevhy6AgBGgXtln2u2nisaIAomf26BpcWjCfw2xivd5c
pyhzgu6IMHlCf/SW4UgSu0P+VmCpn36ccxmVeLVlYRmDZNWvQEC3QXdTeD1A/wOC
8PyTzO4qZ4ZPPsdQuOTvcgGjzgWvT5w8IRPIzSb1JwWfBX3QtC9vJpUV/SjBbuKw
9CZF6dyox3NQ+WVzKAkGhaaduJMutkpGmkaivwYT7ksuoU2Shfyr5ZfiBppr/Oxf
Ras+zUx2MHA6ffezh9bozlLY4LmusbwNoQCY8B7hdTuRnRLAwGk+cLCnAvq/Nb1f
Ke57Qp/l/mdliBN9ymLHukqfwzdxq72KTkXP7Rjn9sMP/KMSXl96uMj42L6tJqo8
FToIIdAXnqVVxSJ+rTDFp9xKhBM5ARtmh1ON0sHZ6JaIXIUbo4kWFOEYRolZ2iIW
yUqvQ/gV+CSXPF9QJoDvzrwdyg+KAuLftcA9rdzwPT90bg9Zpj9XWzBkrlrMau7A
RIOt7btuG78BMm78vJp89vlKGqdnr7yTZ5cwYuY812IzxiLwnwAk6wZomV0Y0JpM
igAHxfIVimtcI1i2djMg3xEXHly6gir/CUBMSG6TRAPbfAg0BWaewelLJHIY6Zoo
7PkBi1zrMv4Fd5fv0I7H8uPHPWsJndljRivLkXh6Jm/aAwhp/4OAtoAkg3hvFuE4
Zpo97tJ0eAFhsesY6V9vGqS1tjffXaJb/5yjckQQnE8yLzBFkXS4i0fD9JGSpdME
VilhhO4dsBtkMwSUHt+vKKaxtLR9U4EIkPuxbRoTFBLVNtpEJQtXACx9AClg5taC
4lH3Wz/GGuF4Hb+c9DOadrdmMNA6MrFnfB6wsSlENjkCnS+1cFLetKC/YrZZNPZ4
hR+ssROwIPOgWqp6HrwLjht7P85WLSz/uY68qnPvFloHQmUAgJlBrl/icGF1ijJx
Xp6uq377StITaA7LQ+pyvB9pSnXC8gxuw6RIAVsFPxn8mpHFMvzgtDal4SSfb2IF
6FnIOW0nZ3FMumpe5Umd/r6hW5CnEKJrO4IixpERxp9bEftZal/CjMW9lPf/izfM
xFes982S4TsoygAM3bhz8iakTG6EKNZB1yf/ia3hDPLIs78+VITwjFTA/tCqELRh
9v5Ru4SzgnVQHAbUjR5wUIv31g3T9gCIqmJM7DJluIbrOEbAUzCqiIMaodzFmRMa
LSxB71rNH3uCIk9+nfarUOmC3Xj8tpjszPY3Tey/QqlGHcAc9+IIpjx6TlU7L6+j
CuKg923aGjweR1jT/mNEzfveV3fHQN3CaLkqcsWaVFn5C8RZ8eT9dUwVshMJvIx2
RcEPtAf6VG0FUSHK1ASYC9SCixvZtM609vGkNBkHBAqYe1FQ5gGRc5rLKP9NX6Yr
J4yDjEzrBJANn9yPlUAXVo66yhA0FdDNkso3L8zOiECHlmiqD7n7lKo6rn4Lr6Bn
aR0h6V2coWxU4O3sF9sZ+2ShepUCgNy+RdVMGC/iBjPI7jaYEyBRaSSn9xX/Twsm
JueoEHFgSfqdcQeui94pYqgfEoux39m7Z4l3DT83uALL/9DzVz9kHvpC5mY+yeGT
CulmG0Jx+FtWBka3/O357cnS1qudZnN1Ro3YXgSUmeNggKAhD31s8n/Ecg6PSeBd
Y+KQoDswc43NbVn7e9ezvJO9SoLjr5Z+LksQbkbn2RX9XopNqxm0+JQkgUeSRa8q
AFOZInd289ZQQ4w0FRZL86iwNoJPxIq36GWH5Ha7xvD7etKI+PJ8d8vFqX6O8ZuY
JVVMZz4KEy8Qgq2Ad0Y/0qswCD532pRNEx2RSkfXWN6yQYt65WJrfNQ26HoYVFb3
CBiPRUBUpIdtfZ9y3ev2ef9ofsckUHYUQzYaWt1Oq8f9MJSSHuSdH1LE8xcNBGYr
pF8ESgWesr3iUpF14Vx1YAn2zmM0dbXFYzgjsxRrfDF/aaUrh3cxArKmKLxx1sZw
6fgIcwU7dxhrzAqHwTAhcbuOHt/7Gf3ARaKYV0biMpu9DOEIjooC3jSY1YKuAG+g
zRNfzMeefrXn82MCKi6SyqOXkGh9xKJ7yYP13QcXPfjiXX/hk6RDd50Eo2DNFFJZ
V9a3EWmiAHtW/ybnTCkdTdfY0nucj1g0eNYRo6SZxTcurS0IA5cqBAyuaBQNBhir
PTa7ZRHxKaBzeOURL3bjFJTEQHzZu1YjrhagTM+x5JGSQaU6Yp7JMHMf/Cg2wwkc
L9My5Fqd0G28r+GP5rLft16K4ziI1qNFVLAPWRL8MB1xtoOAjAii3NFW1Agca/v4
ykit0wsn6Civ2v9kOTUBrbwurft32BYY5lnBKrhIfHlhreCF+kstA84bterDc7yv
fU1QxdB58U3Z+yGuz+7dvWOKg7u9sUzkB2XTHcQcTaIrQXN4qawnL1tRHJsZPHdT
VJv43fql1dqhsn+0NX82l042GgS2qCCkr+3OKjW3dgv5kE9C65V815a3YWiwsBVa
Xs32EdaTcRcZ5kzdQeQcMmpuBWwKLeFu2WO5pucXEVFYXSqKIYxjIcij8jonib+I
R1wnvzZaTujdzm4djPqj9XB4GN06BM2dGxyJwHdj6ma9ZfEJ3HYrw3tkXQwACefr
XvO3qwOeJUYfqTuOjwUVIOlCQeINgbW3Vb6+1qzRBmFtOPKLz3CRwnfnYkxy/X3n
JRvmeF+HO5DWQQmYVP5nTj9H6fKAh09VzN85PZBpiOhBY27tnaUkN2065OKqQFzN
wHRdzGMS9wQ/yV9+HbCBW1IIwjy39DXl7tuQ09mmSHpzWIPfdPDY2N7x7wOo6EOk
ZDd1snY5XTvyUp17nromoQqExaHRHKvnkJl/sdnBuCn7djqYdNKXvc7jO86TKQVL
Yyxk3heYJ1TZzEEOH0/gHxQIMMi4QsdolM6UsQZIvOYOZ/uGvn0FKNri9Dss5R+N
A8YkQmmbA5/5KAkpjE9F1XFQQWlNQkfs3l2luSLOJtihtt0a0khFPiXgDqTYkTVm
qnccAuOkLepqOIj9v/JTuKXZOSoSi0lGMdjBPl7Eyk4au9eXmAhQbjFelwroUvPO
6G61M4JpnqP/xODOaoEidw7jorBwgAPZhF1XZb3rZlMOwh8Z7QrfLUhoojDk7q8d
/OHBZsczE5fjvgpi9GOZ+UZrc9Ozgtc10iUrUxqioDcbVmDGcoI2981actMaw6f2
SYkjqjTwS8jzNMovAqn4m+QEDkA9g1atophR6FZwHOrqkBzcyw0IT36PkhIpH4/t
RZG+nJfYVTY38cKnOvesQTcBRX/M1ddygLTuJHF9w+DKOIBZXrt9U3mZQPHNv1Qm
z5OJSvz4NL1i1BiNmBFYdaXjsqBwgaBTs0JRucf5JnlJKmFc9CvXXhuMISXYOtmP
1Nm0qg2yBEveelxafcbCEzV5QCH2sNDqXC0Y0/hOsIqZYne9Ml8Q/IXlXDQWd3v8
YKZwOCdKo5QpIl9wVedX12yz9ELXxJCG+9CTFDW7odGf7aXCZ8nWsMbfAK/EcCoB
JhQymyT9peJCnOQ44SW+p5GFU3hB4yw1rfLLwZfs2Zj2vYI4UV0WWWjmTpQydnao
V4qA9y101t7dEcuOtWUqF6cT9/9WTBCaDc3AhzrE+PAxcB6K/+gqxBP5ET4CbHWC
apTr786pGO9bVkBDE+AfqBiNFIFy165nt2J5OeFS45PmjLgSZO3a7x9/HsiYGo1a
My1YS4Qxdh0IWJ5RvudIiCS/1gJw0/edR0FYYD/ApbsfVhhsPLiF76eUIU7Bpt4d
dDxaCgIAZ8wllb62pGYe6L2bgvgeT1RXW0i3pXwOIWUgoUfGmJlsBYwkCtCBKAtF
/97Cz6wGii4T5WDxS9/i7BjyhJP9p8wfCr1Quj7Ui0VZX/FsbFnzv38Xv7WNHYqV
A0SNICsWlnGzJ6zCEyQNBiwitd3uPtL6AOvw96+pMYuuT9voIwaBJ9VtxplgHmzn
smqaaFT118u8s596c3GQ/1brONpIG/Gjw6s6umlzdDf88l/1AdIc5Dyre5SAOjsl
Ny+dKEIsFljSGmoY+sO7aSV8qRTfCU5r9Ne+9Hzk9TtVyNbSSHS0hc9uc/Iig7Kd
x20e16442j+IF2+rtW6igA4qaHKZVFezTylw40H5zdmVfilWpjg4pqluWihMzc+1
l0HtLayPTSKE8cLFZWh+PthUFLBjmjjMxXsUaik6dsApTOhyoVxpO2PVKZpXMOlT
58SXn4VZ2ke+tYZuO9/upyKA+jZpAc4Rl0+MhXexkfOx6HCm+Vw1FrrXJ7iBSS6x
7e3F0yg4Zhy/PzFm8ZO7vRMKYHFkH7OsO0HbBv4boRPcaBtWWio+a0OCoYX/s1WP
cF1NXxykV8kNCkhnGactHpz+mjefzfNr2sQcoiM311MFZc9oOlIaBV/gmRuvqDmW
7jLV/107g2m8Vzn9jllaJ/OF715+qYvE9pnIaEIHaxd38SxWgKMPYlgdH5dwY3tk
qZjTmVVbwXLXNhry1KXgp0h5ZGU1RA5v0UuaYBGzVTcrFx67VY/a6UHmSELOlY8J
ArVpy8riUDkyvscOFqSno/wHFxSTI5ORTQVQRA0w2Eq70aTa6NY45fTqCAmE62cT
7gQvOKz3ar+UyKrqa2nWUYvyciJSex0e+7H4GiZPbvjrCCHgvXagb8L6XEuyEHfX
KnvQnqL8ikCgMdqaeTrutu35HYfxPKOUPpI/sZcK36njVxjx77ikz2i5KIVZlUFJ
Z/hgGJIOL47oiaLtY+JI5I4VxjVU7D8iOlPxROK+VSqxdaxYXxLM7j3zUj5TjNmE
7NvZyvmsTnNrmJu3eefF7BlmsHjcruZZOMjNh9jC9ZESEjf98eNAk1bOrcbcljak
nQ0Tie75aRYoUpXPbxbEM8KAo9gcXcFZ1E02YdeOuHYVYVJf+rmvPjgUiXM2KGMS
Z4i0XikOBN5YBhE5Zu5Wter8h7AQTEr0BZr7JWRxv5jnDI8FkU0hXzVY9c/CZERK
1PXWondODqTKNZiy0zh3bQgvHgEGYKqD1D5o35T8eIQh48MvVG1vGrR8Zp1KtHr5
PrxS1fM/6za/d8txyqeRsv1S4fCIOOspNH9kKBr2KTXmTG91pxNM5TJEk8JK5DUx
F5edyktQI8C7GDwCM7I5oT7TFlTjrUzy3QrQ/198WAdmXfkY1uA52IpyI94RrKgv
6e+ebGt4+s+NSYwxDSFZox4I8k6JxHfhVYgEOBolOuY/MqK8VpfF1FRpeG1Ytko9
EygRrvwEOa+bvxFNnI1B+4cm4vRqWt/CR5QUUWo333UKM6mzOhsx0fM5XlxHlRT4
HsuOKlneeymJkh3rLT/qxORZrK0WdfX0PksazI6MhwbqRVAEz+i/s+K6sb3hH30S
JJ6+NjQlBSpjF2oyl7Y2uSD1dZHZ4jdN01ZUPP6EN16zs1MZ7AFV9/BubGW+mB99
diZ/LNJ2uK5OftAcVKzYu2K4UOeJLPiCPPNYnL6MxvBhoKwwcdU3LA7UGxon3cbi
L8I5CG0rkn1SMrBBVmpi2LAKlurrX9CcyPBvZwR+sHLRotTs8YEam9/VTyMXmtsA
kPKsGtzbH2ri7M/D9vLUpGpt5uj+OS1Li1FgOSdEPjh64y7Lfb0m6S8eC+Pj03un
fT9qvWUy4MFBNsH/BW7VBwej6hpK8GvCOwHkyakH84E1oah5a3id9oxUA8+FBG+t
EB0zKUHcBjEM+VJ7LuL07DwGOdL05wJHgba4ooR3riB6mD9L2kRzJesNqz528DXi
dKhVp1oETRp4liNrCsKbAPvH5j40VRM9NQC4WfktzoOvOttyfIDFrWnZsPITMzBz
Xa3F79vUrFhkwejufvpH/J1kDRLhnid7obDM91oAW2Nvqzm/9zJ5aLNeISaycKGr
7aqUGf0ssbRBEsQ1n1d8pji4+yUmInbq2vve2m51eAr22Rh6qNkZGwt3L6PLdh6x
IZYzsooYRMeXNkgw+ztcJtMe4UvuRAQO6AHj42da7/V2P6tLVKbAW8Aw+QJ7ions
RBZxJoQMwyonQCOJ1WrC23hmxZuIaI1fQKAtaCUp89Qk1cNve3ScIcDIn0imNBr0
6HQai5PRdo24YMJLryBc/8FQpvyQy7gMlnWfr37dtAoA3JuSGptTOJ2BrI2qTvu3
la4XbRHI9rxCguR/0Hp3U7UBgGT16ECJkKiwktbla4QwUnUpcuE/tK0CPBKMLm9O
z96XkGL/YAhNdHesfrM9+QfzL90WtO72yY8HSNku9jX9QrHFKj02SokcSivPiXjY
0hqYEkAL5Tb329dVD4GSoS/LqZUwQ4r8oggUYmd1oxX7lrmcV7UJQkdHjUUqjiqt
Wljm8KEYchhbD2fRwbM5xo+y3LX9/sgw6rxNxCB9toR3JIH7Mps7dw4QkrnHRraS
LkoCdSwqxEqtgQfglgcSSafdK7TYM8/LX0QhespPK/Jpzm6QpBGS/By8JB3R4PCz
m5qQvohge2iJxrF3X1DoPn6r+Drw5Afn83i8r3r4hgdR1W4pI2+Vs4r4kkPgAkm0
Br8WSvzuvE6SM+CX1fCfB634C3z+5gWcSwZ9z+TcqlyRRSa+udzG7FWh6uV+9wpi
+ysJd+fzIE0RSZ11uTs28hbf8V3Rc9252D602EAFzIuGWj2jh0ODSK7P0Y23ypno
XiXz30NxvT8kGF8U8l5Xlvy+IWgjrg4ea2OkPD+e25y8rQV9EdMoRmquYwMWGPdW
OCXv6F7hkXexoAwJX3Sqnv2zTRq+f0PuSatqz/gDW8vpXsxXcll5EwKEx7LR2/XT
GGyCNnLOqVlKNuRVPAY0PQ8Ro2Y361fbd1yBCKboBgBCc/hCcTjd05Q8JJXeHq17
1Q0+CY6f+r9lO1k+DvHNRDxHJvRIdhqnImzNgsc4Xs3x+68XZqK7PDbF6m7hGGpZ
bkWShOkLKYoT97tqJsP7YXhL1dowdcLF2mg2wfX9AWQAnMwcu+rptADAbgMl1eSJ
BJLVPcHofNlTya4oPlCKb0hYDBa8pN1kFQ+raIdvXH1o8OKY6WHcs0B62sHyrle4
bRBHUw1gHHkokbbJ7lPm0xRRDXcmG4obZ/UxdWsSBUYXe1VVa73to0U+3ATo9Ztn
xne4/hxVqe0bZ4Oe4KEjt7LLx5958qPytedV5HaGiGejkWNrYS9UL/vzfNULQrVH
WioCvr3f2k8g7hbyntj0/5UcJm4M1fvUrOkbr1ZyztL0QPR1Z3Al2MRNb5grmOf0
TgPvLG9mOfQ/2Biu2FFL2xemlUyIl408MF8fkEQjwwc6UnsK1bNZ11yp3e1VuPZq
aiKls/fuPBOzO2F0KIeXTU/BtELRqS+5FiWMJn2ha/lkTnXhR+JAE6mcwcT52jOp
Fgc++1dkKPK6vECX4X5vilD76pVMVUW5/tLSvn2XTLR57hj/ycYsqKSWJNOF9PnR
W93aW6T+VmK0sC6WcXx8HOi9Px54Sojin2sc/ln6gSAx7n9AG+yzMEAAYrWxDxZG
4gT+EuffZdAN7GAlQKgfa1hwlKLmanJz+yUEGYgVbY9z/ou713IbZ3BorzK4BDMo
O6bPEQ+VyXqIT+nOYC69q2dtmDhIUQH/119AmaI55qWov+4+zZGErAyTdvmv7d9l
8+zYpHNS9wUg77RaDGVh61JW1dWyqIDyWXfFqrDQuHZ+m8QBqI/BtbiyNEeR2KRV
IpCsC4aVtX32sPndM9ERjMO1nf1vASrEHUy2jIxVsNMq17DdWYuPQzlmLn3CUKkf
H9unDMeExiq7ftowMG9QAv4wW6BRzVKELvKT8nF5pUYDUmH+0lN8ABGmwjipbWLd
n5lrrbAYE7CI613OsrQp546XRD/wYTibl+YpZRBeTdsH4iHv3o6CHeWVMyHI9B/s
I+HjvJtbay7SF+26cJplHUMscc729EX9ezpH3V7oTloJ5Wx+lR08m1CDY3XNpR/0
mg5rZZyDPMR/DzI5FNmFkNCz/jBLvNys8oHR+PpGB+jdr2C25rriA8Y02aUnR/tl
Hoc47znmuPVl6DaouLOcPT7Hdouid5pgi29C6H3+0Rcg6/xnlH7IscXFTLhOk6gt
5Aed8YrW5+XSLjXZH1TlrWj+c0eLWWvZyM7WufmmYOpSN+Yi6LxQks2zJAygNoim
HegFY6Asij6VqYnsfZU4VcnMRml8jyUrrLPxS9IoGROFF4S0RCxGv0s43lsIf/7+
ebbTqSigLTGDHMPRY47QKlBL44Kg9giU2HVwvHczV5CDuKGNMq687RMowk5hCc5r
OdiwXCd4vvAMx4vO36K5RMICeJrcOflhwia8fog7lmUbX/RdJpMUb938mHSJODLi
d1W4cCC1kKPVNutWr1lexGAJ7hzX7enG4Rgsow0Jnp+UKDorbHpTKT27Hz9Nam6q
8BmoqqY/nKUVjKMgcICSnfj/MFM/9uqrnHSMkwIBkfU7wbojRUBXDtp0aj+8hdQY
g0ze47B4Q36t96ninH1x84e0z+Dki/Jk7s/xgcbQ0LyhVRsONYXyEe+jOkNbRke/
uhfe8nULc9hwADpPfDlOdTZyCreRk1MS8PycpUUEiLNPgAZA4249QZq6GisWiN/2
HR6RSFNNPUsg8k6OtmJ9Bnv7qI12HR8vO0og8bdZC3FmPMNOy3hEbn13HR+keKgl
5LZq3Xiug58s3rrRaHft97+W3zNod1b27KPQP1PktfqD8LScX8J+Sp2tW6Ly+7aD
bPTrhjvrLuuFM9RJHXTMiX+cHtyPY+2JO2S6GZQrNcCBTUaX2vWwmb5UfSOySoea
1SLUMyf+CbdCUio44Sg5Ig+yXKW9dU2R3B6vig5FM4w2Gvg55VvMs2yjPx/qXSld
vwV0wCNECcrt9bJloS4PCcreeAlvKb7O4sA0GWMUnqsSwfyobJoaqoNuH8CraLd9
aHdGNuYP6ingaHoMj3UimWSYgd3zXsw9AGWvrT7n2EIfs4p7C54llPZtyO3/gg+q
9oTp3fbIHpKFMqJ82QlQAHHNd1mUVlWgkyCczJHhl6fZxOM0IywjdAreENKqxtH1
1LxYQhckaZHjuG4EODVigddstfgPMacs+6zwTOEkQ+Jr6MR2opEezVS5eSk1DXdm
51IbAa/dgJa9zVNR5QbNm0XEBUsz9lknH+bD/ej+Ghz7LemmtTw86qfK4S/AJ0Xd
6mQnexX1a/SLK7ZLzaecwQ92BGapOFgFZJFxdUszjlqcJ4Xm+3Nmk/Vi7NaInHmZ
wrF0CCuSctnOKrObNIZGay+fTPoRzUMxz3dLodPr69BFPxwX7Lq7AmszfVj+K8dq
EiKu4spdA/N0nqCc00RfBn5DJ4HMv/Qfa1NSlc0+UCgiwDExKcuO06zKvp+nYmW3
n+PD6qPF63X3fdFzBZFsb+ivrovs4L4GCj/UkHyULV/CTRRjHd22Ao9kdwhdhfxq
e1pZCDtd3Qr2u66Qd3zBGzHWRDiL+JugVwDq+vf/+SuNF3Jh7uNlCikp3x0/CVSW
uF0vb45F80ND9tPccqdPSkaa0fzXpcXT5jVKliLaeUjgkVe2BuV99e0HRpzLr7sI
x1csfan6csn7FPHL4V6OoKNd9n7c8cyNwhZ4KKb8yk0qiMOn/BO1Yo05UV/jP1Qi
Ze0PSGZ4Wp5/TCqszE8QNC5R1zqffto2hn6FVwDMfQT+sMilAsoMwo/v+/so7ebz
DQItoKdZB/9ZZtQlCo5RzPLkmL43f76EFVJSO4AEG494Zip7SGyM4ktj1o5RHb7I
QyTpRxWUVqL/t2Nx9GjeQtqZ8yXFrusHhVlDs7FHgUnnFbV8nzbaJosgwV0xYmbJ
vzN+A4EAejQ9DUl+3Kf+7qW0Z3umH3RdCGihRJi3+QduekwtF2zGCpnezr06m+Xs
l1J3ZE19eG33fpN/Lvads2jr+9ep3WfhaxUNPb9r7WNfcoX26V4XJfuiqS9UXp6z
Pdwc+tOySUlv+4HmCAIlLXuG8l2I98ZJDK4It2jctVrLgnVMEQXkgyJFLCVTeV1G
AaiFfphOa9MwOrY+Gyvrizl2Rn2nB5tFM9tVBKK36IMbf9wln80R1q4pQVb/jAh9
BBKi9YOPLXpykoSglDberJR6ievcG21C5x92pACU4NickEL1g4qOi/WbFBkWlEOc
k03ljvEDfHsxnO5DvZz48KZQlHUW8U5f7Rj1SPWMYoPsLFi1s2g6Ef0kVKvkX3Ft
YbFjjVJKQnxyA1XbFjWMnoN2JaqXoRMmgy6j6Uor+UswAtObIPLgIQo2+ZSKrkJ/
4TbECqn8901Mj0YkR3lU3L/NcFMEa0ocbp6r2dRaBHXGJEzstLtDv0d+i7ZXQx06
/YayBdVeR1pphaq4XjLEzzO8sypiw5KHfAEG/xwrdJ6mOx0s7BhH1bswqAPR/JHM
pgr0qvfgPpvdehQaG/yjMBCZ/+O0iCBsVhQf9mAKV2mPsp2EWdeNnC4K0Ekl4brC
hg+0DZx3Dnqt60VbTAG+Kq++ZEJAMs0QWhn7OLNHFkXLsw2lrFldHQS6jdI/+OYv
oIqWQt1U1sh3Sj3NcvnXabRq76aYep+ftlRuvU90RCu4YnhURhNbs+ZGhoWd1AQH
yZy0/UhMTOVP/RqcPO9uzQb6BKjrJAIkBzd0D4zgMsl2QsVZITBtiFqwvPBweiii
YW0+iw9oqFX6gHXeW4uUtlBNsUxJMwHT5TPtz1VAGzqno7rE+34iPl9+5LeQkPxt
dWhBbrT4D7C+Eh88Aod0dOv94bKPflEqiRA4VK7Gut3l1nRiPasfmK7HLJ/WR8P/
36FboBbW1q6Bf3k4cNNnHT9//5uL5FgULTXdgHdpLKwna1fhy77C3nSk7lWSH1DO
qUlX9QRfU1P8aPiJlKZ8lvk5CJw7ALjTjLlz2P1WXUTRlnNosjiUdqcruf5ck+oL
twcIkPIPP9LCI6sbC9dBz2g3Qs465z3u9jXT6Bn7AUMcDRlDi4wliCaWiZc4JFts
S+vN8nsGev/qvQ9DrAvG6iQf2ekZGWwF5Dn+BxQj8+bMjW7oYKWlV7lT0J8OcNIZ
smAuMKRDjK3g6T52Hw1j/ckG8PL194IdjFgIRKLYaWXfl/kRdLRBNTNUwm6Q6nIF
ueLdKs/6/tJb8mLMi7bLrqlvejfQNnHvPJRE57Yp2Pm435276zH2S5Y9st2HFvgJ
dvycITBl5pM/LP/Sy38CFGkNT3EBgYmiTsuU/MVB1VZ2I/rpoRp3anjUQM/t7jb5
9bkaeANm4Jl03DobtusfRiGMABd+94DFoZUEf2N9jWr2Ffb0cL09QpgSLqoJwOFv
s7Cjty5fWTvPeqAkMo+JPoh3+Bt8TAJTad3Sjl6d4/EcKAatwuEUVJXT+qM3t35b
R3Fzivcw6Wy2EubiahDrnfr/S5WTY/8ekZYreepgEwsrC/+Dc63HezcMMy0xUfkp
zJAed1i+gftZkD0V2B1ID2qrTXfl5JIa+BeJfJ9sXdIhOHDD7IMj2eTs1f8iCoMX
FfCgdYRT1vVWpyfMTwtSuj8T1wi04OM3nOFCknwArl/tcXZ2x/rZT6w4wowrrB3V
rb012dU3MMyR5sjlaXEGNTlRVb7T0XRNBndP85z2DV85iIT9iUu1t5IwEk/caiK6
1GPU585LFrdky2VmgWCjtExFaWcFjVjI93mtsDH9EjZAJpA1oVvNSEp/qrwnXbXo
rp+M18EFefDSWQligWKvQBmFiQibWEAv0tEaRJXDN38JWDaK/2lVYJlDHpqKMkWr
xXZmhSMdMDP9Onlox95zaSjdiXwLKfA+QwuONqIq41zf9N7V3fyiQ8bRL4wAPMBY
pgp0bdz8LAB+E7P9kpsGDS0h4kGkxaKWec0LNsv8YD8ucSlOvq4kUbpVyDhcKBs4
CiGbhHGwvGeCVQl7q21JYpxBkwjN3ZbrE/7row3oXy7WhIu89/CJmKUQfRQ/9HmD
ILqc69mTX7RdG7MefPt9rcxG0otsSHVggU4JV7NZANIBBUWsDbJVHd8t+nVygMQ4
1a/qyUbwRUEdaCj6fJEQSoGgiapHIj+HgMwtvPejSZ4o0sbeiJIkG30THpO8OGS4
NT0duYteor8NY++TPDJZmPyk2CzsncUWy7gaxi/Jb0df2zyXyWe/m+kRhO9FWLzn
EcDUzSZmnYuWE3SMUz0W5UYSEto0vMD/cOsipPA9/sLM8hAJ2P+joxfZ9wRWoDd4
vDvrkffg64dqjyMhKYDCn5Yvr2gHAA2LICmxwNe18neFGhAOP/por1G2KgheJ5ZW
1LIqsfV5nx3/7AkdBbOdE7ehdNR3SIbs6/VNMYVUMyHG28YBVbLD7PpI2MMKdG8m
nw7EO7oI/ztUdjo3F9nyP7gd4Z9DQNpBnDNSTb/kn6NYPcX+z5nAlM/bmKk8ayq1
RbTalcMUq3tdB1x7nDilutLcbzWQE7SWnARRB0NMeeLQFzRjPp3Kr7o44OyTjC4p
mHrI+p4tjH0lUAVEgxH+0bZmKpW0ayKKlNfPPDEBwYj/atWr67elmepH2zebMOOb
apg8RKYE/R495VEasdzBcL3aPio30R7r4qqjuReenNEeGReuCmzDGmb0fR6cLD7c
HHGcIbKDBVLpPpm2YvtQfk/ZvTwB3rbQ7jf5AANR2lCtOibGDE4yYO+ql4zZEvBJ
LRF/hNbVNDR/iBEbCvN5HQE88vom3mZcezgkZ5qXHp4U7dflIoqtixqusQtCnxOi
vDySyg1027/yIxttNUEAD6i+nbleJj46LwZ6iTHpaps/hKNXboYmRmdROqJL0gJw
n6fDZKnpym3SjPuoTP0GclGJxe99usQm2IZyDzYSUiH7vMhCcw7lQ1rhSeMxznjD
7KNO6TGXaM+KtHr/MenGBrb3UksV/cE04PGaf99kBOGBuR2U7WfyfqSBVkd0Ly77
pWtJhWpVa9fXj4YWka3Am10f3OkBsFJL8/mLuQLN8gO19RSRJlUQwFSKJAR5TxN8
z4ffJcHIyj+lkQBMSy8i8TVBv7vFK0L8Ya4zzWs+vCR+cggKcn8FK2pNbKtduPtc
PS6vs1Y77fJmM20eQB0zoxnz7bJnuNovz/qQkVKRwg/Ox1HSqNIyhRjqmNAA/O1+
Dr18wZkTBKiLFbw3huxNAhc8E11ESIdBxz8Y8Ff1mk/GAbo17xXZnneYafZUcIcM
5SvC+Sv6ZEoN9xLVtOknZed0faJbtuXLpYc8xzKI5TbEZgb5BMA0XhxvfKqBKeLI
IdpJgszmqnlQMTm0q2BiXeAJrLLCqspEwxn3xm96I+J+qmX/tcnOY1EyOkg16lXY
P+GhKxY+83165dGeCEWW+y0G2nsqnfyPE9m/id2rHIMSMiyN/YL6LOYha0J7v4MW
CeehLdqdU21J6y9kN/mcgjA37rxG7KMvGr/JvC24Go3jRx2c1ZhDy66mDYasZ/9Z
S2C25uezSa09lKcfZ0sO0AGUUMv2UV5SXtry3AWabgD3na5PjCE7Vzhka2TTMtj1
G0e1gVg34Pi6nwMfQLQXtPZ3d41waOxYJM1oTnrLEok0ScNV1VneMEPq+rAHI0IW
MGnKOoSf2jsgrORq+sRREVoANGPMompgucmm+yQb89sYr+yPcThiwfEAZV65eGj5
/XdZIn3RbFJ+XMate3q/shokka4nG/AAi+WnDmLnqUhtpNGpCs4l9ILzoNBdSaZf
+WLnyLooUbTx/Fw0O9gdY9JsuBd66B1wlhCXwpFsaHqt6vQMAgq5WizQcrbledsV
b1Wzg6hOMw0SXEgC2vhIW80196+roQTvZ9lws1q0LUZT7SHDkoy31Xv7r/y3rPrn
WPltTPAc0v1lRsogAbR2Je28XvxA3c3QxYlvCZiHoxcsSH0M8SYBqnYic6nedAX+
Tpo1Pld1gOEkq5OPqhvFiXmyBIHpYnvUaiQcNq267Yt6HtOIxI0e6/0JJpIcEwFn
4uj7Bunr0SRM+Oza0umiDhgyz7bEnPXuOuonNHhocMX3hYRHih5I49DqSaTjLB8Z
NOjK8czj8VzhtnfZjHF6VtEBDlz9/l2Ii7RdOoLVyuhcroQtAt+r+8MDJw5FxKOR
ibrRpBV7u130cRTS+d3N7T7AhjgtH9+WCYlZytNLsp+1ODC+dUgfV6zGtGTDL/Sh
ngERy3LehHl6UmZ2aCbBQG8fvjtVoCQvpc8tJ2F2lU8h/MMOVhGi7Go2TMTCP4X2
lJZSIDwHKvmk2yQbo6mhWchVsih8BxkvSi0CLDw10TgIhunmj+UYfSc2MmKziqVe
GnFCjjfWeqdXQQCz0YAdI58XCwb+TP1j92kOZF8Jd/X2HE+dDQMdMLKs++8L/Y90
HEAYGJBESDYDZurny7ut0sg/fFtkSaWyS3Gk7sZ6kv7Xc6nXWol9Z+J98AhwVW/Z
xjwFVdaPJvvaUfVC81OLBw0Q+mdnbi2BMzocQsSiOJ+GWTjZmDFH9RJ/DuH7PmQn
HdElsJyBttxrBxCT7zUIepmTey2yB6/nzvBmusojyCptjtXzTM7WhjyxgZRBHo/N
OMSog5ij4yUDq+KKaDESkH6RkXMUO1Su4wpQQfUPZn57fpLlBz+ZXMFBwZLEYxC0
tWmNNMHfnRiAx5FAgKsa87OmEuGwwWzL7On2yEwt+PdNBm1zv4A0grh+rgohoufZ
B1olvQfrXYcrLo1pwQq2wCZgMYaXXVY6U6e8Yhsw/hwZCj+sUQf1aGa4EiTGjZ/v
4bl8J3veykTnChZjiicyiHZFt+gIuV7dX2nt6nNjyQyf2J51zRN68/kRtZbemt+O
CJFtWgrHbd6UfByxiSEUdM9378KNxW/KkInqfFGVO+welsn6AH4nYbKpzIXH9fW8
dRIg1hanh76mSkwuY2bUrKX/0M79+SHef8Ukz/GC4t+lC5CRI++3uUFBM054oEHt
Q4nJCle2t8z1pMV4BtKuSMjgLvaCSiOaECA5BVVeBPcf/z8tYu8ABNK3kOOgCF/6
jFSpU8LHU1zcDXZJHvvbLI+zzo1Kqz4cxPMnRlHQ2jd8EUS38ottgrA1aXmEEHw9
3W8lhxDbYL/zYfveVMzVMKbgY+mWMPtEtdt9p1H38LguoB4dxd8PHVfssYdQmnH6
2q7MGlDmXNh5SAhZccTn6muQVdIzhh68rv3sIxn7TKAgYdrC1ScacXR8ISF3IVIA
OP5izV7TLOr82MK39kCNrVJbS6bCJYWKF612DhIwCkoTwt6q2zqXDeB8SWnFcHRY
eRWyuHROA1X+WtAdHCAaHd11fRtpl8/Bjcgc2sPnw1sM66O+NTd4T9gl89/zqRQ0
Fcgw2BnRHfp+F/Siy62CgkLyXGHPXnJwds8yTGeSLGH7ggbhfj6TJuUc/BczsXCI
5A20xQHx+aZ1qAYP7o1rLtfKTfZxTbpirHW8+mfPkB6qFHl/XcF4crivQk2mdJUd
lOGoUK932Vqbi3gG7o8GxrlM77pJ4Sbl+DMiqV619Oi459srtXv/vM6dbfnrcG1e
JXV0X7Q5F7OF/6jXzA/1lyrUJ3f5jOd+Xpy2cluMZtWGBv/mfPkrBZLyh7Iq8UhC
wiULh63WwrsrpeXojm86fgfpR8xvGJIz8ObX0B6zXDsM2EFhn2nv0rSq6nOA7PPy
BATAJiTUD2B/zXtXlZvcrjodB9hzJ7IGd8Il4GYtwv0ptzsRZtKHg8n7x8vAA3Ux
mi5kXRAIQB4XubSAU0VgKtZkid7VAkF4YHQnMwm+ZBM3S2hnvqmIZRO2qKld8Qer
xAtR00kfaYai+6fEa/NubSUIBvC3/gFmRyjkKH7ka53+lG98KqU6sf54MwLeeIhX
yr/c3o+3Z2oY2wWtE7W8WRoZ23ywUeiraYxzNouXjK2ziLRGjshmn5wALnod1iOx
BWvSWuTLYcWKqIoJembaOhoXtQiHPdOpqt3zZSpCti/JVKcrY0QErP456eyGpK+m
ElmRTA6ixl5pIz2H4mM/UxtmFyTiyeSEMk0MebDbkmwkaX2O9OU6z8n94LAf8VnX
a3lo85pQa6n0I544PkNhCJAhDjTUkoNGaRJ8jmeXWkrKQLPikNjCqeu60DZiouM/
XnsVuyu4XvOlmBH802jR95qMdz0TTEfB4Oqiloa68bEj5F7TFPiwnqF3a2h+gHLd
NxkiPeY+JtICB1DGoTv5nr3C0n8a3wDT1yj4Y1RC6QZ8JBWJo8Y4BhbizjEiWY1s
QB3kBRcv1mDYDm04mwQe58CvYCu+g9ro4ZzVU0Lh7SgMViYi7u+n/vfihm6aGaSr
lqObtqsax3EuvIvpInpYNr8J1WWH253Oa58ev61SOan6vt2nFsPcmpsulBenbfYn
sodZoBi7r9zV94ywBqa+jrpaJsBg6818hJE7KO54DAdffSGcG26s9xgDSeR6D/95
5wVgOlWw1qfEFDeUWbo4Oqod7iDtzsHy+WBeQGuyQhUCdAfhcmw0CUPSoobQHADd
2ScZ0ZNs1vZmo+KJWgPRNnUlTENcH0Udfjl4quH7tnWc59NL8fSG9M4zjqrtuO1X
RH3VH2PLt25ObfZP7S2oHZID+Ophif5DwES4hMFLfeCnClZvKl2Idfv9EQ6sWLMX
wkJDbD1n0Nd+juo+ee5w6BKGD4D/Ntgeva+vlgZc0v6o/0IDetKIlnAN60YbWYd1
AWzuu6X54JhO4tU0YoMozpMA/0bWdy5YAurhiSFxSqN3YJZKmUye5m5a9NZ3NQ/E
M1mX1TrrP3r68bwH1xL68dS6wYzFZMvkuQaF61b9f5lD5E3JKTOteHuZ6WcfhBB2
CzvKL+h1RK4ypjvAGJlkwCHWDd4kD+CT2E7tS8/eTeh3rGsAHksJNh4Qzfly/9wc
C0c3zzsr4Al99B3BoipYr0hvXjOe0qSQ0jfX6XQzn3oNz+cG+YUzI2EQDIkMGv6Z
MeiFcXflTNJ0/ONfeNt4qdrUFkOneDne31dbCCD6w5ei4ENix+DH4g72Yi507GjP
YblQkJlI6Qky0e7m8yz3dasKnvdpcStsw9Dr7SQCOftuSD4pN3krG3VV6SjPvKsR
0dTeKFcWGxmSd1ZW8k/vmXAdYr2ll46ytTnpgzTJcFdRhT3ja96h1nwn6EGGwJuL
sHbuA7lGzTzHOvBqqZd4FMHgIbgkUz9b24a/aX8U81bxGcQ3hvnc6gxaeTjIuzIR
/j2Uqk1SQaW9s0YqreY4Sw7xZz0q0pwOZ+uOVpe768fp80FLQJYdN8r83Ug1/jSg
7xigfwg/gTrGB4lBogOXQpRCQiqgpYUHnDMUShEV2SatxDO0kgAils4qYNtK1C6V
hnIrIZsAfT9JS99qhvWUlxura1CI6uQwDgdX4m1B5q4U7eG/HHn+OZxMqAViuKX+
c343h5sfwzY3IAVx4T8a/sfQtD9c3vIdbjIPLkLGlSwad84FK4XkgJzqR20g72eh
d+TrP/rIqvdBzc89GEDxactDL2OwYMqcjvuYY8qSvzNKUVefr20gdmIte9HIord0
OYCKAYaKigDw9bJw7SjrlX+eRcjNKCyH4I0YKRnkmpRuOwW0iurq7imj4FhFsOqb
WPQKXE1J+Z5muL4OEXPyZLO3NA8TpqCFetIDXQskW5TH5GjOm0Wb9NeNh1ojyz0L
C1zwt5hOxVe3yq5j16wnxKvLGuw2Thv0MXxRESmc0jgbCEz5xjkb+3QVBLJVADb+
K694hylfKIB4twG2RZaMpssCYuvtG4QOolId2uV4raLrryg/hf2TwOp1xVY5iagv
+dh6QqSOnz5URf7xZ5uDDuEnNoEFCiRm0MsfedqQTjXgVVhRpEIiEgR9O1yEYYtd
p/E7SZpEDSpCId/vRQlDyCrfpeUEdIv+J524T776H3CPSuVccSE8g/FuRa7O7SeK
wn+fKxrPdBX3Gkp581UIazV6YslTuguocVh/yT9/csaE1qey9I0+wytdq/qbOSPk
6m7ZNtU2FFqPbq58IZJ0//LKIICgCeXPAW0utUnagLV3lmecD4zYIOsThZ56OQ4+
Hhazu39gQ1zNt8t6MGbGlZopbEzeA9CVmQyljqHjzsDmNkks6b/QLsf3Zh9no2ea
wz2yxpnkFHyKbnf3kE2llO1ze9DoFc0MVu7bS6JMtbLopwufao6eV1ymXRhRjNWY
xntQPKeglmGzcw+OojSnAsXX5/RxU9kSgn90uLyxwLIEWuXQtL0S1Wdq6Cv1exOv
0JFLPcVMUmrR4jJmlZonNEQLDLnaXHewmLRKnRhBgY2uygtQgSkcbGJU9eb8r6xD
KMMqIraVeRgI7awPgizEYi/UvW/RlSGab/VWzRu3co7t06VRelBsHyWrK6ruUwMe
lRkK7tc/iHpelOYtUPvTZeG6A7FHSFfgbJM34dux1ooLqcEj7FQydzMoMdIrT3GK
50Yba41beqmNqBJtD7N4Qy9nLVedBkAr9SwjcNe4f7kTk2GYdXN7i0+jEQ+QkGY6
boIT1cWxYdgnOsei9ZF0WtwvwWI1hkZfwC9nY8MaobRTCq7iKN1MhIUTDZuT6m+o
PLYE+/Hy5K3Pr67d8OavxRledCCU9qeO/FRGXM3OEVfM6Pf8Sl6FXc8hO13vFAG4
7JkUCUwwg0Sm+YCelH1uBS2rxmCjjmG5Ilo7Qd3ws8RDKxnmLRUGY4Ut4Avbtlxi
+1urGnn4RhxvxpE8vo4PSNgp/uKLvLqkx9A5HgZ3WsRs9cU1gofe7gtTfVmFQcnq
WPxIJeOCm/4mqNZi6FIMD5EIVhSU9loXhPqk6LgFUrN64rByBSrbg9IfJRoUWdfz
KXl8KqydM7ok5dQ+GdPHR3uXVNWTzxjDND9WJnx3IPBlVJx/rBnk48lKt7/oVjBk
OtevpavEUb9Ay4YYjrY3mIKxwsZFYlY62h0NK61W1SGVaFJT8zUdaXqqcRjtiuij
td+gbQaBMH57L7ioSt3H3+lzHtDA/eD44koMJ2UaZmt0GYkgBXEFNkvG0OWs+6Qe
/qaUpUe5qD10vfnwhDSR+WfKL2hquNSW0OZ0EsMntxB3uOmC0t+1HE0wIzI45O7w
dpuUP0Zo7B0PngeZnT/Yfln6twq66IxQaRbUGSFeg90Gh4f8iveT/Lw4uIIaEZmO
NfAoHxT3ZG+jPndWDdop/na3Qc680nrbavDMiq35JnYKNj2Sw1bvR1iqpkP35HGe
+V3pXAR++6898v31pJnDkjOTbmOqB2dF0aAYZIXFj618MQMvBzN33Q9tdeipTq1v
nH54IUC67oXHadOs+h0egNMXuuXJGEBLgTcyMzMS/YVitPdDFI44btnplq9vpVZo
4QO4TYfjnPtjD/zODNxAvw1hvCvioMm9X3NzvNsYEhK2i0O5S/uGKrSpxMYKrPBs
vSNruNkoVXdGdNW/D6y09imKcok0yAOCSO9pF536rVmIPJbHNEr2vrskwHbxnbgv
LzuFJPLAPSkLc++lmwgpe6S3Mh1SVWtg8apiJtqbcLZN9WeObN6quuI+lzKzjmVa
YLxtBdH6T7dc+AtPwsfli73yNHbTtCj0GlxWzW0sYUstI87La6+1Wav9jv42stLB
prFAJ4UjX/aWWPxiWSyai5LPJpBve9GBS+hCoFx/tXxivhKDQBas1y/tt8cXu6DC
232qYBQjYmllQI215NB1KRJp5BedZVeF2WhSlaMNW+bciF1HB1Pht5dtgrsMqTSg
jAjXV8mbbKDlvlVbkQEMvu1o74Fd6suiJKpOiAFRI9C/cUZbNwOFCf0SxWbSuyFM
X2YBoeR/FTfajtzlViIZnUfGWciCLVvyf6jOcnreuCm9iruzU1UFrKf0N5gdRB/S
nGd4SWzox00bfb0Kc03WpMeLz7KBytoOvMzkOyJ35tFQTa61bHUhpEoNtgwOmx98
PLcrxde/cQhwspe70bGHM8lzJIOy1gt6ExuvnC5llNhkBxKu4ye7b3o+B+RK24RI
8bKkyNyrYmnWWkDmB8SoYS98bTPNzfMrVFoHbnOBe99lhb8NEO0zTQ4H/eSb2aTI
szEW/Uxq73UZ940qxJLE5FsceEr004sH/4d4GjTDANpDQNtvM1qhi67WbwTP6K8x
8AOAG4BX1nkl0I5nl18FdYAdp3+6xLOscxBneJFja7LYaB/mTmuInIkuW8+FdnoH
ka5eObRtu095KZp85PjU62TKIppMDGKAFpBxCw2MoiOAKQUFf7yB5l2fsUy2j4KA
fjhBgGYXHItXt6yIr6UBZ0ZovhXqH9J/lmtH6juG2Sqb3sPzDOrpIuOHL9zV3i8L
6nGRP90w9nijKJwwqRLROfT+uHWw9G5G0C5mOk3eMAzMj01BcI0RHQgzsRMLZu+t
CUh7VKdaHVVODp1ccwl/+qrQFsi95olDQW+Kjnehxv/lAOp5HWr9Mh2ey/oROD8Z
7kkz+9RosJ69q7ypdjvB3EiaWhgtPJt5Rx/S9hjNRhpJ8ZSYG/3TWqGn1KFDUJH0
I3c6S5XnGcw70InSIYXf3l8wrBl1G3A3Z6ua3Zv/Enf8ZIOqeeD4jdcu9GTrbbe7
I3xFtrgAApEHvncP40tr19XEh4H8P8iVJMNAhXUp/QY8L8+uHjlL/XlZ04o7SVri
nw3XS2mJAzHnu+CAuzZOdmn1SuePoQmm4fyT78kFf14ftJuKMBO1qYOrU63skHsw
0LE9JWaRRt8idCd5AwHq35j2EIL68w7YvD0p4PZI16BD6gzvApl+0ulih1Q6Zcgi
DKbV7rO6BwYj7Ep3HpU2vQ7pH2A1Xigb8pz13pP7aDXf3k9aYBuRg6NI+9Xm1bLc
YvK6unMmj6DV6CAuwp5CH2jyIzz54i49bh8Dc3WYt/6QIOVxPzf8eH3SY5ECB/5C
z4408ByjWL18HsBoN/y8uuJ2s/ROhoR+A+j2wcSiLc2aMYfgx8/jEhqUYKgoW350
dMnHIIQr/IGe7+5Jawu6qXz2OMIAr/LoKWvuhdF3X5+PUWcBf4PtesGYWn2Pqw/S
dP5+QSNtPLrBburijcc8xyTnYsCVOcSCUEbHTv0Eh2dOzEDAYLZMXzC+xvKUmnZe
ubFEXjNVQssUYPjHbRP6LzPbFwbYHToUi1LywsePaulQard13jR+YgwdwZ+QjiOR
ndyftKZTHbLT7uOXeMG9T247Xug6+z4O5Kl0x9uuSG+EVLcVC+PSNUX/Dz/GWlf/
IyJry755Vfof2k3xcOuWwOr1c1CssxyTmqZOFfGTPUKdKrp8UZkdsCAVGlmcxuXw
usf0dXgCUTN8JUKVzPlAwx92FRhfRcIGhujTK97QuluOGY4qkwtqtVjMXwjTbdxf
0DcpvUR9Oy7d7tQEJVMoz+KXf0CeWE7oN24C/MDnRMc6gkICrBA1PDMSx/D24V0a
hIOfpjerxG9rfUHZhZUeXfvc81TUNFKJNernMVOnRJzar3uokuM8in0PFu2jcchg
GPRfwS+zWoz/kN4cc0T0VQGyGzoh5xP4WCUnRgKYGEI83M7jKm3ygRG4JwkeOZ5m
ua9kmrDPqWQjaq0nQaQTfz23MhctD1YUltGaSR47DiPEQk9LXw90qZQF9nGyNxzX
aTWCmfYxy5TboRCCzEVQFcxdriSpzu7pk8RT6dcfycE6iv/VvJ9zBPxyMoiakL+8
LXbBqK51vXLYkHHHPHtqHBTVBO/as2EK/2HWITkTXcvVuHz3u/hquYl4ItXfxPkX
QUguqBzD8dMLIQp+loPlgOkvmAKg0mKtKRXhQAsM9g0BXQXTTltRJ4u6YZ9f3t9q
/K3PmjaNfC/pEHJ0clg2dMgjPK15UMOzZTKBG1oGeTJ7WQJnGcVY6QPSfPC/sI6p
1J0HMoLz+y7fbGidD5y2ECOs3fpWrTjawer5TnfWvpKZ3vpjSGpk+7faLEEZq9sg
nRjSh6meGRAT+rTGLuMgcNtWV4AKC0kKLy/Cz04GNnflRLFM9FSysv8ANS/sxFgL
u9CTwptfRvx5USUJKJPRw/23Cd0G7MqctumrJzDcYYNq5aX2G0fL0Xvd0Qp4eri4
4fIoqnvtnHAPbLml1CfUatS5IT6qd/S2LExa/YcQzLjXrqoqjdNmJMkSp01p0lv+
R2DZvB9J6r4WZA1ZOx8p+NbrgZ6L52GlYRi2LTRHo4+F7BaxLEl5dDT3Bmp3h8DT
+0qrVFc0jOL9sA/ZLzimDWQwpE8osrR0y9DFTACw3VRfr7H9U/LagPKqoSGZARWB
9QqmtYsMNJ3aSiu4r3jUsWZjscR9Bkp7fz/0e8z08oeUpwKWDA4zDFAz3vvNpisE
q934+qc1qct1WK7uAR3Z4QEATuGtPTfR3dcjt02uv+umlU1/afOTFYyN4gfV2Mng
BORgKNP93XrkSzw3lIMw1F2T+mWxcWDEUXVxJeSCyx9NOXdn2snjVZnJQUtrFB9x
ojU/J1zrjnBjEvChBQA2DGwtNZGf76MH1VAyflQbQmlJOI81h/V7JNRjOb3sGFRB
MPVoknaGZmVaDD635R2owjntPvoFMhHl6gxmNpcTY6gTOio3ceDEO/TKfKfFWWXE
TSIIcS0JT59MjQ/7MXNowUHjeFUGHqcV16OWtzrLxWdSHKtnfEjgbPWp3v0Eo9kY
3YRDwm8I479o4fg0RZacafuH+7vweF1uE5tqAyWrgzwIfOMqzcrcr2TBoBMmaHwN
Fc0LuNSE3Ab9YOkubla1GYrGaXzFcZDOePmL7lw3ArR6I+zPOzZ6GNA048jW+cnq
WGDalTJgB74y+WdW3rYuJioidpxH3QVr+cIeetr+Xgop1DEtcgxZk8xM6yZ9B0lO
P7aayN4FGV/SMZdVk1ZWKW4vus+yIo218MbjHjcu9fIOfAenehMUsLRmnFqUi5iD
uh/QfEkUlBLa6W+48leBjxc1gk1ef4EMZuqynTUvTm8QVF15PdUPQq8bdeFAOIMZ
3tVZC8E2qT78hQZ6x7WkTQgpfalD4wiZQvpadsyxrmj2aZ5sEoQ6jGdk4BzlVB+c
QczUTE40df4qHNPFz50zVYzaiiKFJq4BvcQ6W9ErJ5wT7pYkW0kflwLwE3YmmYgQ
+n20QVxk5uWd5QYpFiax1pxbzBLlabZV6jRKKJ+3qpctWRHu8FgaYy3xMBOQxDmU
tzVUQgJQYNtbSFsk9o2/HxGHPQAJtS90v7z9f4CNXSWE+ME0FTGpmneVYZy731W9
uv95ZF18TK9+xIwe1hustLofvFKxQJ6eLb+iSJ5vEZzHWRbrpEyEgOCQSTv4eX2K
wWMglMMSTC9W1qutv1uk8EALTTAQY36jgzM43h3SkGs3NTLb5D04mEN/LfOJwgzU
c9nKEr5j7Q3OvECQGIOHvIbD+dSHLyo7mBTRJvLR9GeV6LmkFCqjouoojuw1rKoK
huZDcB+NDodmpwvwAucgSr8Vs+gDjfCJSOHG1Y/zvW5SWURXE/UMBxENfEsCGzEd
8aA0iEndRTjR7WeKcUDyf3dqrzaVDvGZOZs/x/ycUYGsB8OAq5TjrTbzNqo6Getm
d4LbkqPaijMGqVLp2Msk9K6tbb3MYyLZpBrJN0dHPaoYrelZGUkKeaad/EY/6lmm
mLTejpCXdR/GdvCc1czJ3Bd7Cqkxjw4tIsGtfc97IdJA8VT9eqx3u58eWPyvFN+k
DlAVeEP1udwKckS5WYHsAHdiK4wqsZ7ZSv/aaBC0uSDmSgY9HVEX8QIFjM3YLIMH
iVbkMj+BJPzCbyMxmO4TQG2IktqN+HkmaBS7iJHOW77g6BWkUP3hhx67gHFMZrfS
WdQhbMTHtlIVr5/y4AbhlBTwzbt/ndzhZFFJv6nnKe6rHCk1qD+wmIBkvoio/A6s
BHifwIJJ8T26G4/lvPKiNHcKEkwXn0CJKaH+h0BNS13zZw86//f+w+xPAOonYPeI
dIj81h7G5TNA3y7xGBY07RqNNt6gXP8lANAfepItAAHkZsyaemQf53ZKIJanf2Wi
InWUOQ7lrFuuqTeT8BgbOrGUTeAW5jZXmixpfVwHCTOXopSHdc5u4inNPyafU5et
SqRYtYLi9Mf6Nj/2U6T8Nyxe55m+DgMNh0UaY2ffwFh3/wdntW0W4+i4lapze4zU
L8EENZj93vFv9toeCrmSEaDhXmGx25UaWiIhUx3Xav6GcEq2vwm+Jr0wFl/3p+xq
KaTJvEQDjlt/QX6Kfbl4kXdsUIO1NZy6Wi08FJmDs54MSMsG6/JsCEUBP7l2EFRY
8h1Oy/K3SmMW5KNVX8SOxaLD7pn9u5q6ybK6ZBrBjT3TahoK1dgoA5fVc/mpChSz
f/asUBmDmgurbaH+iMqDS6IpZ3joR+kmdYxv7oyt4QwdEA/d24Hj2BQwNTLlGinX
U4taYc2/3YjBmfweEMKyGht19xc/OQfDa2PskcK2cV284GRudkH2ndMgr0hQdYcQ
CXG8Ob3tB3CyoBATtaT9vrYYooYQs9PIRtyLJphi1Cabnz5ok1tUnlj1Ndp6ihft
lVj+8Iu0iPbm0gsLG9yIdeAXDzup23YnpsXJJp231Mcn9ak/qKrC5uOFxKm4Pr50
da/I568O2GkFqKV3rWukikgZcnH65tnrWnhji7TvGb6ffv3eM/KnXrQkgekFQnRV
UCuv8ae+CIRk/D3DoHCvyVqu6uw08A8ATLf0QzL049iuqkcR2sUfYCGOa1Y0y0kS
vCqgc+pULUfAvynpwp6SHocDcQjDnzpsIdjqdbmQAbH5yauDmKTtvoQGTLI76UcN
NnYWmIyWDZq/gCqn9HxWjwJMD7vrm0w/qEvRWqQacq4Zzd+C7UnDgQXNK/dvpvDO
4fmEt3aSW7C/hwG3SIF9yHfYbK+ZpGRW1y2oZSIVQbTQb/Br0aYBx1ebnUbpDCS5
X8YVU5TGADxtPS+WQ1j2v6F254QHYYxrsgfS3iwPlPc42E1ZWQTvKGvxonecV5kE
8LLXiFVmNZ9WCHIQk+Dk7mgA2nLBDwC69heqmVEgtiCFBwH8BkLyLjlKDLlW+NM+
pIio3Uf2f+WcK73ft3wBPzdnjbul4MF7G9HFWBOG6e+a+/TTadbEneM7t4OeIfFF
UKllwddJPGao453dBw3RCBI8KEDsBYx5h5StqfWs9TF/vmpvS5y2oLuDvv3Sy9Cz
iOvU8DHlh0XLpexPcTR8MLgi18umOHHHU6UWB9UjxR5+oq9RsrUlk+6sA5+oduOQ
AiLBLfdU1uhJwfQKMJ5oD2srnZaXld8Eo1zcPZx6oNg8VOsIT5r/POR59mkyQubR
L9QZRQKt0h8oRs7tPR7bs4lWeHgQuBsQWUKeRiDWM0nNTcicVS2qJXJ4Q8ZA2EV+
YlMyRZDSMww0Oqnmoelgo4UAMgYMHPtUccYD8J9riEx1wJyRwsowdYrox7v7P2jg
Ag71IU81wkJjl7j82N4P0yqLfYOd3V1tA7boUpxAFcmrUX9C34zGvSLU5JM35djx
yBpdZa0ZHQbbUjblGQiwup4IEqhSz+TL8Dnh9QbzUMn0meDPyui3T0kuzSQ5d56q
ajjccZjeH45OTFeEgNxAv9SdJmcyjxEWD5XjjS06SwtxPWdHe17nMuTDi8SL936F
cmI8n2XtHpsBRZxlOrm+o0YYMf2rRGoE+ieHXvrkdWz3HQj0D6RpvZAQNgCtbifV
BWP9wEzWj5U9qm6trclgrGM+xf7w7Qw1//frt+twLhT3HZ60CJtLNpFTCS61PEpB
ysza0lBAg7u90ieIMtztEmA8jvXi8u8XPdz3dzrWf72vZyNIuBsz7UdfJZVqcIXT
dzIcVRy+kUsqs8JblkFdsW1qjmhypukR8GWvHq2h+WkEeBOC4HtQTPyu7I9uCRc5
EHu6wluIOFjEzVBkwuhXV9Mi+30D3X772PEDxdiMP2tq+fEk+3a/f011poW2i/5c
txWNFEf2A6ryB9b27JsXUnpvD4WAJ1hpbkJiEdMGe83V/c1akcQFCowusNmxtikx
lEgYzF2NcWjL9J/s2YZHar2KJGuZwnHHtIrzmoLdo1gFehapK+dOM6Si+qXLS5wn
riZqTp8gQNMYhSNBlD1pYXlprRXVJhSAuEsnErcs3g/g9dSKEzT0/2+JWFOUQaOQ
36ziDrxaLzHjZs8p4qS4xnPZu8y9UjLzRiRO8r2+RpIbgxFixywVgRMv5FFQPtDR
Tc3MEHGFmOVZU6yEp1gSZbJ5ul4fsGhK0tnMOk770aIL4qEN8EfTS1I7WSvbVZO9
lTWSh3PZAu5Fv7BP1luavwPszPJMxWUGZFeD7BdiKWn88bh/o59qMke/HjoYCQtE
wIw9N1o8hwWyl806v/PxnpADChonbFMj4TtSRgh/G7kqdUTKOQD3iWINEz9VQybM
Ccs7kLBkFsy/MYCfYuP20KdkUHzpfkNNu2BucdK+QqB/AscQymz2wHnIL8QiSpk7
FJY0ehKemiGuhqxSMxBlzrGA6xHxSmAOGxlcwxIcH5DkJM534N3JXi0fkjm243mh
dgE4UEwpsF2Ij3xRVzsl7SJ19Pv2XQcRcykEnvI8QqKcp0bXfPl104dwvIv6SgBL
kHtaFs3LlWy9q5/7HgVFsGfVPaunhMeH9ii3ChMziFn+BUSHgwrm4DcU/H/QQ1O/
4a/KiQCMpAv58nSQXed9bppGA3/XhQI3aLE6u+GWb/UM14JZNdWhqKz3iV/Qsg+R
q2e2lPN7m7FTY5S8xkxKQM+VGRFXrenQjaVIamqqcgn2XotDTiU2U9L4ObrL49rz
T70MFpnJrn/pn4CNwNdDsGjW6GcD5s65eaErsaPCjaXd/a0saEVtJq20/pM2Yrw7
hrvWKEHQMzsPcBO1GlKwzoGbvbKn7y34o5P+bqmExvSOYUW80Zn6PCcujKuJuXdQ
y4AvQRCZyP8Crwq+wZ6usARmF8oOjqfZwWB0CHItEUW417k/+pGX40Y6mqgimdTv
fUhioTtjvrTEpJlxZUr4nMJMPyyPHb1C1zqN3Bybs0s/mMfAgvTZTnP2Av5AJiTl
yC92L7EW4YyhCvOlREaP7N7yj3gLfiQIU3DYRo30y/XrlvDqdTeM4E4WvToQ3XZz
SwTEuzY/e3RrrGA3FEk0kd5AhgXfhJq9gSEUFpBJCx6TOdg+4vHALsaudnUaAFqG
xzoqMCO1qRp+vt0e6jcuMsbLYH9AEhaj1JR24TkoIHJX4SfFhYbw2l3GPXENrnYx
psy+ifn3Ta6M1xdkJFa2g5+77Mez4oQQniM2DiqMXJNW9UtZ4ripENPMdzqL5nhM
VveeJ28LjVqz3xKBvTCtWXtnaXnSGoaEKUkccJ7Fu6FIZy6YGYTKPhtpqJXQ9eYD
pjhO7NFEXLue3wn8tHNNcptv4m0Ww7GHyZWeQ64Ip/IUGcR9ymAbfNnDjKfyvnBs
SE2CIipA5gFEx6BypuTuqcUxgm2R7Dj5cGjhk2DGo4FEy2rRceKsj++BdzF76eX0
FumOwwfvLZppY6BU0l/5efsXTR3Ex5sSVs9mKnfHIsatYn1yqaEEoClkuOGUZtpM
Cf8zImmuYFsAOvjpDJgW/MULpJ5/pLVLc7gOvyzBwNATju1eYHn1/oXILbnR6hEV
G7mAx9Vw3l33bUSne1XMYo1dK4+F+qgaoAJbFVLqdr9WubARfqzo5MNfbkkySPni
brz31PvaIo91gfRHJMr//8umlL20h3910cACdwvl8maKk/4YGLwQdlwp+Et7nfkF
fvIs20w2UJ9WXtPQ50bYts5EWMTZQJq1GB+63xYXVDlKlm4/07eWDmSx+WtLj0mM
jPQkfpWXMqWSMfkM9Rn5Ix7JxQKgT4y3hjsHyDdPnBjaYKcDad7eq3myBDS57IqH
llmpkTjywg5WL/mBdXH0icIdUkr35yRJEJZoBsPyZ2+FN38yh/VRy085/q5GWTY6
mVy4VuawvGSW4+rnSHG7t0vKXT9O9QkF73RWNDopuS0vWTEKKjdWIHZV76oCUKUJ
CBUJGqG3CM51joPTjOX2AvRZxtvlxf5GVy+XFj3T2VKBzi1Pn510t6ydvssO9Vew
6BmsgoA12R94gBJkgwA0istDxC+B/3xaza0sNL5OY8Per+3AkF0Ilymyzg87uBMT
l5F3kF4lF9EDZNRcRdU634jdDP/kGXDTsU6DVaS2qW2d78RlysjDRooIZsnccxLI
i66BbYv29D/miWrPlhKdlIxKy7MPnQgEw595yPY5PzB+/NlIfX37K3xC5xarzl6k
GKocBLQtQUqhP+MpDYIfb8Q0nkhwjrzOb2MWdZ3hQZRWmrPh/539XmLY9NR0i43b
OQ4OBhYeSM0cJTUT9VJxggNPFLRXkVE4PftP/ooRuDMYcqaOrmOL1XJh912kkUWy
VYGWqdikEfdbLQnsETiTC+uuGvNM9tEg/MFKXJT7aI5jp4S1PAFp/WJS3pme9Lzl
prOBwyRlePhpvxAUFtw3hOQl1hgZK3Sbu4jbn0CZSiro9FksN4qK81darGtwIyCG
iJmMqz89AtXhIZp9f0WUvGUiQVBA2GKCCmuUhPDNas4D3rzFLYK9HYe+G7qpTlNu
e/pzwJoB1wKgHMMadHz4uNzadeQzQIkVJmSjaMFcWaC8+MTEreijt8+F3zC4VWKX
vrfbK1bBHlCnlssnTX3fbFMaYF+EnD1z/scTBZq/H6EfEqkE5MrgfaHe3spkc9V4
JrqQPsXzLImy17Odk+wGXTkFu+Z0I47k6xKyK8WE5zTc5tveE4XctA6r82JHTezd
KxVm2rfcuqXLomByFV5FggC85s73aHOoSz3TcFXOG8qOB35IsCG67GWsQNZP7lpl
agEk+O4hT979hhDNtHP8RdS7QmQXXPwLfx4Tcc2JKQRXuFyjSBEsOswmWSL+MOwW
edXM3B0+X4bcAznRnDZ6b3akJmRFHrzpPvrgc/zG9HeDIKDeWNxUYP5GeFkQ/G2o
fSRCq9Fr0EopHVgpEmkm8YLajJulf2jcQ84gsPKjgFPW0KUjFU3zmt03YSPY9MaA
RvZ5XE2zKcIDmfYOjfXFo0OmMFEuW3KR6MJ+BCzUXwngF5UDy1Dxfk1ArRtWfZZc
7+AQouzRuhhb0qWl97j3qJZVWrQG19P65RKrGwZG7KGJuBINkvJO5OhH00ZBIQXh
+vN7FQqrxLts+JLnk9QKhLvteWl66uN4awm8Ueol4oAMD6G86Kz17MYLYY+6b804
K6Zol8E0q3h55Nac2OVtVckVJiInUKS7BfBaeWRhEY59AGClC3ppPxp7vOYCzqPt
FiepIWMZXCvXpESgoLiru8hTis46BarQtOiGIRYgQd6oKj3zQq6W27nT/K5859AP
nle3b9J9B3TBGqiiZ7yTEIPM2SgK8zzKDbxLGV/aQ2YJ3d2A7/zUgvEPAed/WlZt
r46R0OMnqBArXXIQb746v3rG/5yYHMWjGm61Ld+S5/45ANFQOtqTYynNcvYHK9d3
ezzpZao6HNtbUnOs4famJ27dZqu4gH0EarJa/eXIxzhA3lXisGcA06KzCW1JbddH
CpJEI2Lv01vXDuuJOHTqirCOPC9nIMdelW5NJ2YCWA2R+hSP0ddeIKYyZGTv/VTL
qV/HQUluu1V0hK7XfOLluh3Hf93C8o11SY9iePzJv94YlYrxcNimxLqPlZctgXwl
rCfOFVoQ6Avs/xtp4Hrj2ImpOqMMeMFfPnYgHxQxgQRgrEpNDI6vbGk3Bp6AdT/m
5LEcu2hEnvtArXiZSDNhk6XMXRXZtDDFDA9Wjo7GRGIOpBcCozfjAOSNlFdbMr2X
GaYItdOMd5SMANMkQRiNa8Lyt+Gy42LHuUGMz7BHlcFq7SlzQJuKTSI4sapXXccw
Nkwm7xs/OSTKcii1SzH3wo+FP5gO/VJSOyKa1E3iMOIvq/ZvjTNfBGIEDYm+Q3Zn
Dn50FNvzImguj6QEjlKonR23FQI0n7TLyrvNOvETf7GlRoW8futz4e7TTH8qgWfG
LKqqcU5XpkO6XPzy7Lx9Kkm8cg0427IKRAnAi+8peXjRTVhbdUFoTt9EQ6Lid8WC
HBvdntEwe5352jniqk4ID29nrZgED1TXxbWDaioGGRAplrVsuQZT9wJ+Ollu/jF1
JzFHo8rigG/U4BXx/t6xUwCrewjDcBeE4Suggu4ZoSBLLbrvuQdQmGjiXTOv0v9n
UwSWio5Ej0mwn+sTniaQxr/M0uDdtcdTRjQ/lSNbvvga4qgR/WHtjIkh8TgVvMm7
Iox9BIa1y0c9N30+8SvaRLkGJA61ok3BonWoc13gN+tA471y+so6UkTvWKzEAYqr
8PnejGe69YgseGworGd+0HtoQ/osu7ddHrmxvOOTCIgDhONpKMgU9h9Ifbc4siHu
ruJke/snYV39fsWUsJnZM8gWi7R7VD04ahauJ3Fg++z5HVwL2v+W+CFfqRTFbZWk
g178oVd3dkYvBGFxz94f2AjLIAHwHfQ2oLvE8CBqX74pnXJnI1dau6Rgn/9kO5GB
Q4qnBR0YbDfYJT8h8ZU0I/wlRzRcV8eble1y/9zw2Ty2ogbYwGYZTdg0q0RVKx8j
dDjGYHELdJVfT+0KSdVXf+j2L+xD/O5anJN3l4KBJggnHYNrP0EJhXsCPcCZRt7G
y8CHlgeJFN+Q4TjjJWg8YypOXuURm3g/rA0S6k+2q/CHlK1DdTyynNkvp0Tmw4w4
zDNOocOSQ0ig02BEARPyQuGimiBavPoOTRDSJ3mUIWoCpLBiGWf7re4Gcn6ZX6fd
8SAX3y95PRlzox4UxlAThHEZaMHnpkH+VSxDjyb+nufR8RwjSKXuyPwo7ZykSrPg
LKp3jpmVS0Leky19vY7X8ykdoVkFVtXIQ7tz4nntMtOkQX79PxzNFTeyt9MSk02D
mRYojkihU42O+2+VwniR7nsyGpWTxTIu6jVwhqw0NH2mcUNWDQQjCrg/9n5mf5Id
jTnIVVigeQ2kPR6LGlSzXUnuBLKCG5I7C1opbYTV+Fhbo1jYJpUxjrVSBU1Pxu48
r6oAV26NWFFu/CXP+RlLbHfIocnr6VBs2CdZYTWQG5lYeU2CHyBBlZkMhZ5kk5D1
6Ds9roiZGvjyu5/moEsolnuZUNfid0wRpKDZ5QVCosogWrTvnLeQ7cbzVfjnI6y1
RfTMjTJNxjbZ1GTmqRvhQJZs/G87h19Xv8dFdNKTy3id2uPw79wT7m78EJO5HbKN
QmSsKZfrP88whHkJ32zwU9ANZgI/mmeAI6zr3t/LlduodA23gaL0MtiHy1vsgm1d
r49V6RQ8KmcN3h466hLe7p6hdLsu7c/qIbKPZcoUofVP18buzAWJAw5DluUso52z
1+zkGXaEj4mpBY2Ogdbu8mJo74fxhj9UUk2uwPO4LZ3+IxzI72sPtVwTilttbJeW
XmV60wPNre+bIagik08PyoZt2CcEPgMLmDsNr8uMnMnuCY1u/aizyN99ujUF7iXK
kqJfZn3bpH1uPHph6ssACS5b1P9IPzs/Fk2DImB+NFTQg3y94VT5jncQMW0zFfXq
9Fq5nytc6sIRxeBtKIE7bliKXRqjKfmwz+xKq3my/uAl1DEH6yxXl80IuPLX3bER
2+6L3+D1F/ZBwSCCQ+87DDd/Me0BfdbtG6YoVVhoWX7OKKKnN7clSGyx3MLmTGMd
w9SUKc4HZq6GBeO2ajPR4hyryoG+gaDhJlsBb8S4VSz+2c6P47BbsVs6jhVdPiuf
20eU1tneDZu058SdYx4tcteZVXxgHumX/UPiZ1xgRd+pNgg7L9jDmK/AHFy8q3r8
yz1AdBnoSB3+P3gYtEv0ZiO9+xK9bIlziX6ZGntel8LwZnKWhJpTirE1DAAtZFgm
vGtvIDojm3Eg0u4+3qr1arqRRejinoKInOEB24QDizagBeSlH+vMiVSwIqli/7WP
1Wah6hLtZ9K8ypre16B8y8QZ3udFd6GVphlZW7qwjBtEgUnKKVM1dI4mhQcg4oUB
kemWQNLELwgST7OPvA8i2fbrlfVc48IAphIsxq/GCrV6pWZkol+cEAmMvpasfvye
44m3rhTq2gIfqEE6z/yHSHHMUlMkEH76QEvZEfirtdA4xyPL+LrXcizK16fkzxfJ
+lWWddqd59FhG9scq+ZJSvZQ3e2BQYTK1D4gypV91fK9NiqapC3EtTfZORFrVq/w
X3s9yDUy+/3D4r6vqItpuwcZ63S6IcwsyauJVUH60NMejNCuXpOPBWE6pWcvQVI/
R9bL85khS6Qqc7Bph5DFWrwGLyb31S4jRdsBT5r8MhJUuXd+8KtlXL15h6o1Ix5l
NeWMx2PObjeoNqgB0Y4KFnPJioO9fc75eBxliw1R8XWjDj00sNMTd2Od84bttM9b
/K3BR1fvDyx+HXpcA6D4cQ73KSqlhSTaMOdUOBTfdrzh3Fu/8cQyDA9Z7nysHcsA
zEVV4a+SdtkUEaDPjAu7G3SFqmURpeTJurNvjwxpV0EU/ltp65QseLXAkuZW5Oao
OHf0rK2pY5353lR5sk7QZsDS/QNdTotQ261vHP9gIJeC+KbWmAErbvNta3Iq18Py
wrfvoymqQJqb7Ttftc6gC4gZNx2USyUGAwU9tcL3Dt2QWRJCH4A45XWSwfvmt2cx
aRc/9tuZwDGBLOh8Qgy4Qg/5ePv296uR1b7VdJnCQ+rTS9pKy5iHS+g7TPJAMPdX
6Mn7cTY8z83NaG60gq4z/yiH21z83PLl84lc0l2wdcTTA0c1TELNggHRaB3YWnPQ
ZeTCy9G3r2/FvggpgpBM6HqaouE8C0xC0jlz3PBcSD/Efyy6G983HXYP+AFazMZd
mt3Qg9vAtn9f1KmnFQILYhBuS4MSz86DHefAs7Gipsiz+olcZHTOZ1ne1Fk7PgaY
aiPLsKQvk5unZjYuKS7vdlt97Va9qJqR6VW6goMI3Y44rPcoYbQlcbAorpZV/3jn
6mP5y/c+pq4b25TWYgsXMyfLfp7/25v+oMBaio6QsGIl1tAINm3LUopDM3Wc9uAc
b4gNqcxMncycq7cxz2pBLRPoToaAl0udUsJeCF1iv0qFnme80IgUWVMUsO/YVcvf
xTH/l6+Lc89m6zS6DcsrUFUsZYIHuf/bFkYts7UBuKJ7f78w7uO+vbpzd0LEcvAr
QHoJxrEaM5NCmRthCeL5LT2gL9t2J1DJW+fuHwHeKn6p7AX366zwFff6WSG3wsiw
puXmx1xy1HW5uh7C8F8Ce5pa7CKh6Hnkk0gRqjHjuujuvhQ+3kY5DmGvHvVfnmPr
OldTAGiR//Ey3PRp+rAJC1qKp3mD4AbMXK4Oym6A0M12Jp+yqR8PYkcgeljkeoIA
NOu2N/2EkZVp2+UnpupOiX31WKVHec9mvY63Z7wzn9SzjTjYx3g8TnBZIJGMXjFE
fkUKF2MIfMAND1YRQmAjz/+ky+nz2uHmhsvRd0Na/yHUy6THmthKT3VsSM9XkYZX
azylgqIhRTi3nFt7Led9SeKbCxPTJ79W0pBY14/KiMNeGuqxu42UXkZoXy6UCrfU
bkHae1QRX1AERZmNSxnnZmSGua1MUOulOeh+SLIk4YKnguOdatVI06jMOtICvi9L
hnSGkg/oV8/Ubj3+sjBwqNYtyxGXUQMWGu/3gF7rdCHg3cbv2Qhj+fkA3a7TR3Ky
T6u8wOFAMVzOZY+82NF0rkkQNm6HcoUsqtx3QssuvmkNtwz+BbU8AOUYUO6uoBwM
6QWZIUr88ZRfdvOdl4LKlT0mXkJKdGcxHDqcia/O+94H9prpxon5wfqoam36dzkI
8H5qQBDVWdpsW1FOBtWAAePpSNWZw+LV1Vjt2hWUL3gg2h9hsyP8fPZ9k1jaByK9
pT/pbYW6zu1iZ8zwKCL3C8TxNTNr28t4zrh9iz7eoOce0Jke82jfsZSQUi28Sywo
vjotq2PZRjFNL6/iioLzGMuBi4aGA90SYYYQy2Dj/uTxCp2bWzgxmynQV1aw8RNz
2iZd5k93byLr/AKphiKbuaGSqu9/LHzV051lZU4LRqHRSwsfr4TikcUH1VSf+Ob6
5qKNAWWDGWNWKgDgkwl7UnrDa0Nj16rArKoyigf85WWmXzaOY4sAxUtUxkCuyJXV
cjgZ0JGDbrW9MGGQLI7d7WhBkuE1xmTrKYOAEj3OsKe0oofo77KVvz918s2Uwc7j
yMhEaJUA1KWHEWTJoC4z2xU98BEnCjemvYZnr4ETCMOXbISa+c1Evt5TXcvCeMz9
xlu1WPpt9Xu4xM6d+zX2EnBJiyo6BpSuCui80qbaYAXIunaTnum4nxo6/kl3jQn1
eHDAkMkezTKNtUPbkQCNdNRC9J7N0ifIF1PYfTOCM5y8fLO064O/rp+iSNLMxYJF
8r9heqHvXVZtvmuJ7C4ojrgSHU6aOwcaPdx3Sc3DiVuocn++afU5EFhia0a5wm4Y
7X8BmYUElg/DnxKLRbCsV3nklKDrLHPHOxdwBza6L1Rytt4o5FyD65kjDufpUkep
GVuz22N46pdDAO1LZtLK+zeZfGhC3wdqutf0B+H0NSCkYrUkhcBzdZwSFXWR/9rc
0OyjaBUgIBe8kx8K+Gxvp7FiTCB8gcpN3CarG7gwxQ7spQWQoC83k+v2Bi9mZJ0e
M6nD2oRNhWk2emSzlqnYABA65ODFm81SeofMT+CPMevroUYWYPXgUAci86ilTNBd
mvobN/KQXZ0hyVEQwuJf/hwOpWBv6BnvOar8Fc78uTHfkQzyyKCTjC4CePeiyziZ
3RWhg2+lIUmSxlyMn8qyA9fzXNGqJLjIsFEuziKP73AhbM2f3cDkdhgb9l1w4stD
cFIGEFJw4DN/17tARrOtCpXbaU2cefCO+TYO7fuuPUEFtjdKIvSoBAq457b5uICR
f8MWqnun79QkmNB3tzAqwUud209WTg6lcbtuqp6LCTM+HPaNOKfVxHexBdhuP0gJ
nZsfCkMYZkM10iaSbtQ8/FAPfp50VuYPejHIbidAfiaDL7CUU8+JAvvVAH43Ddgm
ggjoCZ2mO6FhN0xjyo36xzcBSUp/wT4FNSv/Gbdz6UTZGoCfJK73bBVuUpq81v2x
po2TNloPrB/Vh0NS80xhVS0kx4Ct/JD8PnXiOsm9Uxn9Yyx5kpXgJI9JSherhkPO
LkT6khyBRBicd2RIEAa40ucICzKcMvWn+8u/hwa3QSRqrLkC2rDNg42jsYCL1NBd
cfWxUnu5vPmPzLqGksyW3B/lppHJaYBaH1VnEtI+vdiZCBuQTs8eCz6KsTo5QO8o
1MfzIA5U4HTuPTE+8SZ8vHl7LfmCNBLCk/YHpkEKiqzUKmcv3xOoudSj1OWhhVlJ
gdTW8n92F8wrnwPG78sg8FTmJ+2XsPBxFJSa4gDBDFt2SoLtWXPtXTa/Widn0UJ0
9j9pSrP2kfS6ZBH+GFrYzcYUcfdpyz2sQd5DZ3g5eoDoAVwHk5s8nbh/PlL2zRVo
HJA8M+pRChPmVXbyx3r66/+0ogu8qy/eCrdNyHwqf5Dkauhy9amIQDJ7Ed2iq1um
liOsV/Nn0BLp5wOAsIyv/YeKcK0RrQLa5DY/gac5KW4F8FZ/kbSNy7E3pPs6WuNE
k1LKoeqM0LaCFZouUih0Te9PgttPj8c+4d6ktdCkXRkZtfnikUklKsl+iI/yeL+t
oy/BKWfigcoJNQXheAV+TPBrHwVJVJ1GxV1JqvaEQOnyFupg2ReXlFIRaLKXapfJ
yj+0CAmbgfGqo6pOWsIwMSrv7ML1V74gABJyhyhc0ShbuohVeLvYA9VDm3WjTb4j
L2WQepyhvv7Mw9iyTiykJiBjk4L6laPQtBodI0zUsUL534jFphfUwfqC1WgMKpo8
FZKsIuG74KYYNrpHQTBWFRb/E2WRl2y+zbnvxPE+1rrJzypJVOxpy0RvvUqCEV/I
NfCarlQ5MZIZ0DeikGjQtnerztaxbrSsUQDeEEr0vsFiIydU25EBstI5d/F6uFry
nOCxfAPqG9IQLjDwtMxgN4omwCs1dX7vP0uPAzxx3iA90xS25UGrVahAPzkEzrww
Au7ctJ+6tHd96EZDiUQFBWd9jd4q26mcULDUZrNaRHqnYqwo+j6ZEM5ZYofEYxEw
xLKhgeSxmaqSMAhxoXjyAckVHSz1iubTt51Kr3q7T6qrLmvj6i7nCV507zEKgSmM
RNjN6RM3sbNBX5B5x1E8QwmGyV4PNB57lKtedn9eNUCmSg+XJRwW/VLio4NH8Zvw
eigUSpe5ofqqEfFm6L7oDpz+mloHkciy38aNGV6H2dj+jJ9hDJcboYnf2wDNb4WK
6ywqLrCkuRO54MfxWtlfdgyHYdd4oSl5dG2i4c6Euu7TP3Ns7d9RqYa9uGK9A7T3
FkD2oEEm3b06ZTkqVIBHnaRBQE8kaZ0en1S1209V3b1E25EF0WMEUUEUwj1Wl2Uu
r+KtSID/7g6SJ3k54MRyadwl+FPrmPyOux50w4T9l16fODVVsnGw/twLgykY5EWa
qYIQNK+o82YMvdxnn5oahl3UnI0JNe+AnWKAfehfHi/u4s64iE87XhmweV42xgLI
f6SBbGNi5DxLQ3Vez7jB+N+JL31qnCtMfdAiLPUlOpLENgz2lJ2Ww6ZemrmKL54Y
hY7/gR6eMj7W/LIJMvo6ndKs1W0n1hLWTKm7DKHqxh/p2YQEp2E0c2nroPPLCYLI
4wPZsWDUfgsnv0KYIlfGI5oS7zF+Oca/bWf/Z/9/siY24nHpmPjTsgRRySbUZIsx
WMEo4yztGt0xsEPbzoAt/CZdjHkXxkIl0sGnPRRYRTRunY6gmBY4ClgmbDvlsTqC
O9fqmqz4pgqpIdvcGI7rShBu88MOsd+L00XG92TnaBYxnCH3ZRPtZAqsLaIYYrgp
97fOyUjwmbr4u2PA5lFL94qFUqxXYlLxJYorMVWKwLHUA2lgAxwKFAVUOW1vfOBL
O2dg+ksXgr25ahLdSEbZyus//sO+9wEYlYGVIHDfD1Ye5r/FyiV28p3fYdhWJfsS
vKu7gZX/TCiXceGobGpYrYXty1GR7ugblll2GDQ490VkG3DEajvSFCcy7trWRb+9
ZOcc2g5aqWi6HuIuPX681XJfWMXHSF0ljsiem0GnNG6IZxYADy/rVQzqCO0xmVUr
ulNQKDHuhCGVk0Klq3YYONfxYtfJUfE4O/Mc1edqoG+MTTT/hmMwHEAxWtEOh+kl
JuXa6wKUu7jeW25amFeN1y5V+NKfWXCbxWZG7m15P/0rmF+XvEKe5nMNJTbLnGJH
D8Knx3RP/985vDfY9f3KiImsje1vPqgxE6ZoTEG5+kmuxQgIpe4YIa34lchmUto1
2XkVfNRO2+32VVQX1LfQMzAPIaMiVV57c7E3yFvW9t4lGNM2ObzbNAKtfaaX4Ql1
2giHFk2LvyVx7K40PEUfUK7dp7iAatFSnRXDK+YuDFU9V+w7kMqvStB7qr+B1aAE
UusOF3RLyZrm4eWdGDPoS4Do/ZeydrxCnLbzUGy3VNThpUyEVo/uhtREiePS30Je
gs6c8tca9EI1OyJbMw3VZSvn7hhl1rCBCv8PjymybcBV/pMJMN/g8dn9xCERLZsT
x34P73i2+9CHdhBsrG/QJtnroiAcIA6o0cERN+i1q3D7OyiETO7QBFhzHaJHSpZg
mDA9ShUt+FeEI9UgNzZT0swOIDWIwFwxRWGneCEu0/j56fILqaLa/dkaFXKEcLLX
ile+CIaNPlyTkGysHNt9fhoy6jnQ1zo1omRl7HBvsuvLwqR0Qpa7J6XAhwPgaupO
MukS9Mxvmno9Q2EpNnqMBciBp0j25wpxJXaRjv8OVOaZIG47hLzZTBPrFjoAUN1L
oD42vUsvRCO+CMEklPxa6lN2bPHBp1vGsKc2aKVFZAK9MmngOd95ysoCJ3Q8Zhw1
W6M0QomiTtzqXBmVYOstKCL1D38FkcpV6FmreGGU2hYHgQ4H0mS3hk1V0uMVc7FO
+3rJEUILjxQsU4cdzOPIAFGfjPP1Z+RbqUyp9aiTlzMYLf8CNuB888anQBJ5T4Fl
GuoBRpvVIBHPL0hSJm87dpd7E4dtwo5Da1mbyyJnp2J/cOl3Wp8kaA5yn++MI2JT
bJDj4h8+GnclliNwOlNuxyNFEtpnNFo67UaLodPY7XQu/XcSh13TpTd9uB2eo02n
BT/n3Cbdny3OwFpJMC0q+LAWDMExsh4IeqGknab/miFmAwD64w/oPkV2iMvIMhIw
TyB3wAgQ9xrkA258CxMYgRtvXBRYzuzLZ3rdlnmq2QFoxmOTYpY18St+J2IatpTb
CL2w0+M1abknZ0DZQK7vuwbwV+rnTkcKnWPI/kgo989pf+qbsrdoaiJrtlr7/ffy
K8coBHwIJlC/mgyeI+vx9Vs0Oi6aJIykFO6kg9u+2TsCxcB7Y46LIH5LqLDiZpJ7
Dt5SzME8WHOWFYZcsG6lTxr9GsFjCfc0uTH/N4ValY3BNyxlUkBU2SW3s9N3NH7u
D1c48/isk6wFnOeLMkRcsysXS6pzk7XHycB23wuYy4lwJjHMn+c6ekQaOK/HTNo9
xbSxxbxZwCiyXsbpw7O7ApTRtc2d0C+wwBy9ZnUhB8dE5r+zP6S6P3RblkHm9lz5
fYH1cgqsKUAVJd+xqnFHPTQvLqf2vLBFwnQySe+aMSS1XW4MQQpJEjA+2ogoDk7U
tzzlVhIDyB8PxCj5xkUI1WckpJ27Ip5L4cgSvvrpHafRZAQoPjPLmj/GBVyzHCK5
BmmrajB4+A7WlUK5rPTcziBaUBlBjRXXUobpslgf0d+3qyf34TQePTatscrbojVq
3BTfaW7QiTlKICcgsAI+cB5DfeOapwUGlJVTJU80BOL7b/HS2WNLW6UJXmWUu6cF
Wni0AxKThVQvJx0GUEHSpcxcy/PiAIIWznxeKDEu4KracWmoVgi3NGBmvTFKpsXn
4NcLR2glwQuEVkWDUCGQnt1str0y9pVgQWWZgcfbkrXzGRPMDQUeFn9hb3VhzQUh
bOZETV6f+ETe3PYqX3SLeUsAQZUAw9b2GeLUVjZNsvBCk/kFAGDU/8nZzqJk93Os
pdQ49YhFhPjS0MhdsA1prY04WBKSv0Q37zWQOOSmOqQOshHWVUeL/xIINUUNK/8a
79vrUfV0xL2G7j0MwKI3q3EBrvdyjYCcLujNOYshAf60mMp1N1t9o5FpK5508lKJ
nitewh1KF6/6BnfbaFtgTgzv7pk27YodDfj98LwVsB9rIMxqPgAjF5cip4UXejfr
WUS4jf3CL1VFjqF8FrFD6cmXNgmja1HFoKV/DVdIu/S7g/VIC5VBlji3qako6EWB
djvjvJ6orGCdRL+maBTU7rqnZnjxDdQzTme9NOluHZCAAW36SCC3rB+FRjAi++EL
BWA4ybTE7fE7kmp9ecGzPJx7k+YiRVkpuzRbb2PD/syEWyt1rReM6QJ3So3E/oam
JSQYONTETomGx2NCF6+lugd+xt1ldyXxM3XIWuB4LUlDhgtWcoX+1hCkBtENVF8U
YYe1vuKgwb+NBrHrGxcFBhsyKhDrPMQtw24owSZge7wvYOdsHjKT/ARunNDBwAwt
kecfrFi/96omriIr/iNHp4cj6auySegx71rrJQVwsnrfKsxXUOPGjCf/cffGzt97
3W2jNiRsaI2siwpWx7IROn/kJkTPgHCdXYgCPpnhmxsd2zsp8FqSlsZDadICk9bW
N6yKnrbGo6LaBb5QUuMzcYPWolEuAeuHBm1Z7NGnHDm8Q+CSUqa3AYpFcfGXiZJO
/ABBMF+Oy3e0EdKjK2+sX4rmsn+KmqG2RroEcC6xfvCtDRbOoLO81zP7qRhYuKo9
N0o9lPbhgzhZI1lF0CW5RH9vosNe59+NC8hUoIkaOEim09+U7v7JOh6MPbtPmJ8l
p39nfZhtU/5uY9xYiYBYCRfGgRLftXeqrGN5gN5olCLk1TVO2920l77P6m656J+2
i5lE4ABgUsvvB3nfmg3LrKPB3uYl1hTmoF0XhNb1lpb70UvFMg42x9N/Sw+LjX6m
jiMMlKNzMHcac96cuK7E2c/QbYNJRiPvDy9OH9Ryi366tGall7NQ4aJk8NZqWNpY
4pEijv7OHXN53AoBE5C6t3iA9zRXZK71mzrNKrXAm6r6DekLoGg5X2jiN9k6TlFp
phrdXJBbDNXOeiQ2pBTou9lHs9rnDe52zBRDniSrjmEuK4fxbNaVc5RUt33vdWIs
BoQDavW3diVRyly5QL6o6Tp3hIYupwqJbmK06C9gqJVe9ziWktb4+jzNJzkfEFJU
4ADuWbJBx175ORJ2Es+MQQXd5Hr5qDsvmUOv2+AzhmTH4asHJwXVI/ZTvZCab8ZJ
EItSV/yX/yXLnGsW+ppZMouI2N2lUGuZo3EXTAYuR5zMtfPX9JlW9h2vKLJNubZ7
sXqLPHexqSGdXySTXHk4jz2Ol0+472sWDxiFNno8NRaLEKztjYViXXlJlhF5xt7d
oXn+f9RTTHYu8hWG/lWwtp8OBF/+zCZrWmfPxh9yPYmM40nGc3UEXkFWuYoqpFWK
wTUyQYS2jXswqs8QbiV3DbEUGPdQZUM0TAnpmOe6L129coaDFXA334f+UYc+nkcf
IPTARRZKEpFAWZNmmliU0LtwUT8Rnsn4TfqE6uDceND5yalXtoNhDwNatBJSFns7
Hd+usE4RAjeO7zckHXdJK3WqQWMjnfhNWI/N2OqUlfiQ+nEoIxD81ggAHnokUt5g
UmTGvTk0hBlfBKTqODh1VY0/Cwn1jyDPo0xCN0C0bbDkbQHwrNVBGdtMzNrmQiIr
vMGQDF2CR90HBJZHJSvqjJnjb1JEcB0ym3H48hQkzmOHrdFRfgsKDuP7IOHHCs9P
le/YqGGJn//o6TCeMsjouHP9sKA2tYBM9xgljlPcP8C4lNl3nqtrn6fG01CG9Dx5
GhXEhTcZ6RpdkZX4mVkOdmr3Z33QyADQV3t+FkgD3mvIKqcIgQnl8AOtdDzBJ4Xl
0dDfqOrq/fiLXdk7IB99s808X/rI3Fvm2CQe1wpxz7SjRKh+EmPHyHkEDq7BDWw8
l2YdCrqGIGazNseFtkj9zyQRSi6FlUy4X2eYp34jjCpZXvE+UCRK5ynojAtzydHU
sxjqjKXToLeLzn9+sADrZ7DCQ6Vj13YGw+yDnn1sKtW5hDZxb40kYd1FWGQA6csO
N+a66MFnwhDKYD18Y2me01TDA0WstR+v31VroRe6MJZFKdxBEuIvvsGGAWP8fh7v
TuZAYS7WoPFqd+cdAj0HGAcam4CtrjWNr55XK88E4MnOMgY5GTIiUBfkgO5cqfxO
d51gYsw7sFUugN9c5utJNWNC83Q2ptepeCV6Tn3aN7QKdKl5T+tW/48hREDgUspN
T2OdDKuUlAEd2DxBlpUF2vYRsGCIN4VH7JCTb+gZ9dwrZNoTYSIf8Xob0e6+vg97
ZMpb6uVbFwXWuJYnjZtYGLDFArBE+emcgENd9FuElE2XrkfC3mUC7O5OGkSSqjLy
tkeDpzi4/TkUF0xTd2HiRlp5EBieJ8c+7GUlrg5InprGrHwJuh9chq1lq5mPcl35
RF09VrGAT+MSda8TuW7zO+399jMowjjI/jdOUSxcxqdwODz7xsBfDkr6NziumBnr
NbQnV5qTBmhZvovtOu9j8DqNOLISbZw7lglJ7YpLitMfMQw2UpuKnPrPd8EBDIq7
x/jG04kGnX82CQgRHHUvFqGWW3U9EpVIBeuxESnTA/Tbu7eFtCuH+IZnRCzBGhru
AxojxJCDghv570Y1zvPtCFUgIH1XHyJhTA6idH/oaMipKec6yN1vC+4ZzEdnZthd
vbz1yLAJE4ej0NFP2zz2OL6/PTXVzOk5pIHilunDDHAvApvHwmQHhHlm36NhEzu+
7GLgHaYGRknsGORsXOkDZB3Os/JvM6yRI/UeG69sEF7Kb05Wx5gj3iJ0FR3zuviS
UijZhukEk7qzKlZVMJXweIrZxkqVz5U9bReD8YPQCBpCJ0JqvKF2r88Hpw7UWrZN
u4HpNS7NRdpKz3niyD1MP1Lj6CgKVaZefUYlJgqx5XGsxQFptq0JNhlpuWOCC8qq
qrMcHqbzZnQQHkGsRcXqkSnllwHXvcwJuiNy1EVvY+aKvI13jN+C6eVrFyqh6qIC
PzPT1I1svf9544kP5znkaw==

`pragma protect end_protected
