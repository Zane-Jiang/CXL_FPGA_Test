// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0MBWKtjiFcDa7TFbkSW4Ux8pXVZ1UmRsI6D1jA8D9tKHFSSul/Tq5CXZjL3V
XPaScBJUmkXOnLqabiehX2dHe6koSfsQQg3zUDYQal5y+t7IyuKLpdUpbcNO
obOKNvO23Dp+UGKXwOLdkDAJSN1+zJHa2TKDzSFmLMt07N9zK5AhLykQK1fy
fItYpvjDsd7J/bZV/E8mNlaevybaHIhvpGVa/jD/EhO4bgpvsq0YSDsoJMhP
CM9YdAdLVWzd25joFcLO0SZwTux6QmUvKJbdBRtXOsWCrrNSFusMocu8yA2d
ydUkZ37bJ+5Jn+DwFkd5DMxaoPUdoWgm2e4954eoNg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xh9Dm5VFovmk3VgyzmF03CF0D+On8DOQXcDM8BygjLZGUbuBtRrraMcRqPSL
Ag4Esh9m5oFCZVOjrSasBbyt1Whq6lOL8rnh5LZDxeYNYBHv5hmVnuYPUTwq
QQntKzB8lCuMLgM36Ia2hPZmdGArITUVDe8n3oRBZSAHomzEovbTecIlqR5n
kOY3CWcaVg5ZRj6kP76rMYKEPQIKJHaeRK9c6lt8qv2s9+K6xCjQK0YvJWgo
UBgA5rKqHIZyheEw4QkQbnl8XNlwlLJeqqR6ESaxy1tSiuFs3b7JgjzMuK8N
bnAeJK66ah6DZp65BglsmryYpwZWw1e3ilXTGQc1/A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
f/n0iwczAu0oWfrRmZUXTjzxBGlihyo/PcVuNw1kLwmGBJCwrY7TBISKc0x3
rh2V5hMYP2RskSW3BOyth702u/l9PRn9mm8ytj3Fd6dGdOstEbF29B7bt5kZ
DegXk4SWCBPiGFGACqHlwV2JMMP/s1XyQUArCttxPibrdRDdGsR8BjKtOa4b
vwFi1JYqBpaw/KM42be8FClJ8kdRSkXT3bjhXd3GrwxoGt3eTYHN+Bao+VWW
JTBddIdhDCi4N0M3Hsg97Qx1/tsXY4Iay6em+iieRgb1WKfMRJ8rAQEIhbfO
IyuECenDqG5wVPXFCNVZM9FFC/fXxD8XXKSBKlDpWQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cZeGogiY726uFlcuvmMg6NBlbxNrXknm1YKXrFd3oCrxZZMr2BkrnbabRVof
t2x1xQ2o6tUPeeDaMomZ9A1Lcu0ORBGtTLkcFj0sUTG+ABGQgAQ6nUW74MnS
UVs3h+P6JFowhTxeTiBIsFba0U42QeGTaM33WbPdLgZiO4jW8R8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rJOsaxOoV5xIqt6BESLU4tI4IsW0L3xwvQ0FmDrY6RO0tuBHt4CPS9+Ld4ZW
k0RtVTQyPtMtORcEp3hAeQEPsDnlIU1Iihmj3XoBOBRq1HCNzsIe5OC+7WzM
PM7pnE4PCF0lbnghd2bo5WA0ZhZEmGTXMWD/JVSUxo4gf38OF9FMrq3jNLgQ
VPKdc3pxKpY/JL/xuGYGTZ1d47SNMCNoQ5XiMN6OLkTtPFWMhKw0XhoaybjZ
2u5EwQe3yuOo65iJ9o/r8aHEfxRO32enk+Yk1/aDyPE1dIJuCh/36geRmmHn
/2vrJcL1QEjluU91yVQeV02JJtSfqOBjBfspD1CjjBGy9C6HyHGm3iWH35IM
braWHtLCMXQId/jS+YsRCDbe9owExuAlM0OUiBlvUtgGzLSfn/+HkIdHlg6v
2iFTUrtGmGhcXDE+CUxRM9YW70ATanC16AZz4prpRBxJz3qWXQSsU80Aze1G
5klXA2DlQ/q0senyh8kjmvnWC6TCdNH1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jGI14j7vmDr2/jivGQ1rCONXgsIt5Shdem5v0JaoNXKbElc2capZ/TmgG9QY
4yVePphPmGQsq758UxAOUELZuHUsMRGRfAdOUAiFQOgRJnvJEFOOYxxt4mVI
WyOf0rzuYXHbtVZO4twdcyLC6Rgghs9Xys7ctWg5aiceY1irwdg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Gimix7uzj8fZ4G/h761f2zmzAMbmnrdMwHw9nxRiZwkDOyVxuTqTqlMWw0Gy
E/eGQjgdzS3V1fyJkIijKLYxzw2iwOudP7XVhxkaqmuj2u3fv2XLlNagj6hX
PbaYTHv+ZPkQFlIPfiMDin8ZR99UiXjcD2AvRAqGTgwPc4BRJ94=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3264)
`pragma protect data_block
m26qknWgn2q3zwMn/RcmHb+Ca4nzmp5CLVM+xhgbr8YgXcZ6QFEbnvu3HvdG
PLeIPNxdfVsKHTHJhkm+wmfNVVAAkvis5RY2fLiCcB1euEvfvE5HyP1sziYa
pl+/8GezgCH1tQ7K0sX+r5x0Ax0jxlC0MvpoRgAckN8HQ2Ix4H3TJoQx6L6d
oRzP2ngqHnv46x4DIBk2/6bRg3YoC03hhaVbtJFjW8dSaRoss67Rg7YHiFiP
XZ7QDkUxoWn8E+g9oU2ify4mJwhEsEVo9HiZFmMmBBD1y22kiXM5cL+J0uQN
cSwzyNX1y7Z93JkdkpwmaCi8DOfQsl79nkxfh714KJZ5c1OZNyDaj0P20NYj
QsR61vZjeg05WOnoPR6kSFpeb2JopUy8ZnXIlIhI0x+a2tRZhMG2IaxYl0aw
BaQbWB3EbgZCjpBAjqbaF2kaoL82fC5LzxVXUOBi6PUbWqXwFxMigXed6cwL
rgENIP6JELx/WKFj3GSGzNUm09xZqn5aYCvYOuwFloOYWc43KvL+Oqyx2EvM
ogTqzkyhwit3VxBnBBuydQDeQMdekGfxaCPTGDxTYaq/rNLHTralEqAOxSqr
64/K1SZUflBpL8muzp5D9vgyFMDktOJUu4HOuubIXGaeX9P4kcKVZKFwvDU1
j/gsnhrzYQWkkr8X5cogNv2z+l3EG+yQ8kZgWmC0KePAfwxkrv4Jd9514wiW
fc6VIQgEKm4vgNFEQ11DANMM1Eukq5X/gzHSxYy7Isy6YocJnkYtCqd+mgRo
FxEa+Vlw5iZpSSBA5buER5znu8vaPjLlLZsV8Vox06qpo/SAxGRwxkxHtGxg
m5dGSONIEvaCYCpNdDMHY1IoYCV1Y6tYlctnSQFy0nQk0QBrH7O77lYV4WyY
zcaLqIndMtPCd0Io0nGSYq37kCnxcoQ5+VlgCXDVrbZYZ+J0ITyXAxzYdOuQ
+5ocXJleDSu83E+bbnK88POekDYYU9izjRZNDXGl9eMIfbA+jvf5z6DSPVZo
/TSnm2zeNlD7rBd/sCF73jpknD7eINiF+N66SvgIyAxpYgSm8Iz5LFX1/KGw
A8VGBhCisPf3YmeC25WGfzr0SudqctHTWh9cO0oxAdn31Jk6De5Ye1f4EU2G
emiCwNeeveXaxzb7b38ST3dJXzs9KsH6HbSnpx2uI5PQZl7I7ic+GHsB1YEW
UtZROshL8Ka/CzFrf1+m9G+5fZdaD0gAg8WZv5z12/Ie/mZ3kwXn6HiCAJGg
O2ECqHxXe3y+GZavuw4s+Ijwkd3Alx0cZfc0pVE9f8PbhfsbiuqW/VGtShAy
lR74vtqgSVNhrXg0z+LrOfwWi142U3yDRdnngKHFKm0T6H1wM7hKCot/+Wbr
O8zEp7n+N6dA8omHWgiH03I7lGPczJ4MBXs13GX0nr0yf40vNkA4TelNXMaI
fLC6opD0MY390gIsdR5KXN0D1JDYYfQVM7LGs/gLsP8Zlh5U2mQlr03IFDu2
8Bt6mhsK++G1VQXugBTVNRpMYq7QbWleiZBQkyx/JyNIthRiqXPKwg9Vm35k
VxsmsWzKnzIl7bsRd1MPagRF0bNR7AHq1kNM7ZCvc+N4rEdqJqLppY1avL4c
EQCATQxlA+tvT4IhRc6+5GNDZnmMT54HcrbD42OctENHsapZuZgOigRLJLIQ
x24LYFsK5tnrhDGLa0H1XPXMYiGU/APs072xpi3uRPqg7iuhvqo0l1ifc5Qy
hpKiEtR7Xc5gGl7OgoDFtkHg/idXh7wXieDXS3J1Fh69q3mL+3ulVa8hrjtu
46vx5sY5SOEBVzJIDDVJlT54j522i9+yz+e3hjLAoDOES3EdpwYF8st/vRCk
ruWdEAawXdzmcTaqaTWJOvWNw+WzLj0BDRkaf9yCQO07rzY+OzGKYj4pt8Bt
Ib6e5TZus1rJxp355Abw20zn8ucVZ195rxvmKAOJLsmo/AtE45DmAwEFGm9c
qvV6pbCqi1VYGYu/mHKgHiVBag1qeMBRXfb+INLdUoGPkXZNHQA0PSu6ukRB
SNe2SOR8FQpYof4GMCkDKPqpHjX4n1qiPY6Y23vZOq506Q5UM758OvgjB7hO
Y3IHdom7luC1lbQEE+ieNRL66LjQcvkUPe/kgi/cN7jml84VlSrMyKfBj3fP
NM0aYMEg83Hk0qXtbTt4G4x9uF9ptoR441D/kQddtVu3Q5eaoMv6WqJ8yTvZ
RO/PIOOT4aZa3KiH+PhRx/xnDf7n0OJFmQtZxtWhH/z6KmsDwymEMdQNJIhg
dTadMOjdmOioxNqWdwDGMBAzzoO/4Uz71zA1aMdTmjjbCfyBuPwWGeWJeOsW
/zy4tMUS+U7Vr7iEFxSRq5gA2khHZK2hKnIaUHR665gLCNKYRYK3JEU5bKO7
JbX/Zha3CGTWX7iUxM03iObs2ittS/V4Af2hsCn5L7cAccBT9bbtUPJdYVUR
iZrNJsCQtL7u6nTFlGBECbjF0DfWIcSO2s4xcAVL8cbk4SmZ3xl1wHVc3ktq
aaa0PKNquY9uzq0FXIHjwcxWS6S0L3CvqZkQe4nVn4GVaoXLVDHfM/OEiqGs
aoJKS+BpjRHWVPt1lGSd59Nh62/m2GEGvgPzEixA3o/b+wFhvWLtB+41c7RX
Q7hWAH77P+fJ+MFkmRvw/1EMbB4Hcq2PdFJ15vMiQ2VbF2ytABCxfuwHRDtk
DjZY7JKg+ZyGiNR7ZJJ/HppRia3YYwXRNH9GtnmdlNFVSACHgMpvxHBlpzKa
Jfg6FVI5hFSXVJEbLUMvi5DEUh6g2EUy0xR9+S0DcJ2TY4gw4vjjyGguCrZ2
eMzWt5Q5TXFRHE5o0OFFjsQupqhkvlPHHSv/GiteowkxUmgNUIYcGYZ0vmlw
FhDXJQRhee7S3uQmwg75YvvmtFhvWqpFfGH7vLOTBVvPg3oIXWLkl9ys39hN
n+QFS3ZQfjPawQ4UP+Tvpuz7NVT3z2QoyE7+R/6vx4UEJEZ8cLg49m5AtOoX
KA4eMyz7tWfY+lgJuLZcDC7kdpaVOsei1kC/s+eldd9MGal9BLfno4tx3/5b
E5Q/0q9vQjyLD2uSOWzy/43iauFFhh21D0TKHUl0RdVRsndRW5rK91zwV0Ls
yYFBwAgRo65htpj2qpOO34V2DyXABXJjinuRK8k3n715+GgQjbL6NPqc6+Mk
qOGFaeALoEfkSLmuYvpU1ROHS8JWx+A6nt6tYsHRsGjk+7Rc+IyePhLj+pPs
N6S/zUjr3VbFxDoCviGvR5JxQS8Rqh8W9dayEB0WrF6tszcYAeb0+X7M3YbM
Mb66l+5wjkmHBNziLLKvxFPG5IjoYjlO79E6WOXzQT6n+t/AUhFaOiA5Fgv0
jYwVW3pQ4h7MDYBQAIYq8xjDalC4579pIq7ZtphFPJ+85+ofpe8R9SzY7lrd
aLAlahPXbyQzHNQoFVJstK415cuUjdyDDXu369DzyNIHGLtz8ZU1mYIIaG56
lEtZZh6xVBM1LpWQCPXP5s6TIAjUFPAtM08ksLBfOESmuP70YzCJFVosZsY5
sT4ozH5hQq476TI/NX0w3IdRIy0HsSZTgaaG/50Hg8K1gAZb6NMb431ovG8I
GVz1dVCuTabAfF1/BWUDUsogFcE3B2h3H+h1cNE9wZN33zmDTvGfGL57Nkwz
ZTGXxbB8UuqTiT2CV3Y2N9p9rbHnkeLIAgYGWxNqJ8Q8gPuzJ/ZqqOa9cU8u
MkPvwZEyWmlrpsRuLyrY+Iw6QLTJxtY4aqMQM+piYb+NmMMzogLO0Y7Gfdz8
HYsVPjYbOWKVTWbn7ZACF1e8McmqS+arHUn8k6+HyvtGV1oiT0mK1EqPBZ+A
9DqR4smjScl5zxQAxvz41Qa56CWo59YdT0Fr8e8zsjj6pkq2xaWisyEvE+ja
gZaVokdSdVpGD/MreBJdvobD1e/PPd2grtHZFWdlNS5qmV7T+I01ITvyt/4w
TjC01t9TqfH0f504nXsaqj+jMfU37E2XdqQ6AwaxPrDBcx4RRlYo+DUjAbPK
rkwpQH54/es1Yqj/+fYIg57tM4JFEVsKrcVCeq3+Ic+B88zhWLTKpZDWB8/e
TkAQiqLSNUtdRfLc+Cu4+A27dUoS742ejh9QQ5xUvE0AS59LdnwPDnCwKFi6
uqfYzCX8vbrB2DZ2EHKmI019kY7Bk8exmP1v5uapmY4tlmkBV88b9/Z6wFt4
N9vQ+vDXlhj7lBtEw38dZ5GXXOf2QTDZVYfmBReuy2Qtrq7SjV8EnL4wMuv8
l8bDBWdo7aFQ+0Qe6TWDj9eGWOMQULL8E0U7SS7e9ZxMqiAyKWJvhXyuoYzi
bhqZcQnLWlVFA0Qc5TK6ZC5FYe51nMVJ

`pragma protect end_protected
