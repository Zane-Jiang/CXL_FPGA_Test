// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qcVN+EpYyrlGppUwwmPEXNS4Z8Ai+muD0Qw9C93RzTfTxoFaNBD1PBA5DcfPfYoIK1QFEHfSNZGw
w6f1KrCvTtZ4PR8AzXTdgqWYmMmYBuD6f11yVSw7bmVe8+G9Qi7PHTxT8m2tjWMTl79eTljyPuq2
hlAYMzcnEdK/cVm/WzFP/VTpio7SAMT+Y/f/BGyx8RCnVGxkAvfXHOcuzWVPnWppxXI6GRgBDdGB
x3pHOxrChu+h68zN59TXXTHhAcbsfb0WtgABACMqfy48ukgC373dH/SA3rYrK6IeT4d9vFVyVJK0
4GPNZyE9w4TwVz8AlAcPedShFTe6HfVd2m8qsw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1152)
c05QcFXGY5UXnULN+OzIZzZQG9/WZzNrN5bvU21IzPThaFg8NHhm++UyVAmOKP02qmnFtrr9jn7a
IPxVpWa/GDtK3uHOVZrDF5ht5OzSU4Rxab7YJxBg72tUX9qCIYZHR6W2agtd+akRsuaTa18aKXrT
euKWAdRfknmb6FWhBeq8Etk+QUMrVtLUrFx2bEMWupHZCxu7xpmQ0J8CP1mbn7pzGKP1MTw9pvZl
mjGKe7YrPHa7XY3NJ3meEVz/PBIfELBaNlO8q3T9vScC40dLbUdaxYaQC6rWazb4DTaGTPebw8yh
bag+7vkMNXedvtitr9vbF3XQCLeHC3zT7spq2eYdvPHEqeLkla+Hm0dc5XjvQ1o2MvwI+5tt6+/M
ZZ/hr/Gnpdjzz1SYWhyx/xqGDjX3RVv8YE6z2WdYvQ6GHMDiR0c4hypiI2pJup1E9KMTDrWof6qo
Hy0YrlUCUdJXshcpkg0J7KaxKdAShQDEIwrF8jC/Z6MiwhS1PmbNykdvp63wh0Pc1EHHdcwx8jO1
tjdQO9dbQMhAgFqejwEZ4yzfLCAE48GdWyOOTcT97ZktfzxDbNj0CEjIjQaWPct8YaTOCwYoD8pc
r4DIBkf+iBgvOGw34nd4rQB7V0I95Z4DnF94kPYbNHCKf9HByyCnNlDTjMOhAxt5NK4bvAjqjFW0
iafnLRzMEzkoMfRW1gWf6U5oUTYRyH5RnZCyFPVqf5NIWD9YbqusOtqvkxEqMaxenZvt4UFMdZ9c
3mJND33isUTCSczmUtTlNBdHr6HpKk0rIdawaFgccUP7MgwsP+XuW/Ndcw+HIqrmExjBBdT1y1mo
9tRNAQIXa3fczXdq74pz2lHUXVV03qbAYaO5YcD+5aJ4t1L5QJmFtrfW7JgRY5qMUElCL+JvR7Uc
pCrgipNZkz+1T/4u6EyJfZNRAADjqa0nTEzi1wdzOT+TYviLkT1ilrAyrzhe+kpbHblHugJt2M/j
rjWIxKSf7ejvY/swtVE33+XeJv+tepCcU61wpgm4rTjO9mLu+LuB3FsWJllHopzzZkYQJCns/Rlj
f3HfLVxWkTkBplf8L8RWB+xSFkDmeB4WUh0lb38xHtOILmWp2eOie9qSjzCloQmesc4RN5ozO2UX
ZtL5MXkn2W6cc5iPpVKhtgcJGw8t7/rgD1lgqYXYSggMEOkEimm96/4+A0/eyQ/xGByHKN0kzTFv
9kACher08El6e5pXYFbb2wIjvqnZ/IumzESiIgVMklHjWhaq5MMBM5emwz/8zSgnds0ENnuUHhps
yA6oZA9cco8/8r8e3VZN1v0zfmPwM7nI/LWSPUVQXHbY7ttoyUhlHaqQrzLMexj5rzm9rUnNrvZ0
ACgwuTu0dAQ6DSV5u25vofMXz4ZMyUa/pkkoBAXyr6l8R+ryPXmKS9xUVdJSETiIhhRPAPvWE9RN
/7B1YGi1lQvzKAGJJsAVLlUyS+D+Rto7DEYn6zDLIqnJeU8F4+K61GRFFy/xbcBpmUAUYOepVYQw
TaX+Q0rUw2Z5vw/Z
`pragma protect end_protected
