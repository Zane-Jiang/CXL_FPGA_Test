// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
yueeaHa8ZS5mCpBH1wAs8XipdGS1AGrLmLzB6eciHvo7ZVodLGTHX10D2gHsof3acweZiZG7Lu7R
QkX/kPYChXwd2i1FFkeB5D7ECRKydPo2Ie5w+vPHBwg6h7lV8A5b47CMcVmgP7iArFItEwWDlRcL
6tHG5eR36PH/625lcp6zkwgBFuj18g+jCLISDZhE+WQLZS02fzFb1LAqnr7srUNSsHHSiAUjoXM1
V9Z9iv7r/THxkjpBLpqTcY9AcfqqwiVdE60HYOm8iC/ZoDCXI3jhRkesw/OYXV00zKbrOFb3ww+9
/PcUznH5kgBaAgrYGOL0S6QAUVtUrbK4svPqRQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10512)
5dwpe/4LOW378pa3XeIdOhFvS7j0cVYlnN/HSS8utf8z8FJbcNE9B5u7M9gQrMtvaH9Z0bfrA0ZO
DFV+tdvSpAKyQhRRM0ksnMZ3nh4pSq1GtPRjhnA6gz731LI1Pq07u+XiJJnX5ivXOEneiVLf9Xpg
82/vhq7fyJw7x03fddYVXCspmXUe5yvzePWnR5thRPKZBP3Jc7Cf1+OOJ0BG+JRTtKtahtBPImw7
3hcoN+azpR6KXNTtruLguuPStxwxSrt8aUBoREWl6I4Pu0uBI9/uBXsfXDedW6lbyHX9pSTskD7N
rscLnqK3bcwzSEN6iW0wijeBv22mpKD0gkRfz5/HDeXubuCwMNnEhldases1DkncnyCz1Vmba9XR
/0UA/DneM0h5U/j4XkLxfTo2qzIVz/ydpnBethFPzJVgGAiC/MaWsNg7Y2ISdXeHyqD7Dha73+dj
DGZCMNLVvUQHqCABjKklJjo1Vb6H1W/XDGOV3lplqpZAAj1bDAoFkLC0MKrYffG7KmmX9nttMiv4
H+3ByBJyKj7xrZPBGZMmlvgZZ+thJc59PCDNQwfU5H+D9nMi1ot6JUMQFcJUr2kg9WlQhpy4lABW
yPI2GwQ395SVW+YXly9fluXkwZr1pWcdA+nDNpFnZMkCNZvMNKaTyEvS8aMs9JKhB9vTPyu9oBEI
XJGDDwcHFJynWYfbPvfYCDglPn0U995vzXl+mp6v9qCWWp//tsFrI/ymfRAjCm6r+9XSlGoyY+9R
dpaRibMgZkj0TQRLoR+hM2U7dBlNR2cOq++RJ8M7r8GxD+60CN7ucil21kSBHgcJOFGzEJx/zt8E
a+dZU8hVKqGJPFXm18MUWHTVFVMkxN9m6X9DJX6qxivlfTjkmALmuZwFx1m36cacZDQlqwzx+UT2
t1oVpxQSOxb7XK4MqhJ/lZA10cebsRb/6Ww6zch1vJGrgT2MXwXeOUHnXhg2cVJ829j16gZKbNB3
h2oundT2hDGpNFFqP6mYqk13Li5gcJIpfuyAHjdPaAuRGtZhVZRlGH20yzcJMypmgUuaOcA868dg
j2Fu6y4R0z64qR837NjRSc+inSZDYR628Z0Hm9s1kAWnXq2gn0eF76EpkgNWOKrw3uzvfA5GtYlm
66xYWbenDYtWSlZ6v41A8zSNPFadFXRyuu/GC2Eo4moRg+gMOhkoPmE7fx/bMem5opUy/sjvXqzE
Q7FMaGuGUY1dURpPRPFrpHMzt3hkihpaf3Vk9vCVbBg8IwCpWev9yEJEbrE/ZXjAVmRlP+FxrdYt
EO4dfM1SlW7gi8nEFRbkqTY+AS282OqfcXAQjDMO/j9qz8hkR+JgN/9gO+oTCd0/ZSlwCdZMR6di
Dvwrh5N1vKMjpBx/y9mVLiWMhWNvPTWB3v1SGyBKZfb81w2pEuTlDw6EBu0jkd1SSKlyX0EHsjtg
uxtNcA52O/Rud5SYyXZdmIfT9uGX3lXaicvd7KSc3FofhIMTjBcGT2sP5UpVnItbv0bh1JY0uMsw
3dJM43YtPQjdhI6fcXOA/tGnLr7EyEJxVs1D6qPq902OSXL6XSFp155LbyEAYPH0R1sIRxZ+1p+a
IldnGrZ1pUXBbcNALkvbKCKiDlzs06LeeK3ZqSV2SOdnNjd8D2jZu6UcuLwYD9gKkX85mPCG9TVj
mTWq1R2yzi4/M3hHvmHDKkg9qXYuK8be8bUyV3HooiUrdGhGEaR7SyE11NVBlUAa47IJi9D66oEp
ZyF6VtQsaetG3WUvjwu4CdOhEryxdEV3+82RQk1BzwwgndOsArUa0VFaYk+p588gfsdS71Fr0XIS
Bwj/mVUS2srX7LetuLnZs1feAbgL4Wu50z00l7YOrHxJ9RkHBSmo9CTi5e357LEz373zVLiBYsV4
rS0VyZW83NGnguna3ZcLTx4YXQoNM8Y7kmzgDBMKpWO7bxXGG+mheDGQMJri+0kACTXaX+0M5vh5
41VccFqT/kbfnGHE8+lDq9SOt52lGDi7+DljvYxXGnoHa3L6vQlj1aKJ0hqUUWYuKNY355R4g8zz
B8Mc2haidpOqk7UYOnDYVARYrv7UBKwDSUSAfO2lz3FUlsWz5pN8y7AtQ/mA6JAlP31OpOd7rSf2
fu0DIvdQZeW+Ilc3Mjx7mts5BtNvDVE4+aCkAkYv9xFISZyO6kw4GCCNVqi9uEvn/GqjcRXMzi4f
ae3l5HYzQ3rR5cB9rqZppDkkabTqGiUzkjgQt1Ce8MwMdJjEsCJEEXiBZX7PCpu0ClBl1mIggX9s
ARRWttt7th4MDCWMP5+EU0XMqSGTsfxIpw8VRgDhPoOaOSl2i1Vbt1HbPuUZL6UyhaC4UEuBajUt
UEN8NBzbgXaPqeZw/iVdXsZV3Abh1Oruh16oPmbcCdy7PbeyijL2DuRmHokxWEibbwJfD86tTEzi
lEk6RDCDaH7TGHoPA2aAeXNJaSl8DbGYyM0bbY8Rk8D5gGfXM5GZvseDUXDq/fznRGM6qehF+M4w
XllkZpgZAFRnIYWVW4oNyYOqcWLjTl6F9ukdpnJuF+ogLWqpBgkADHZSNiwhu7xjHn0WvimG6qPw
PXP8SJ0Rq2hc9Jdej3BAhFkX0qpDB63GHMQV1eXEHZwOBv4lQ47bgeL4upiVkGq5Ry2C6SkZN1y8
NWV8HkZx+Du02MEBvMFz8XveXpS8QpayHRkdL4JH9x+6Zo6NsFDyttS8JT/cC/sDZiD+UBB6g/jc
uHbEHOEUjLrs0t7ITQgLd/spF+6K95SfhcS3C9jMrj51B4x1CopQHNMaAJ4pI7h2Th/hI1cAEFf1
0zlBk2eETVuNg3i4LnPgkwXV27D7JNf46u1f6PbkI5YGkn/Hm/KIqAVR+4l8lMnbyoFYY4oVY6Xl
OGAN7vl6y+OVIPi8lE3vHqDqraK2ywH7ihsYska35qbP48XFLpJTLrPyDeAeNWiN1/b/+WwjWdKd
sy/Y/q0XKqG0f6vNmTTqLGzKPOxTEM98/d0QcoZ6vw9HMzOCEBg4jwpZKaUzPkvijnnib1n2ok8f
nrX+VDdAAgtKWbYrH6fHOHDTgaSYAzDd5YNmAAxdfKnPMvIor1FF8ooczl0WSRQlthBQ7DgXPJdV
TYJY1VpOIMWOfQ055MElz2XfmHv77YpNlO0USwM6TeWnMGwSu1mFM9ic911iZaXQnMu6KLHzzJTY
YOli3R/OhXxfZxE7tdOqTa0JWKxibMN8niFMih/nV+jEkHDMve7Cftr9ZpmGpqykHfHFCp/sUILA
+NkbZzzSyne51fo1jrqH4P4YyApFD+4Opft13SgsG7ObCgP3Vb+b3FhM7EukHIMiQyVd7/QP+tCP
/S3FBilJzQFrJZkVJFwSVBufrsqiCN9B9+cX3PXctsk3W+bbMDd9uS6JSWozk4G3F4mKOURhwKtq
w9YFxlZWrV0h1g2pGRg/ytvD8GgFaKpquAZvkQ2g2Pdz1Uv07NtDUNScYCSGAxRz78Oh04/w5jv5
Cg7oVfqvqlUxn4uRh3gRyniO4Er8BTTBAmnT4KRoAsFXpNfFhxvYapykQ1M2r674dBzAl9MkyDX/
ikUOliq8LVqMttbTYiz0pW5PadKm9Vml7Id3oPwWeX8+XGkteotJMNOOe6YnnCxrBqqnf/K2/A5X
2ZFVwy973tZhKCYhbnfU4SdasmM+I5p3lSLtnN5XxCY4GrSzJn9qD1doFYz46G/xqFpOduQp5QDo
dcqaLTMJ5L9K0Bo4kzrvCk9dQe+iGPg+ASu3wBye0xTrAxcyLLaFXbzXseOubhHfavoyTmzDUSko
5g64mDelCHunUjoFENutPgxwD4EoCRCCOXs4gXJKpGgrFhA6CScS6iJ/B49Xuri2FDCRAVuATYtr
6kh3w3NHdDGk+CasWsyOd+NjBPD9Iai4UkTfMn2JofxQ2EFOLFBNHrTNYsc/eRToZCRv6qQYqvIV
InJFE/Zes+vaxqFgBedqtzjjSsoy34tpN7w8nAuPumEINAE7bVn/UjG2AOQ0uvRF/iNJIDt3vZod
8O34Bf9JCvu1GqXm3mPFkVxs462/hLZRMQxFwhAUNZBU1sPfjCvOWn1KOdvFK4f1qrMov5VxQ8Wv
M5BrQ+zyJECGMjkCncnUCfS3tubzQlV6zYdpupXlTA16K28YZST6j7wLqsH18qYxBJlUMs9fDOPs
LjiQSCkRph9bm0SbGYdAsZn2FtG0MMkSUb3qyvStmyPjwlYRd5XjiA8aIcoXr8wQiA23RkGlcAhw
TJE62x84RmZ3dhT93y9fJ6ACNLxXenPj+SJdNCEVDk3swuHwrWWbPKimLEKN6XpnHdj0GNufb3ey
13HyrITfJmXRyqm04lFyymOe6xC970pnFt/OjLvK6N9eBrQH+kK3y0GyawfxLApU0+3w9C1rFgz/
hS8qm3HCzYbXkw0E8QZ5F8sGItdLA/5kJZHcdGJCmYMz+EB2spEzsk96FvBnyyeAx2kRVug2dnBW
whcDJaw2m5LZwOnOafUBxVyPnR3l7iFRddDes+DdEOL+w2xOAwEBiRWB3HL5I10NcVUOdd8DPlEd
tOhG/e1TziAgSOorlW4FMhOJvTrvOIVUrQieDOyP55ZSizY+YllgjQOxmWK3A/50rdmfqyXxaeQ9
Jr5BRwNTua2/JnHm/KP6jvZcTx6bPvnVIUHOCyfKMRzmeCKL3/vWvmWKBC3iitlN/INW+tJnAhdo
WzDWveYG2L5f3aYkMYZGOA+VbF/gnNTyoC1XZRSMMhrD3V1X4N5HWSy8xTPN/MkEObooxpdch8QC
D2lcDBNSvdrIrzLhep1sBJcZ37FJL1RWMwGUVX5Xf2Nxjyh8e3Sh+jOsYsSlNRbVMfHMllVFMICS
qmc5sMQSBxL07n/vltu2n8pHYnvKApJvTbwpBGBPHwKTpxzTWq6RXSw4h680EP9v48kh8+6ie+GH
sd4Ww5N6l+IFLXwI4KZza227grR623hlOVn7PRz/S94MSbOTAIEoTLadBdBX6HFyoSUN428qbebk
IsIWGZT8jhTTJZ492WTsVjn2MeP43BAnSdXrGBmH4d+8pHZ3KF+FGpMEVBUjn2618o/IxoeOEFHr
qPzv1Q31MktFrtEMIdvhFu0n/B3mUMyKBhrjV+KeQaHfDde+Giw0nrkeGtu1F8GmYFqtq0x2FWe1
Nw9fPS7/1ELwZT1sZs5weMpdmhkVFdBGH/5D5nOzHkqTyFKmBa95Wq805dFB/IrlblCHyYbZJNpt
Z2OVg9wykAY3kvQUfq1C7/tSTYUjDBUWZVtRwF0B/uMSWRWPHijIoYwYy3TPEyZb6bZ4Rn5Umbgq
1UCKnilC3U2LeMVQUZRjxEaGbsAVXx9lPr0BrK7gh48BmDlkfxNPxpv+tjq3NQUyaplTEC0XksVW
3zuwQspy26Z7n69TBdZIN4voaKFm86LR2FFCHrTPpEwNDPgEnXTnTBvN4GjUjvqD2KJ4bgHtOYkj
kX1OheCLrx+4mLbqEnxv5CcXZt2eRdNPO1ew8KKqazJbtgPgzRlDNyTFykljDivIBGivPfTvAfFD
MGdxsAkiOkwrjSiVRAgZvNOl9hC6lA/qfk7wZpKUBzn67KWhQFnw8MAxHpLJkw1XGsrmJhZBh4ge
DG9rhj4B+zCj4PBc+tj9zEIlo4ceDrNnITaan8ybSUK/KfJP+U96PdR3S2Ut0dvX2LXuHDtlmyU/
A1ha+xwGnu/ncTb18BiZRPpM+EG1ob+FA4QjIydEbh4QXH0fiqd+KQ5086Y897MUOu5gl5Ugl7tj
Fj62hClKxFC+hvo5913+KXv4iemvcj04L0w8jT0c99WW+F/mx3rF/XQ5qQre4k898KpG9rR5H2fV
JQZo4duUQwnBcNK5sTJjOjLp/NLBjkK32FDIm8uIC+hrUoreFpK5m56+iYk43c/wBjx9V5wComDA
SPO0l8bMQiAK2aXwypZHEc6mj1GUQyril0aVxoOw4xSAKphUbiXIImQ97DXXCjcB8bFSU0nB8fjF
XzRAt+qo7dHoulgLfyWdDrzobj4yWOwEWTT79b/0Gvd7ByzK5UEJm/52i/OIhg9MryLxbZGZUwIB
BklxLiMj1pmDnYXhNf8Jk9LZscI1Pfo06oXKR0qL4iMiyKMJtO3iHtR8c4n2PNUNU7q+gJZDefYh
ScyAUQuD3DaZ+9JU6h9w6CzM0m7BL5oH4ocA2BsCklJSxGMKxFUK27WbJ5RPlLS6v0ggPndfSO0M
tQV91W2TN2FJ9z2KmbYzr4Gov5/fvLTr1JhdAFSFxQDmblz2o8JZLPTCE5YYRIk08gHoAh20btmE
WveJM1HXmyg1OkqgXrm3lFvEC0X/7NsxTFiO2ChEy0m4i2u/wlcaO3NYyuQdbTjO6WJZMV+bXI64
8cS2RPRdtAldEBVR+RtVmLuDkQJXIv70E4sn+0l7jBr2u+5cP8VmMsbBi5Z1SFbPtMBW+ITrdg+n
3JeqoHIO9M36RrzV4U9HPJhup9Uoj5NtXmTehn9WSs1tvMDlowvPcWXD5BrjJrdva8DRqhssaZtc
/jVOaPWWA7c8DE5ESFSePtAe8ogCrFOYf4OCR7i4gnTzh55UkVCrVeZNFfzE3BC2OBG2bR1T0/zn
I0MBjOvRUqZJ2QSEF6KyWAoWYYusZpkqQ6wllYl/Y6WnYJB5RhfJH7di4+aYJM1C1/8YKBDcxXzz
sPVfjcp2HcEQGowajVweM9Lun3fNFhzdiVQE0o9eCLwgmy59u29GNGWuaHC+fd65+vUrju8SeDOI
3SazWGpMr1+jlILVvtLAgFmX6idRbvpPePquXioZvRHoeLemIYcOF0EtMs1p+Znraw38G38KpYaL
MhMCzsQribDipyIR2qua1qfuMGln9/VDI5CIguVsY2DwwN0L+PeParmimyKhKpPNTXgkUqwh3+5K
22Tc1TbD5tOAVxkYpFuCWkiTAo4/nVKaaF75/VO0Fw9kTNH/jMW6bqtUVM/In6wRNWN2GCY7Svh+
JhcvB2FNddQ26sZqTi1OrB2PU4dSdrAjxIJ6VCHax5IyE7DUInU7/J2XijVj9E7KF3ZEtiK89J2n
BZPUXgfwVasxdOEftbIJ+ctfixZk/izBN3mPxl6e3hb2coMd/a6IWuJ5N1NOzqpkIk/n9iQGfnGS
ADuE2nmFTmRkq3qGEPXxc5VqmyhIny1aDv5aVkIc/eDpMkRLUw9/gycvxlcG716xjhlDQ/DAs3mU
8Uu2uwASx0395/aAgxf7VWM9/X8HrtOV+iagd+f5bXY3RooO7OI0QIyV8pRM4LzKsbgYmZJ4IyZ6
OYQlZ4c1m0j+qkvQGziVXdEcO+x0y6aE683AwhZuIXRUrxC6tnAeKpOcXZX0SnJS76rPGkc2JSMM
u6juQhBzdVdRv45gmZM9ycpy0/+Q7ZaX2TqYAallQ5Wr2KWwklAMkzkkBWniCqR/UjRxxsFufv5h
Y8BYv33wZyMHnrhMwX2G76Up+QNslz8Q1l2TY2Q0TUsrsLgkd3wn9GAa8euvFw4SS/++kDLOH3rY
ckbsdFIawz7dhB0HQGZGaezsQr+qADznsHbRb6plNE3IGFLSr1M06Zn9bxDBP7zyzVC41x6ijgoA
Lz9hXoQKb8M8Es3vDy2kcWNYBxLnr2tsjzjQ1zx8AHC2QPGs43vSDW6OIdD7rAxu+olnnX1EVug4
y95nY87N22anBEQW11qvKMjmD0CFXNJPEUYUYO8uSMeCZuE3CgSSn7HX/zS4Sj3be0g/y/DTAWWz
tj7lEOF6G1/AJhrd6bRJTlqdMjf7oPrBb/KIFt7IUihu1P1lUQTWk6zilInfpyn4vw9HAKKsP0vL
FDSBU+XH9pXfX4psF+tVkOC2vP9qQUieYfr3hLRbvFVAVaKTxkoKr2bbjs7HXplo/NhsM+Sk6Y/H
858bPcp61mwkrluKu0ZPNR/PGoELwqbR1PMIb7LEOqtOw610mH7EJt/6ODTNNdpp1MyvMiQiGvTw
EfRjMLBm1+TVW5+mHdSezLDaSUM5XCpUKcmIg0qoU/1JnoG4RWTSg0qkB+elMAeLjUXcIot5qCDJ
9EGihqwbD1k5WErEVKfLB33yPALfJLFK7OT8SX/tMVP3kD7tHGOlEIcCYIKiBg4AAr/jU2vBIbfG
SA3Gbm9JDMfafIQw3ZY2UZazyUHOl+xCk3SpF+341pkxM4lqczlEQNcGFrltdYMk2+HBjwo6E7cC
BdHO5wfxoPWFCQgKbo2I+LUnsrjMsGpslbITwHKS7YuT9cpgpn4rUx6E7ghO7p7oGgujSMIrUTSe
oH2K+usQ0yJFiOJPmovC4RyAmmg9Ili+vOYuQrjVEElsZZCFAyITbgwznT1FqzgYQdZc9cu2+3dp
1pI/Q9vJanJyNcH20lro0UXweCMlwDnnm/Dbe539hlWu0RDml9KcMPBf25UUikIG0V8gbyWAU5yc
L9IIVx83wkq5BjSYmEks1cnQGC3rw97DgEX6lWlL257GTKUSXo1YU+w6ye21akUX8w8inVgXRrlx
AW8MlVL+vhF4OA+TrIo4s8El6kKgIewcDYNFequ/4P5OjRqS+D0fgBPYtAh2rb67xHz3abqeXjFX
fn++EdSxaYX3zC8DEAPVsCNkeTDZLjmdhuYeLMt0mKZ+OT0Y/fawjnDZFVVNzzemQtSNWdqTtF+z
cp+43uVbdhiQ76bbviinZJtMD3er8Qy/Yzn6Zfh3L6X/ZO0bTGVFECgjt7dE6YZZwezqPqrI5Rbf
ICiJ5eUiZwESND1HICqk1xTJIhhWhomG/z+7qkq2rKkOVUnSlezow67T7Gejb2fFdDmeQFpIq64q
XaM4dMril1Tb/2F804Sih9ArFG9jB5shghFHuhT4Sc0YT6qmtGTl303K5hxxw1SADabHlwzDl2X9
zlVvGdgBRmM3hprdl1D5n9gaovaGed2GdpUbCFxtgIQIdzhv9MlVbz9Si3EbFTiJ5Tib1b+6xfat
a6mr9sMYWNNF73oeJTcgbdRt4SNcLoQxlgwOHvVIx7eOwc/GFZyzC2BN3Y6zIQddFWrqrSrqMVD6
Am5PZRgobDdB4sreZFTJaHvzSaOn4XoamkTlPGmZJw8eIVlQ3KrziZqfQYyykX8q4ECT+w0aW5Y5
0EQ6cYpmVmpwf97rfVp16SowshXos62gYHxoWT6W+lzdejuKwwAZgOz0d6mpqBFo9dzB0xZQx9nz
e51q65NXJDF2X4j6LSkuwYUGIWYO0zY2JrxIIHv/HFzjRaylF0km4RWXiZf2ngYiXUxOj1/0/eo0
5l/xw6CgkpugaNC32qpCyT8lQWzS0Ydz4sWMo2Jiqjb5xsQKBRspGDJQ+fJYE7xLtsXFnwLxC37O
MtGeuzEK0MfgHWs7rYOe03k1WxWt6XUKSicPFclIuuXYZKBxIVwzsB6R+rhL2wqs2pBLCSxMA9V2
kacXU7MvnbFfbeZY2fw5WDQHdE12V5eZBbuSaMK9AS/xctp2l6Oo3TZXfhDZru4Sq3hZ+2LLiibb
iNP7+xG8jKf5EYOBRBnOVpWwe/XcHs5KEsCzax8a1sNzzPAzF5kAhNtVw+Hu8jtP67EXayafvBgh
YOLV0cvpCY7Bkc7EwO2PfIbbtwoQ6P8BODI/Zw7JqrixMoyXN31YwgjoPfn9BaxujvJUdLq/MDSw
QtsH+BbY4SvG3S6oLWCx6RTUu0ipyOkYIzW8nx5kymsr6OFAsBjbQ7vcRsTSVsUOjdl4zRifQ5Jo
mpWpCXgVYKSnco1I0LG1MJPQQJioddABbhvole+prPZW1HQkz7LkhuYjxVILy6q8w5AmyMgOlo6R
cc3mGkR2oN2drj2JJSTi9DMZ3tc69+nSgqzXYIXDZHRSASJwEl2kE6VusoCNaMMgVJh9IMCqGyPy
7KMYbXQcFcz5+QKQmnX9o9xiWN3vvVJD2awxDHO9GSOpHPVSpjjO6DXGpXyxg+VR7McUCAgA4wD7
HhiOwAl/FVs+f+wSBG1heGI9edh1VfuCi53NjqmHPKSMOGTAZc2LHjwT6aLhhdvZ7AQzax8GVCM1
0ab7j0bauTQLRmiL+bP/zY6u2gdOE4IsXCgxkxF8JTluaY7KeMjMxC41rFqe4fLZuoh6dnIKrsin
r0uO9sDRqWddyiOjPXnvb1rL2DEby/oQ/oLGqpGuD3/K3i/l7sKybQA6lm5AIlRKLY582j54Y+g5
kz/DcT9mocSGwyYmYqNO8kp3buSql8ZXjgHc8IRYFm9RbNKCvd54ppW5Ggj3bd7DdguERbxMhNaU
nlZgDcJShIQmYTW5vqmdrVGB3XVKKRhC4BPJOOy+W2HlxStiTEvMsRicP5j8R4XNHZMvnA3bkz9v
Qs3G1P3Uwl+qFLef9E6087rxY07PkK2c3Md9h0vUX1Y6yeil8dKscov2AWQHQeqSzCtlgZk42atK
gP/EB6IH9fbkwt/qDc10ZeVL7xZFSvMYHhelCPYECw1jNfb7+yU97lNVnKWHu3/zw+wrHX1WhnTA
O0xinPIRqe5KqBaWwkRLJd+Vn15L5VCw22lZDuFnPsjJj1ZkCCPj/3UNbJCZZQp1OJcrG3CVMKa6
VG4gmUsGGR8V9z8jMyxSI45V23emNJ1moamGWfKeOHthrHTDOUjqwD0wFPToq6pbFwWDmPFkVatE
WAdlHrpGBKUQ406azLo79AD5OEgseBF3fB5+9UIf8LCarLExo+ycpfam0Hyxkw/gzLK/vYJnc9M5
yyIAlbj1EWbjhBgKlFwG7Vpgj4H+oZC5osZDBTIWwLbm8tT2Lth5+WiLHy+m289LA/g1TrcEWAA6
e+1/hJlWxZzcJKLH0vzzCoLu+0RLrjvloHU+/19OlWUd+mvcC8kIRsTZefYNCV2lIq4O0konlBQW
4mwuffF5l59s3xUzT2cqg2simXKX3LB8ImQDn8OwQtRXtKr/ZvTzX1kYbU+bHPTjuk22w08L2vD6
F6JtYxICOnuIBdif46jtRIN+CVwzhzU6UpnEzYxfaKa9ktmM4zyU0rarGMJv8NtrdqXpLU/6qXOu
+M6c+Vb5NbV8TE49c1kLpkXTtok0KA122CCR77ydYjU4KzycQ13yRQyIAG4R30t3PY/iEKZAj/t4
2lQgIM6JYGao7oNu2NoqWgA0lze2BOgpNoYlvccv9FWmJ2+6p8ASWhPjYgNhfnrHiENzWH6DbRWI
2dF7UZf+Mo3LKJtHd6FE7/CoahxTXZom2MhHCGo5mf5jCdQsOy2yzrqFyPa2FUcJFI5Tum8qfyzt
sZ119zWdyU16oeVQwDQxHXb4SGEDod5UCe2nEuMaPjnMUUfi7M4e0nCh201Iv79Q9HdHXQG8BLEV
SJK4Fw9TPvAEZ7hfbmxR26XFl8xMkzseHuVYmubAc+yah6WrQqQI+ZJRZW6iTgf9NeZYGm5BquKu
BMubtID1rqwBaMDnozfCwZF0EyCS4jW7lfJp4tje8t/kvzj6rv/iO9AiP3QFcmg23rnuSnyVg9AC
bVjeggF0EQRQo1N+pIKLMHPOpJBtXSLYTfKqxunxqG1pttHpcKMn2QiJVAugQZhP1SGGupndoiPG
J3OR7oTCn2yOpUYSKPnm57uCZ6cWBJHK+3eCCeh35zCvBWyttqlw6FL3LTfZtAn5Mdn3KKZZKyuE
jsgtUzwmT9Wh073FjA83ZCMT8OZJ+QiVQSZL6v8g6z0IhUcpNuc+YEdl2ZftJ3MNTOV3uYfEN9vZ
3orpU3WTuQ3+cjizGQVGJttG9kIjKsd9E9dq267AQpVZ1k2u+zdxvETrKVFwZm1lKnCKux8pK0Ml
LTIUXAZtyuFKE8ZiI9K4rr5NPcjcZ3drwG2syPBYjCb8iIObAphobHTt3tD6zrIjDtX2J4zahOqf
c3K9E6JknH2v2rvf4exG3d+tOFpwInngafyxhZLiguUlVgwGSPf98pguYLD9BDEVR5jm1xyvncoF
8qd96qGBtSb+qwEW1sq3z4HQ8K65aqBT6t+yeT+FWrGdI7wriHrRWkVBLfropF4PcCiuelUcWCVq
yMo3D8qnZRNGn73Hn3/Om9cfqqo/RkSWvjjB8odDEj+GD1Qt94uJhpuKZCdi8I5jb5Jk7Le8Uw5X
39calDPlo2uPqVvASS9Cw06Ia9lHlxFB6Y0+djX1R0mTREx8jZY8pjCi1cpTgeSmPp+l72jOuoDc
y2xXlYSBikE6QbNtJhiIO8X7njiUkHdSM5BerSyB2gWHclfJc2KfGxdPWQlzfD4JnjvfZmo9kFlK
/Lo1Uud/b+89T5pDtkgcKahSHbE53Tbtt1u92eivZ+RvxpvLlY/CjarksWVRq/vzhNe9TrzoW4e2
Ssp8JLmmw7mtdS1lF3HaKJ04TNghresfBcLDLDa8AB7GFKy5rQDHx5D+6JYqmCQeF9k37PDWcfNM
I1GBF+VaSjVqmpfhM2HCEp31Y9CNxGxDuDaoQBEHLdDlAGgbIGxS3ltTkJPVMrtkLCInUgTvKf1U
ciqDuGnAd432OOR716KBmAzePhkBqSzzevbYFEK/R/IIjfNRezrdX6K5JrOSEEPDob1UkAw2gm0s
H2Nosn+uvskqqa+805LTVMrBxIRCZb4ZFWjnlMJVEJK4exm7ZZZcONfYFALy+IStzb/YDYuf6CZI
Es+Zj+WjMPWYiecPzB4VXDbrfoKsEn8DiTGZkCfL26B2z9UlLuZog8rhjxsprivzONQh9MtZgkcw
YfN0hMqnRso65CYk0PnIZu+e4LW/8deydmeQqdct1LojcoHIc7X7PeMCT5VuTBkg4oxlOMZEU1H9
03xsPW3syQrzGKYE6B/ZybS6Zd3X/RD4kfHa57VAeDho1gIwGGYdpKHQa+Vb5RKcXll9kuvqcE99
KJSCTwmooACXYogm97JpedeIxOYyoEwpLFu5IUcigj9+wtmRbyoFU1DQdXgFxK15q3+taP7aY8pW
BDeHmKjQ3WF4jerElwFcXMM+mFG3051FFa5vqA6Iek8UKluW1YeHM7zKMiiemeHc0gS7arNJU97j
Ek4U3m4dl7wB8mDTq/TCPfthAR7i8RjTMUc/6DdXLhUqyV4a+4VefhjiLugpeDNAInDlFq8/ouJ3
9VOwsSWU+jP+U1oTigLa9BBolcy68OiYavvMzmX3fMEsQFWAK/E349CUpiGzsHwg+YftrGOmDDej
6uIGzTFvf/P/VQWYNzn5cPlaQ+m0WImS2y3g6QRkYF8OlCSoLQxmUAjmBkpwW9/OX3CFIkolMtkY
+UbKsCtjtctKW+av42hE1rdfRcfObPyvKJaEGLOtsOdY2ev4UoZ/aI9XSGSpylKkHFOUO3yvm3Bg
/vFJ8RqNIFWXq+q4OSCDNakDbmBIlf1kCj9Qz/Th3W6iVmDnUiay4+b9ZkkgV/miBi6FKRT+6Owf
UGh1qm1y+cn16pMKqrxyuyFu/WzZIlLIHjkoLWDSKVLQD1cV0q9NomYgu1pBPKC8LgmeDSACFE85
8DSi6RfPap2Uer8QfvGDgcqrUmtKXWwi9e4Y5yM6okpxaLEIt1NYlKmC3/BlqvgTeXw5tcl/fynP
+x43zCoE6bE5oK6oMztM9Rrp52PlmCxAm/oSMov5XKq2bPxIi4dR6dS6/fiaoaQP3Cccf4ubl+wz
kB/SYdkYGcbPwE37KgXCaSXND9DGGsnTL6I3qIZ9hHYQM5t+Y6VJaRwxWmcnBIEWSmi0fMjxq+y+
MSHutzfH5oSQEopUpvrWrsOapIzmP/MaaSqGfnITm9C9Uzt44dZUQyZKfoeOyhJyD7JcOukSdw+L
xNhkfKPzUkwNzox9R1E3MLS23X90kuxUOTP9q4aVLKG3XZHtxwuD/k3HYMroBZ1Rw0re8jgLRpXd
e7NtfzGBx+amYyxmTS84vYadcht9rHF1EXCLN9YwK+OhJpOYasqeB1/cpIfjgU31UqAO92/I0/iv
FtsP8CidcX4eJwszQogk1Y56x9HxKezpZJ1AyTzgSwPOMpy6AmRKPrt0Y6/faEKkcMZyjilrxbJZ
jmzntXQ21v/YAEKq/R3FtIrGHB3YF3QR
`pragma protect end_protected
