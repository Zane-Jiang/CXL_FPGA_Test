// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
eVjeHPbZGh990J5NZBAtc+ZWMuAfl6ydiSxFLsNYNg6VnZHbAo0n+eAjp1RVNyNP
hxZ+rVDwzAC/x9ASa8wW3VSKZL23yOTO+Vmw76KwSR2OSq5sp0D5HKLp557jv9jP
zNq0xIVXjYhOMohCVSMIqW+lqj21RNwH7qsrKnNiOLM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10576 )
`pragma protect data_block
ANqg/md7ZFDXpZbWfzW3sC7IQ3XI4XWtJ5kYuJJ50CrOzI5yYYWaR4Bj0SVNLrDp
RBJSxSjkFT30Od4VKI+FSGLgoZ0Hih2X3waaQZRLfZ80V3G2uLzDZ+BFkIpkHu0X
DnSqDSmEaWDo4zAFslJfqI487YEevJ32xzlAvBOuME1d8CJL4nus6kjLlzumseVE
WfXx+Jv9UQP9rUGfxE+PPD7m1Cc/x0wiaybVw5yaMay3DyQDfKCBqyNYJylGWNxu
JFVdvL39aa6at+2UTikE60O8qLfHxsP0oxblCjybC5OjMTjetfKx3JgnYl+PDw6r
7zwLfDXP7gwUtGxWtmeLphU0mc2g5tQUyC23hix5W25kptC5bshsThZisS3sOV1x
L3W3Jc9r6qgHBvbYSKicN33JxbJPYYrBZQmsS/FTI3Ty26tGuZOdHK5ZbCyKCkOx
y5n4UDldTmooLpPWE0VR7b2wA904Vl3oiWSdh5amgIbIiCeTE0Btnu/n7KnNhyTK
HLQEvCXjKMpY4ppiwgcenFZLL4PMGsQeHLCZ6I30+SyU8CIWZU7iNPIA9yPrOrko
c5dIptrBKks9gyehXd4COkHhfEirnjV4LKUxYJTs1od2FbSsMvF2bReJF8c6v2+x
yfqntQHNEY2X8JwUBJw2vr3pMAdXly64WIQzwaqbPhg2OUYg751zc7LsnAjXPBku
8dQ/uHQNhcqDC2HSRhzvuFta2GCJHJ44Et+ZvqP0UX9PySVK8nVyjCu6+/MI1IoI
Rc567YfJ4HG0797mwwLgcffugdRxjhfX2PXagJfnMcJ8GjWTB1Twk4CqNc+p/iyi
GNCmAsvS8CyxpmVRNmfNGrFAsjmRklOhcZyL71bS0Tp4zhINB3jvRUiJAz7NZN3+
T3h6fMrg7TsTD+xmbbyBQb/oHmJXHedcACO+QHP8wWjhYu7WBJMUtO9Wd8HpkXKu
SW5zIlttdDWjaZe1/9u5zShEhnhR8Ar4uYxV7Nw850XlMuAghPc7G24HwZ6rUkN7
UOBOaxHwVMh8bgLgjYgXM2QaismZg+QOfhuNnXHjxbcc+8VsvsmuUcERqWDO94SK
hxgEMJ2uUaATRFdkxOF37SAYBwAW/HUkgbBix9O9Ct5LnfQSvx1y5jb/xec3AfxS
txFXMdHUmuuzzVt34S+XG63/t3MeoVnxB2LPOBF0Uu25mX7egru2ebu2jGqEIphN
T5/mmapVYNMBAfkEK/XIMtLItTolvnt3gDQkVU4ZpD68mQDMJ5ckS+EkKX5/G7AZ
7zowtRmhEjiQ1WN1OARvX8/vBs5ZzYgW0rS9ZVXiOJ9gJEwr3Ys3P0lP4ZCQu2nA
mcCwz/h2v8ndTadEIHOOamCBY6Wz+M25OnW2GB9w6wxvmq4FvV7J3Jpmmy2YV7RX
yHPQlP9G2U5JN7lL2VTNVtk28l7nbdilWO/EwclPd3sfbvjA7U8EmHoc8q8c1M2l
DaiJgp9yTGkgLOLtvUfDs0Hj84CrUvZPV3GuRmMTSD+XfkIYc62g61hOB1KJMDzj
+WKoDlFQbM9n+kj+g7Y8DAJdYwnYgyrXRPMZQ06pXhV2xGFBe1naDQqZT3PXiNGh
PC9pEYtWgJyyrxqvk5eJZYijOwPgzNodkNns615wAVOXPM4SgYsBCA3LRGFMkL3H
MWBIyyz5OMIgeBtjAvPrlHxzeTj/ab0YQa17DzIO67TYekV6WUrEIiCaTblH7zAu
HNCwqdk/KyXEVjwNg5yuLHBd/ZCAUJ396bjQhn7KtfQufphY6jnhONsVZMWiQOTi
7nN/GRFYJzWtzoe3muWl07FaBxcH6ruvbYEr7nMYBR54iA8pyjS7XgZHIH8lCCkC
zqRqcibK3lJf6SaAUcV/EjfLUb5Kafg0d4yFJyZQbX8rZ64lhDSTnYiQuhzDGh/a
CCHpcsSozsMrI/5BHgPReK64XFFtX2TfoaQMkYGOjdw3fLH/VT5F+sYWp5Q0VQGw
IgKMIBg899GR6uy4Dz57NDAaaVIAaTvcPQmtdO6MvZ96SrqEHx6lt3KfZZpTTkd6
E0WXhnw5NkXD52qlWfGsTRAmQRuRZ49qiuyDyLOrRrJ8W9Wgn/lqxuZSxsNF03Tx
L4wY0fBXm1zPbrTRr1ngsF72YAIlgeQDs0l4EWaeJtMV23UCT6KPCL5qaoSrpOMp
9nOTN5bvrxzJHm44OXzMHkQ2jKaNsUiPj0Oe8J5cz0FTdeqwiJwagGAStkVR5+53
GUdpi5VdiGBlReKJqD15+/p9mOUJd8VAXGRqtnIOqLwd+1D8zSqqwRMSOeeO5lfR
ayiWMQ3mCXvmU1oqv5cV6GM1cqBXg+Zpaxv67qnQ0/kXkb4LBulHQ9fh/fqPPy47
Vd9y3mU50z6pD4obp91xws5BK3Dy46xcQIC0nOMQYRNRZQAMsUp2MRkN/5dH3yQN
Fgsz7ct9eSGd3m7yctgFzrNFYvZqF9cHvJ8lYMBTWAo5dACcyK6BaaWPo9/ndxA4
lIvAQA0G1LFlu6Yepa8EA44+ju1rdKA8zOm9BpDbVUvxKdw+CPIcLFQTrP81tGck
u0vGB/l+ZBj3MNNKxs61f6Nl4v9ghya8dDTTKefiOqsflNYgI138uelaK3KLDXDA
2cXSan4drEUF7VKy3iupVlENc9fSgiMaXLu6OYZqdQCeRJLN0ikZtEkdY5ZidCt/
jPOU0MxT0krDRTWFZ25E9ZPllCujUzbWmRxibN+rSRJAmmRXJyNeQ+/a36tZlTV0
bLqz54QpNcuhHuswXrWvv7fjEUiROuPrssqXpMoNY1pzQqIGHyshEi42PnFe/hPE
m8fdrlB72FEApgMWMMmKD2c77a21YpmsAecdbNwnlo9diq4CTnodAapJEoEGyJZJ
Td5O8RxtcsTgNK7+la73JB0OBBWWGtkcY36EYS0ERnMdAf5+oiTgz83YCW8dAyha
wlozBezJO21BNRd4yM2GBIXq9VuoUXx5KKMkGJiLf8dmrgU4gRMd/f4Kx7lEVHd2
aE3SUa2uQzlrFi5xwZ3l9Y2A36nchl1RellkcmZcM/xRt/W4q4I3/HEN0IO7/KY3
hSIwJO9HXIicCj3YN6FhaGZgFXUQbULVX9nEjykIpbv/NSlvy//PWV7lkdsazzRz
rdkwDu0mjGvoJyHAfXdsChIyn4mCeT4yn1fHxZ89uoHVOqoW3KFBL5zpZ0fgbmmm
lQftjS6RrqvanWTnMO75f/+5vFRMxN8/68gvZ/vYaHJ+wK4h39rRIXpp/H/YX9q2
HQDraypwDGN+om5KCVjSG8/G+K6ZU6TCRyd99oKWoI8mMJhkhWSCYRGXxfPtRRFu
2l55GwAUAOWmQsKmbBkAbX9/56JGY08TzXfaoaeIdmUo8irCxLIK0GDm3M4y8Dib
adqxfr1GXeUzvRn8srzFA/o99kiMbgD48nH7p6BRD9UA+ZDBLpNh+/O4IfFmVDWO
d4oPhBBJg16HoudsYJV5OfSSC0C8x9Q56g4ogl43ruGj0L5/+2Mxj+WZw4b+t6KK
61mHvn4ggHibczDNUCJ20Uw49w/PPSBUqixzAoKpnGlYCWhj4YWlNbFamka2f+H0
8khgkPHo1xpBNxdg2j144wRvFC1D5Nleb/AQ9KO+K6TwtudOL8uDL55k7400pz3j
+a3R6BZMk9+ZK8PhhmPIG53BZJ9Ndtmm68tBRhi039CsIsfd4MqSeYmMe9WRZezU
XyvR2+AM5h3jhQ/0IljHqz5COkjsOHzZN43QuZ7bSOwNk54thnoJcqve0ZHLxhZR
rhKL4UJM4UXiygBqvdJ0LOohd4W5TVDv/aR41HAz+HBOxMnP+p06IJJaeR5cP0NK
FQiRnHGpDtOdu+lt02wmR6eQEZGumOaCVjbSn3OwDPTLah29f9f46kt7EIQeJ/rG
8aXl439se/QtT/cztEkJo9G85sn1X1HBolWdDuwQJSgxtabbOV2PnBq6XqmyytOJ
ce9cXY7uqvG6NBTh9Q8bk3IfLn101B3Yi2lmdDu+fVSp8TPBZnvE1psmx4o08r0e
HdLbpmqZ0lvrspnR4A4+FisrYYHzh+HbPleeVo9eh3wWLVQJpNayUGWlugNVLl/d
tYys5gCUru+I4PTpybH/DXrTd+A0l5Klbnjotb/r+hufNLjHBOANVGjby4QGPntI
xl1Y/7wwXHGIV1OhI5lya6mnDpu5Z8V2f7vVCzOVRA9YAI8v8dKqHaSbKd1tliDH
ovdr2l2BEtui/SBeEDLeFRgsIPJ1hI91S3S0qAeOebFJm0Kvt3O0T9f9JhZ+kxI0
DwQZkeMZ89fv0zy74xJV7OgfVs6UQAarFdsRpWpENUx4kazgzWLaEd0jWR8eY9HF
7LLxRp2cR/hSZrJ5Q8BKBfwDzqdIqyEWmjgyKJf0NoAge529stXFK5xOsmUNUGXF
rq9OVMghGsy2KGvJrxoqT7tkr9EM8kQ3qOWtUSu/RUmlnTpg3q3+YFzeDTRNziQU
CP2SwrjcnCT4cBc9B1Ow95Etsj7MYEOlwiWbcaJtUsfpXxpmsF4p0ltAyjw2naC7
iIACdeR0cHb+xzs9v2rsaCcAOZ7H6OJLcnKI+AHRp9vPaNqTxSl6ztYHVvqZWbsI
Ys3AUJ4/6RYnoU2ETHhEDzLuvOhnWuqiTbkD29T+BEQIfKiN9Sp2kxgJjX9/NmU5
YvKC1c4S9YtWVh8QEZ4EO3m5c6z1Y5T0V4FB5UaRbJchtaT7Oy659LdQXHtyT3r5
PHvu9ssgA2nlyKA/UevDlepheuIt+4qffthcqdYWFbAZvjRdeI0XYU6ZlTYqleys
HIsFT1qp2da6gTE3r9cyCNScAk3x7YT29eJH9Gxt6KhK7K233k3LRh2Fq1ZN2Bfm
MhkIy+KfsCOvyPl+HI4HXFmfptQwaNZ3r7e13xsvNaJMhakH6dvOry4paPeAgiLf
OGTTS0n3w35Jja2G7O5QJCvBn+XlNUZTR+NmSaAizQ5FjoM0uC4ZMixcu0vMh5IV
S5ouda6F7rZEg52BV4IYk+ho4zFaaPpI4M/jr5J8BEgeGYlcendSrYzt0Jwuzher
A/8R2YtSeJsBGAFhJ5fkVTtxIQP2Zq5v3JdWYcWWAywPJcSG23fULF+5lOfgPaLk
BHNwvnHNwJE0xHGFoiKRkLXAKeDcpURPO7LTeg1ZnIPqIp+XPPHmClag4MlTbKrE
DjyTuKxHCLyL1fdWdfLDVLsyba0JU/l6EHs9MWuDcxqdK/88wyE4V3v2/aYNw9ZP
Fl5dMjlTIPTY+bmzzLrYnxZYDptjnpH1SF9F3b8VqvlU73w2ZOFmR9OgiFJLogBM
nzTlOlPLyLUaas2F8W6fo1/RmI0AmtmzqEIsa9HDouutUN83FmgKtqWZZvjwzLgw
QQW1axadY1+TbWFoO4zjHbvlG1LppEdj0fuJv2GoQmIaGfaLL57Hgu6qts1dZfiV
zmzySuZureyfPU4263MdIva/N9Bsi9FZFvy4pwWPBvei0MQa96bDvvVYRdl6EIM6
Gtea67Kt3Jv9LM95d5CBhaPf9AbHor5K788hy8t4hm1+rUBG812BM86x3Y20dkT6
c6mmzJpkHx87Bq4+TyYj2FRGc6XyPAjqnh7Vg44d3bQXdWnGBazlKgrXAEYlUXYX
UBMMT8cwWdoNoX28Qg1MmxVSdpC9bC3G0gtYtgDwjIg97wJa4FO8bEtdY6o4K8kf
Isenf5CfKzROsyq39jRUfwHjpSIdSaXssH6rVBeji04BgZ2izYh/mlSmF5dSNIpA
vzsDsoHG+ls5hebtS8+3bbY/En8L2aP17r66hiugcmb6cY9CxIhNjSD6ahizOLCz
12fT15RPtWHjEG7anS8GvdNWlX8MtXetp5QKKIhwGCGvmH15bPOfm+t2nIW4nZ/W
JZs5RLa2pHXOV3EnKBIzWHt6ALRDU4qISWuyyPaut1uXYiIktn4FXiiSEIudMvEP
rJxaEgW4TQ7MEDUD4n1PyhtNuwfqMcMw0a3ootehXgqMFmffEUGaxypimFGd9Orc
PK/4VkU1QGaorOQ2p6/uS/lDZpZmAFOlZbiZp33oFnNYmFJVobKujtET6j/DNeCa
hwYiP9EGgBcxJIWbBdF/lPlVY06zQgT3SPbawE1Z88hAmtVMFoZto1Og+cHOHgf4
sP/T4yn7n4tRDqujN1hHLggSQRAdEVQOe1F9aVgkGrgApNGuXMfu7jELnATvnpvd
i4s2MaST6QUpcDA9qRz02eQC46v6o4c6KEo2Dy3bttLkXnug+J/zmrBYdIhzEvs7
ZVhH5Yiw3g7chFlFuJ1z5gTK17pKnaosDWC9kQicgqs5eeMjxZWwPccC5HOf48Xp
+GAvufsob7HTY6YGIP9/rOv+LKwVcEvxr4XhbDFaFI8XE7nUc4AmrzzTWjHJdIY3
e+p+z7z+6eseld9RIJphPWrAtmhTHhA2BFvatEmTPqn60yRKfPMvVGuazVpGoPX8
FLMah3v+LSWDgRicmUPWyw3oddqtGVFO5y3pNlz0rKWvz5ypPBxcO/gW3oE/PVMf
g2H/yQl6bsgQQrX2SCNKx+VcN+PqxVxU1hpu35PgpJ76liC/BVix0IzS6sDcrV6A
xY8OayQV+rxdU1jtudbrtb2LbkgMjgmVsL6VtvnBrY2ShRcXUYTDhrhngTH5QU2h
Zx3JOKe7jo5E8d/YrLwFv24VEStHtQBuPciI69qw2t1m23k91+PH47KgoeWGZqSk
FE3W4n50eUkdB+ABEOYYSx8JeMWzn16ZopBQetQ7GW0avT/+uo4MB8XHA/XxEat8
6ipOTRhxEhhjpaFRnwK+JtT4lSSzSv7wUHb8nvLzPBA8kM/ukA0Wpek3nTAzoHQg
9+osdUWwEbPVJzJkQMlfaTOfcLm2ey/mG5JUlwCG79hG8K9SyYpWT6TG/8H+fSEK
nMi64wO08fiAxK5p7RTVb3DwFFa9SUxwczQynTwZ0nCJgjejNnxYjHWGvNPYb0vo
oQ+0BU5Jdy0sz0DykpGpHJnHrsdC7v/ISVIkimNjyv+CNGhPUs4mUX0b/mh6NcZd
L8fMSEk43FWiUsV1jygQknin2YUXodJI2fJi7OXs9gmaDRZaYFqBfuU/k7nuCqrF
B7A6n1YicZe8a9bHiiJy0fCuN7hCJLAvb9mEJBT1GFrpEO/kWz3GRMqLXE0r77IJ
AyVZZdTjmELUcDUVrUMi+AE9bYJTOxeIIblkB21t2P60ic+OvgXYUdJLEUJ3INF4
4sfuV6z+84rG3QEfIwr6EmsjWt8wxbit7BDCnEi4HhfTOCq/zBHuOHpGPX9pWZ1m
ed/mEjGntYOHIUyfLboffXmgjoyA5D+bQKlMNgyfRoMRvBDQuNOoJo0iWX8hyuia
SoEbqrXShoU8nkxyLwTnA87xdSkG68JJgi6VNJjnsfWd7a1vLrl2jVjWVuV9krQc
rDTS2XeXiMxWIadlpK1PA+dDJmFNhsNMJkVEZ83f+rqOwC0qAmRDE+tuyxIvpc5K
ew3vcbGLvsmFo6mYo/bsioyUpc4IH36u0nh/siw6M04zZR/gOtQDBJOiJMiJbJCv
MnIQi1irTMxPLjkW0+0YxuZPCEUE3PzDnHyE7ZMjdvPSBJ3B2TNJhvwbOqOxJQGd
AhfsURBlnlydFsiz1fdfYYXmH7/+PfkR65eHVlm3QsodjswJMQ874DUzA0J60Ol1
qHL9Ecsjr9fvKQ6xVMpcJeMiqDu61oQP1b0sXaVrobmAVEbWD6j3Ssfv9a71A7cf
CWQiB9hJOZowOsBHPgNN2RNZJ7GtGrlVYuXdWx4qXaVME7foLHXeWKhsjeFDt76C
fqbhfQ2v9LVE7qK7lD2/AqwqEDCYf0FNKrbhphBzmuIcWQoyELWiIEUMaxirItnd
KAR62v3KPB9oirF2d35LUlt54ZESCiGm8peL5itmTa9BmAIfwzTHgjqUCzCbWNh4
iCyBiGtvr20hxDuD4Xo/Myku3sG0blmHWBZalr6AXuIM+jDNtY6fjpYNhEYKtsA9
Cp1L6WfWhvQYkcF8HyIcN/pSeR/7sLcssF6gIsBIoRD4vPOWw+Q/dKl6q5sd8S+z
kZ+XyGJoeADq/7Fl8hIUN5xlScczVNFTHQ8FsXb/nr2ZWbQRFP0Ht3/DGohGVjLb
rUI+6C7U7FFsEDDM3NUUsi4owLXMFbVtLri7LxLUeuXeA7bNoeaS0wr6QKp+R9KN
UjwiHZC9Ru20X+o6iJ2s2Et35bj3CR2yMs5qaFSkbayt9fu1N3HgegCbXjs7Znum
EJA2ZwG5jXnEl7UzN7S4zWiZ7ZPZR9S/MDlRSKAvW828NKKQ0CuVJYNDkl9w/A1C
4hssjEYawMQQtjLSRRyHW69XSCmLLzOuGQw+RSGS6mQMhIZvOhyeeYYZQtDmI7Za
S1AriMEkdeOGlqfmjSnVFwzx5GBf81h+gR4GJyMaC6cdZSAkySzb72sXDFPvXw5Z
RpZb/Hs5opGrdJBiZBV/35uEaOwic505x2VBnr6Ny4JmJJNXduGDO6V3BPSprhod
WrOiUDAU4yxfvzXxPOudJO5c1zmFMnpmlHqUUCVNjnFZVRUUIbC4GRZ44OdimOVp
85NfDscqnmqCRX0gxd1gY1b/qKGp3hy5arC3woM+vQqBKIld63HDSA4inJ3rT8zI
f0uVwmuNE/Vco4TvIXc9RS4iv57BidHcxjeWs7vgx7LiM0FKyZR9WdI+fPNZOK2a
DXJGiijiTKKC569ZObNDNgsheZ8hTlWuUASXyt+g0+lLkjK+LeGpoNvZS4LEumAB
14aiA/3J+HNQv5nhQMsodkKKJ80np6UOD5k0Irvn1xrVMGitx1wMh5iL0/n49JDn
zjcZeRBAzaKAfItNEegxclW+NOTJq94oH6I1/jtnzG4C9h+6CLSwkO++UI+hf59x
glS04lgMEcj0981aAuBiGgb4kzHzg0mslS3c2wIggbjzv2P9D+EEXOJUTPp9chi0
r/MBoSK2KOWVlfYV+gtpIFmtL7L1+UKbIirnUsi+IDhP4WSDq0C31H5lck+ce6bH
ze8U4Ba6Tol49mzfOg9agJ+3o/c3rL1aaGtdArhzAoEkjZn3MdmlYuWHU43+L/l6
l5b2fwu0W4fINtjKYtjjZfW+P9I0ghw3Z0pgf58XUf5YU6q3xX2IP7qVgRHiaRoR
+AS7oAuTzuFrQj0VKfIOmDhmr3lXZRplYJHGdB4aKl4N3IxWpTCoyDth/Z8q2+Ds
dymGyEWKnpqGYZtdVCjvJShuXOvqnHrLJDl+SAb5YhUgt9xkPCeRvhUJ0jn7ZnD0
PQ20Q2eXtJrlPuh43K/Dc2bUHWBwngxmYyab8hYWD5W4SBIPNusgn3qMCzBf7uLw
XX/lP/lHCemxhHK4FGkHAgrT6LnnH+sPhsqwwrVgLGRbSASLgHMbBIHt8EA7qLE+
e6Yktg03pdc68TF7nGbjhJnXZy8njrbaIaDuDU0TZbBBx5kyhOEZNPHxTh2/qVQ9
byUe93TD6ojY76+78cpfoP6kfUZLwILyX0ApSyncQoiWX1rMCjWG/QB9bLtLLJAN
hRIecdaAciV6WKI+/vDW0Cf6WP3MP2uQRI1SvvmkQFZKX09btbTUnWuumPZ/pZf0
Wh+nDJ5wJS5s25Ju6ub9S4DIunGwSFNaMc1bSnyVkj/FkuLi/rtq9S4M1H72RrX7
FsVfeqzqnnNY+pGJw/Vm/24WZkML9C/y7Flui8GJA5NiNQzdJNe8BSQml4lb6BW/
qi4Hmn/LE+Q3pZAlqUutfaovpzhPbgIJen5IXwtEUYbDtfPpLlV9rSCPmVL6vof8
Q6WzW6gfi7WabaCfKNVtZmyIufyj1jcYFRmiWCxhzDmvogl/IaAsNW/8a9ktC+ud
vxwVmPHZJ5xuvWlRULaLi53njtZe8PmLrB0wb32NF38WWgwjTLdjMvlefrDCOv0q
vpE5QTGnlZoplHMy/ThWtZCSIyLM7Mq8mf1+knnl081sN259E2uW0ohym+tS93zE
4BfNRgTBq34aBeEqJ8d0CdK0pB78TOuP2Bt/Mqy8FbAMi3o736BSHo7N4kI6r4tL
iYGEwlfaTDEJrT4Jffh+57JVp8aNTvTRToyklx1G6cigv5e6ISySRfPV1QpZ4f9r
6reuhhxdl3hbq//8sPFXoifWeVpV87WloRHcXmgOE5RXmF5We0qK7WUYNVEt4br2
AywSdKbD0LsPa2gtLZI8OgEQa+JWfHJiHoykHSUTFyYFM8tNqnKMdIVKPr1zH9Pm
ljm1DbVOG5KsazOAwt1LWhcc9Weu6Czm7YMTHInsruFl6ahWNyZAI9QZ3g5l0LfZ
9bjcbUWvpT/+WRTZ5MbUT9QZgwbZ/q71qYvktObvKzfkdEsoT0sEEUyltZlEWH+I
FedRfqAUA1Py9VZrXS03wCvQBk9KzuJntYAhuUCgYgyXgXvU4KSRU6KxMQNS/5mc
wB5hjwgnEx54JDv4T40l91j/XRIqs6ijSrazf8ogpQN770p2y8IBK6aF9O8j/0/t
ADcz1qioCU/SoRS0Q7xJbKLS7qqW1O2pFBy0Dm0TyxziNRI98philqNGndOs8hzs
FgLUSjqip4CTneokesSwAzX31Manc8hQiOzhTfFLBonEDm+U47rDpKl76NvY6FGK
Bdck/JIw5ja67tHxEqMFooW9DR5JtDyWVIS7Y76v7jui8npF9h6kI/aSy46YAV5e
sxvnEKBiC8SuyADgWVtwIMEQ0IJTF/H/+Fl9NNCOiWV4mfp8ljEm/J992m//X0QW
dl8Bcjh1FXjDQu+/6GA/ycfeob0lKld4XILZSAEwea2UOKyzl/uxwn671gPb7HdY
kzu168c5H7T+ucD2xxe+vygzl8h2M+u+d+a4m0/abussQxh0C1WelCmFEWg3OgkY
vrUlkYPAlJc4cDhCJrUUJveUxAFe6aQp5iQsMmQcUltZ2ggOO+6STbqSyX1dpEH8
q6LAF2nGK9Fwj6Naut02mMaMzxAtMlYKUHneQdqiJ2arB6J/OE72zZyxT7AP2/Ir
qMAkjWHZpy507f4EiUZMTE/LoZByo0i2EEhoY/cVNMJiwQzUKaZ7Y+iAN6m3OxmO
RhUUGjYEmoGk4MNlUUJwryWlYwOZbxjp3OkR+vasUxYXlpDxF8mSwkHWpX2Oo0Mq
ulXC+QAR4PVEhci7OZziekBPHRl1zvQ5MVfx7jDrVHFCPBWA30rK/Vd+LcZn8NaJ
qkrVCJCzm4jovTD4XQycxPn8mtzqj0Vdv/zoVeMgImRkke0VsLP50CfNRyLU77Hk
5mv7BkYsLsx4UG9lb6qaMdXmMMd0ritSOAAClICFsqUJ/TWj02KUeETCNUQJPAyT
/7wB+g0iwANFsqDC+rv/cQkB9VKPhKmVGhDmk+FwWD+ylwKiiW5CoyT3xQ9O0FbZ
l3MfpwjH8nstEmUqGKwBDbLSn98zpT15OdSUg8FYRvEp+W89JjPlv+i6s1LOJa/k
RGrg15qlg2sWfns+amtwu8APXSs1HvoaKR8FKhsdrA+3YO2L5SSI/AW2fTQLVjET
qnCAmrcCrh536C4M+9Sw843nphXJNYF7HDSvrRXi/AhSi6MTJo1EZyaD5F7jtHhQ
EyrMxAAD8EpEKnCT6UY6WyYKSsyN4OmKxTvBuJ453kumo6hpLvUKSc8T3/ArBYZz
nVpMmPb6Z097VzOffR6kLGQgRKNaPwg7+L2g3kWM4gYTnXeuEGVoiPtNtIbb7TBd
m7FsI9p5IoW1HSXBtSlQAQ4LzS9Hcc0irn2rSTSy0XLbM9I5PI4A/Pym+4u618UA
VrrpgYaDC4SCCnBFs600hRAGana9jmJMhvIWfnxMu5V9WEq+3Tyga1GVXVy0/WRs
RK2QYa1TI8aiq43DL2V1OIYVL9jBe16nAxyi1jJb7tNI+GVzUz5JAsA3zfH16Tl0
HRIcles2dixE63cElErDqNjwtdCWZgbg+7MSkiorCKd5E6Sd/927KiqsSGDVkot2
636ab+tqXEUc7QdmoF00pRyop2bYFf4J8Cx18FGkrRyLTEpq3UsYBYbxmHXrx0vV
2baumv+5eg6WnJzkVBwsqP9rPLeQ/dGvayexBlLDv/RP2r6vNmE6TXQRNMuoZf9b
8Rg5acX4Jd6AuTXCXJSSCMscyN0pOzIB9h1yxNblG5LCxq9rea3/qlATw1t6m+/0
QVZlTprT3mbjduCeIckqQn3D4cY+dO84yGbjaTcNnPnWnQddb5Z98NmOMOq5aiud
UKn9DNhIxgazo1F6WGvrU7byMkkmDg1COIw0K7ewvW6dRFcYBnPwR/qK+83HhyT9
YpXBlimCXUIh07Pw5J5pdKqrHu02stequHYj+VSyoNKspQMxha1seurU9wQtrI3R
9Av4Qwb3l48J5OkWpy6qPOLFlFO/eNduiDMNMuWyiIZ7x8EIqc+8YF8rZrbUM4qE
PJl7Z1vDrRBzFCYKeYr3ntIqg0hfEecSa5IZtSec25r9tIMJwMwHTh6Oqzlufhi6
eUmawvDJ4fm6qJ3mK3aKRi5XBeWRQ5AES/JuCMoYuYvdQBAiMqZRAnNjzSQoKG9e
gt4VzYWD984LnCxsJhFmHGdvvnC5CzWklbPtxFKXHBwyvDa3Gii9FKGcH9gsUS35
6F5yy/5Myjw5y9l0aDuf5ZYHSauB6+y/nu2EXvPLsVxsfs2vZdGvEiSLukQQmc19
M5McJYanOwEWDAxp5zTy03COegVsCFV0AylC3tkD8vRZwMuLOy3RAKZ+1/t61g+E
Bv+z7yapMS3rC0SWHsAk8RGzHJQD3EkcwqBJB+E+Yl/Ee9up9TAdDVI6fYxIVADs
Qu5deGtiyBmIDYjnWHbObpUWzoKLEjqAQSZXkIBSkS/7rumN1TPa2Q0E9QwXRs3r
4+TKHtjguGLlhTgCzpPIM3t+Dr+JLq4R7wKXYC2uPqIEkbdeU4HVDgKCsNrPNQ6G
k5bM+jtm9u2+3uk1jAazACFHrsgt4gFkuxkKpaGENHtkqaZL8zb2WyO47bHrB+D1
8yyTLL7FViCGYMRUiBOmgFAAPQmkNXlMnGZfWExS5XfFCuqRqvZ+UDmrT72Mtig1
fCaoHevfPgo3HAEwp8yoJy+Dm37Q89Ny7m33WKHRyBw7bqinXFm11w7QNDM6xmY1
8IVqYF+1XAvjQ9qe2aO+XJalcIIDvHraoYGNFR1ag+ieKofPA0GXxfuKQzzeYT+H
xwoXc1qvXADhwb0k9YqwNURRa2vJtuXJCbCvp6BUX87Nqx58BKo3/K3dMB78aB8P
yNP94JEXm54AkRv+OVP9VhPVOxY4YriCPBIU44kd1Q3TBFr1SrRIRwekALfG8qe8
7NiuJ5DxryEBJ0sBSpn2Ye0JWAySiI0S4Om/zy3NoDUWSBEVOfHCWVWmjQJrDPwB
RI1bcnwEcIqfcRAwlDBdPdm7+xK4iq4qCdo4jYAs8Ap7b6PP9oFvfMJs8EZB6VyU
QfT0Y8l0J10+s+SsLRfTJUAxrln2SnuFoNU3ZKD44f1od/6GVr3IM09gxeNqwgIB
lDV72fLyl2Uu+ZeexahI/tS0B3Tt0v7NPMgpNitUrCns2UHTVmfyDZLOroELpPIF
aRIXF2gTR8XeZSd7uM3Fr9PO6EZSroSrYMTxmRm05/ZvD5wKNppUp07jZnRkGa/l
Bel+bZQger2mBPQXfknN1ES7M/6OyXqshMrLFw/7DN+6Is9K0fV6aVS7RT8wPuJ8
0CII0g6FcfH24L8f+c8wdhYsv0E4E0aom8VqYREDDgbuvjt7QRn0MX349U0oNJ9U
aTxezRA3bvOQH0I8TWJ8n7CESHJrC/oUjEIudE3yVwzLoiVp+isLBLLJwF8MIvak
jnnvJZ8gXpgbHmMQwVKOuZ4S9NCRZB3f4LuYmRZ8CcWCzeU3eOktG80IDHctsJbk
ODzRItf9RpaOy4PdE8Bv2b1cx0/qcEMb6K9pcoqR2hAWPVDfmyjCwHDNdzE3sgZ/
X751x5t0uxYoK8/+TXVu0mlnQbC541gT8eDno3eU38Hyth5IvtDxl/v7IoxsOK9Y
EyCnMk3eODC1j6yCzt74OoA/vI4TYWcsgZcclBY5NtZISxGX2yIP79GlMEyLgkgh
m9Cag5PFP3AHiuJ9b6Yb8Q==

`pragma protect end_protected
