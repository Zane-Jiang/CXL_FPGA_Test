// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I2DEDWXnvP/GBDBlh30fwMmI8AVtyukV95yPIG36+kbmssUYJu0hVWwh44q7
MMPrOsL85uzy2ny2G1N43dqts34t1YK+m//BotVeqq3QZDxgb0tvJLytG5nA
joRZJ4HQbZNvRVG/V1vbNjnV15NRXS9ipvr0LMGNHDMjrb1yaLcod/NAqbSi
qH5fxeisib24LawxYf/KDzDYoGbLXxL55i2dhi5Wah45fJWjSYle7IvLNuMj
4N8inT13wji1AD+IwKDeznS3/YrrGnIuRshFipug3fDQUArY6WTLUd4zqc78
3XDJh2wi+V18bqE39U6hAiEGZub+q8h6gR2una/+wg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gj/iwY9xyOsT4ohybzynWKqFMIjs2MGgHTI2w0A8qbPyFq7GKhZfbImZDkXB
ewA3IGZPRzpbLY9QgeG95Hekn0ynu81dtjPVHZ3jKk/O4r2KqclufMOMx8Uo
n4YEUAhclzzkDMV+todkMYRljDAXrPmfYUIjRVUsaUkqIpnvrsqk7i7Gp0u8
FfOnRL3zrqDtFtCW5wpHBXjHfoKI2qDf9pBEfVCGnuv+ar8EqpxiH5kB2g1s
BGOG4fmw5w11dkwRNKI6ot7BOO8A8Cvb4ncpb7a4RjGCbMRL0Q3MsYLQWQli
0yV2ZLyGDh053WkLed/1g9ga334SGw6MNO4mwtD2SA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Yo/aqPuUqyVfnShg/oLf2/+QYi54Gl+QcNQXFMLVb3UpTIbNOA8qRiq7H8pO
RDsoLxTwrNq66xi0d/wGtlrKOIHLYhmOm1xTbi10CLDGMrxpipRz72Xckq8H
Tc1B2KAoJ/YUDBznDQ+90ZIVTsFCmx7X9h4Bqa9ehRPnh6I4VnubdLXn4IFk
A77jTS+g5AKcYWwrkZszw2AtISzu3jjQYPaWVbPg4/NpWT4KWiqaLNoxWztm
wUQt0FglEtzGGOiSi0x1kblkq5aqc46SV99L/OypOG4xa1gvfVYYE+OaQvrj
CMCZ3+xC8exuzrWP/NcmYHCvH6sUUHENDewZ2FnVhg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pQuFrqTW+T9W+eu3xSd92mz82q5IsM3rroPONTUoXriIkIUDFcR7LsvB70i2
e/V+RlYUGDwivfIh2RSecRTyZIrtb+a6zP7Gp8lw1ByMMAsBm5jmjc0hfh2i
iuTn8k2I8XiM1ON0xlmiz9du0+XmVls2Ey1C4SDyppEQmJ8qx7g=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ks1NxQnIg5NrbGiOLkep09hXJPkUtBMHwg69ntT3E9G/mUmCKCasf0p8L6aq
mVxVN3xYgAfulLcnYIipxpqizqbie1ETHA8LEAxacO4v4xs3bUfAfO9XQuxy
YqRdh7Z4hDOeKOS1qV+hRNulNx07t5ycXbl7rGp5ddBRNvCFYnaWVPhIYfQF
6hw13wr5tnd1c4QHitmJLXUPSqJNN4QO2rlFSuT/27WopgO7k7TdQpCCUa6B
jd1ttdUHnX0+1u3QPSVnO7OWLt3PaTkP1g5m4Ny614CVASuuStaw/c5IJ4CE
3ChGE2YhOSRw+kEL5SJcOt/ZuJtjMXHudAF9LEKBz1yscO7Y7IkASmnZAyij
if42dF0rMN5ZSwF3dHn8/Pzi7XUOgtbyvVXxk91Ubdt27kuplw0DkYJhFO3w
vaW5Do3kWz2MZal3ZEu73re2bmR0hMOLEtfzE5BaMbyy35vLSnhdQr1sPFIN
XWlA0qiC+jSCmoJuM+RKWdhwwGVym0EW


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
htMyBjGhtdCayCvCFlgfEn15EC9GLeCsfQfL2ImiyN2L2mDo8ztXjWM9/q1j
OM4j8tl240Qjw9cxCahlQsX274xExTwQrYEGMnYlV72bqD8mNrqJL2KEfK5U
fo8sLsegviTEz0D6IdufSvaUyz0MfDSUir3V9mZ8cNpucndBPRk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BET61X2JovESrN6kI5gKSCKBYaZr4IbBaMcSiQhuJzb5vjwFCRDhKGstWlrl
cMnu2s2HFSO+dgpRbpewFUugUOHtxon4HEleB5IgUKz9YOmLRUcY5QysQLJJ
gNE/6IcC1pY3tImyQs51e7QiL3uYcaBNfk1F2nOrdc7Q9gRuI8I=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 36048)
`pragma protect data_block
XI53Xk+3gOQwWsfGU5EpGpLH6vtFF9/mkiQbmNTM1U3hs4cPSpJAAp5K5pUI
+h6PwezVSWnVNhJ2FGMnFTI8fyrV/sPXgDRQzvc2nmAgUfsGkqrqJaN02YZr
GRNK9Tr89Wr1PhIH/uB9xMqiSQk1EA5RiXOnYSeww+Cphv0lBAKVjhhfa+/n
ZeEje2M7EE2X8Lm/Aj7lE1r6vVhAXwgqL1kCN0I192wY7Z4Puky3M0OQR/qz
8nS2UjWrNts7hWEECmVDGa/xyiuqD67T9C577s4ZEXDWsswZq8nRVek4NWS7
RX5kJCLydU2+uLn+rKlmld7lORUlAMNCwad9hDedlzWu21Czr9xjzK4cSapE
TtIssix0CtebATtzbiXEpdfCUAJOaSDqvLzE9aamhaKKlLxoxiW9igRh9Vie
ZXU4h+CsCx+0jl58dWmxj/au34CPzUk7MJ7HpLs8dvs852WAG5yCUAwPHuOg
Kv/L1OQFbOKPYB7PbH+3wvBx+irMfRnoDmjCJAc/I9n1a4TyDw9CU6oEuMBo
1KQ5B7lAXmQdhdZpV9Rf+uZI3rQR49lpsJNU2Icr/pWqGkc/hfQHUULKYsum
cdeXUltzXhHedfopK6TRSeCTstDW+p0+ACe4fPk3OpXpqjkSTPwJk20riQ+l
Ld6MqzL6xILA38eXImMWODfPpler4z/DofTClTVzg40fxews/GW1PrsXG7p5
M2kP5X72gx2DVaYKgEqY5wh21rMnLg+cJOz1e56qTFjdlxqdEp/K7bYPYkpe
YlUphGYEKNddIfno3KALVsu8w3XgFuSxpiO8N8GaPl/3JHV/KTO23zp98IEU
dJbmcg5Ecad790QnRn0DB4BgsEIvtBzVizC83ytHHfz5NZrzcdlOBVGTr5Af
uNWBTfAyYHe+4vWvGGfAaPhiJWeTdbY/3w/u7F7OA5EfM+6tfKtV4ADxdcsY
Ec+w6mByS/xjzbfV5VElx2Im+jIubBn+tunSRPAmA5tYaBHqjL9H0zP2bVqd
uTMKGY0ViAu6vMpRSF3NJ6IGl05nrpiJnvh9TuxLVpAacbEweSsSzfwliTw6
BNUiCnf1hi5P6r9MSdY39gqitK8YvmCFT9EdgqcFw9BDqYtbnrEXzf1fE675
dihQqc41iXW7j+Msz0KhM8axr8Fai01EW3WZ0iolshJqU2MMmQGd8Ma3Nug8
7WgID0yHz1HMXeDpWwG9m0PQGP12o3O/vkXpBhR47hDNTqcAKb7gQPmQUJI0
P/QZ5BxnTUPGmKZeH7O9Q5ErcHMISGB9gVVDiPGuXNV5GRLy8RlP9kgwKxK6
zYNiB0YrmhNbKOB+ZcqJk7iAUlTTKepb/ue3LrNj0zxB4N7nqM7oqBy9/wX2
26uhHDYqyYlBOivDSUr9FPRyKpo2NBGpCPqECIvKwCFMfO7SCKcd+dBOWBvc
Ypw5fjHkZH3O0d5CTP5RA+lFrCc0kx2sPZ3vYbsMKkRfwZq/KkamqEfQKJp1
i66bvQtrqd7zg4Wowxffjjmme0KE6pG4r5w6y43ypy4kTcgYS3ti5gW8gQ1e
W1XgqZDCNN8kQJ4hFfPirlk0cq+I0Iefsh+9lrWqmNpXwC+NYZKJfzi/CFCC
KBaBYGJ1fBKTUem2NEPoVcb0w53jZA6kBgCoRjWTOrHXSph/W0YwhhTl3Vae
GxGCkxdoavsudn0KoggnO85PT+OF1kODg/skCHLxv2iPBLDKfjkCQLywNTr1
GETCdtLoGioKDI5EQrQeU0c/F23lR1sfZXNBlbhT8rXrlw2gztfyWpDI0LEc
ZL7k7j/TGt59Uvxxpxbm2sg86Ft8+iKiDWAhkWVwk0+JM/gredBbg8Qc+gav
XQHtPHErsQheUMlIIZB72OHqfOzIbmcO9iQECvi0jv8trUa2jeP0DXOxoLvm
NuqpB6Ilcv/Ekl+7i1kR8Ogn/cp6/3M68YtY/h2vwHYMQIHsIYb/ZT8VRS6Y
6dBxUkqN8Ra2E5YrcL0KrN3eKAWSH+WhdvMJPdi2iNCpb925cshnkT9O0XvL
FlPwN4nNpnkGnEi08ult3YApIt60nfKPvnDzbk/1eWVTVAXR8+/uGdqHHlGS
2QV1O0vB3jIx5MpYYd7O5sO0Jr8Vc69sXYC6Z00F4aggoJPW0ghWDM5IWCXx
cc84fGsFAtDvpV/N8xOz2nchkDh8z2CvKZ1GwrxffvO9gisE/1xM3c9IhFPP
pg9cjn8Mg9abqUAre6HSTKnhmcbzxNlrFhC3djQx+GHUIkFEaQrZTLXZyJnX
9pu3OEbmJZzOStuAqkV4d6aHI4wz2vHszNWj5BVJBpzBucTL7k4caedKelh5
FdPQnO9Di79l0H/V9zOhxFxDJK2oJfoQf3uYx8A12oyMKDxOkjGLm5Ltpoxm
hdI1sQh+eDSgwO4MsicG/kD/rMSwCh5yA//Z+FPlFaCFEMjoZNURWLf/3h0U
jowtqvLedNYK+oYYqylasmTeJDZe1u29ZUNSTMDq5vKW76vkDGOJcDTvM4p4
00CgFqd+oDW4Ls46UJRrAVthbpj0kpCZynvhKU3Vkrs7PD3dfy8BKhJf5FmR
tJ+Heb1W19xdh55xx5TwaFTwaSx5k3gxoOxb4uPrat44tkyJbE1uZSkvnwcm
fbQggzgEGmSWqnj7ES3ptWehHFoKjhWR6rErtpR59w2SwoMtOmjSPypWRgCK
dBNMAQ9dWId9hsWDqYW7kJaqVjlgmPNw+eEFymKd4O4sxo4emboUOdl1dVMp
jZ2nU5DigPjnVM9+uwLt/FSnamWOWa9Mo6X718k7BHT7GYH8P3hMnD789WeW
GHQ07rasxIUFvOb9rcV/VbEljgYedPmuzjHgYs7aqDLUDd6+G/M1uY5q4R/W
B4QkkpaBapQACXy1PqWPIZcwALRpDK9sw/AEfXSQFBaVM8UlBc2PZ8I0sgYd
NzY6iOo6NCJoH5zy400Od2Av5MN9SDTZTEtuL3y/mYB1nuS3D/GeYUgqmLoB
BlrsaRJfy1mjyojfMr9I9eC8TMNxG2ANecRGB+a68jycQvgjFdvWJiKrvYzb
aBvPqmw7ih012uROj1Tp2Czor3hfsaDhmxN1+QLXGy5QV+T5dcGCjOuJ27nN
lTdoVbY2novxqXztSzg0+GjZcaUxt1Uf5fGFhNOjSwBR/SUFXX51Z8YWXKvE
3MzevipveA0w4l7b0opjK03hXs5F40a+YL3vb/DdvhOUzseesc9eIDEBDiFX
esxFGDCDNLbg/4SECmagpl36wzF2J2kkjDwVC+tLY/mvvkw4C7O73CBj/o50
g5dGyDR1fFMyCV3maYVGDgbNZWfHpfZcMfaHply4vVyoIagPv8myvMbn6erK
9s1xZtV35GKLb5J+TxNTFZaRHQeAWc2vZy8KdmOB+Eh+SYjudmHmUdu9zS3S
n1ZYjq//VS/96qnDjaqz2TftEyOsZXevG9q7deZzZ9sz4CoN+y1EqWdMbCkl
mliVixhMpqiKygphqCGHcuWD/N8Ws1OnUWWRYr0jFQTPLub+uKtz2YIcTFf2
zn2zQong5vsspk6ZcQDb/0mb1crixtd2QdhE/02khWmdQp5c0yAFX/mf6nTT
8plhc/sRRBtD9tgs9lRIPR10L2S1eJkO2qHlLUyzyrzf2A9SSeShtt/cjZKP
z4YzrvAxUPbbKu40kvNiIcGvODvWbCrQQJhXGEj5cc7R77vrHSTkkXdKWzgD
B4TT+SqhwOttSC1DSCDJFSsxVsH0LtP3BBUthZByl/3ZFX+6oCi8uYf7lvQ6
G3FnXaaYUAyprfAlbwz6l7CM3ijmXLpwIsHxomaqtChgNijUWlZ8R8/JYxVc
3BtmMFfyD0cYDlJEvtTuwSkmzJ1JdalDq6UUaJGLxY1GLrTzV16jq+19vGNL
hu3UlbOmyX11VSBKQIXZnj9Df38RzSJAvKdQfmrdctbWwu0RQrTRlXOCHS3a
e/V3UUWgSkQZaEq4F+zd4ReWgSgzF3Cy8NIUXCmas8JpVBIxfU1CCgbzfuCG
6qx2uoEqhKMqtf94mgxwcxD92qjBeM5/D0Yj1khzv8Eo4eHx8ANOrKiXI4H0
h2LccI9YFq1eTFP6MVJTr3uXJaF9iFLAYKIVg06ODEFY9edfde7fYI6yCNSY
zpJJ8fog8S7SdGhf0dPCt/5BBSH7gaXWe693MAtw9xqkhhz3cZ+6Ua7u5Oqr
pUit767Rofx9s1BdO1inJL/BLAOMnQ8D/VMsaWy+eK1i03djnay14Rx5wmAx
tUCYgB+Z8nEfY+hqpKWHiXrvCdBIbGadgXsC3yzDgV4a8JlQHpLECIjX4ulc
F/8hgfq/JyXwMHkL4Jy0fd+tciImBa8Sp2xXmcRKItBYoorLrR3gHhRkzKdC
zjX7zr4tZStr1ymNWW7y2gwbuDZr/hpm0xM7aBL7XsF/kRYAoraMAzKhWAhu
fEHKGavPRf2HDGXzoCRx8mM2MWrHrQ8pnecni7Ihm7nuPnp2G0KXgom1LioD
sMbauXl7IaYot99lS5Ds5JVBmA1OCtvqwE9BPCFygnu6qM5kIO9BzXenz/mG
ldbkcWDqverYurEzdLULFidy8Iy5Cc30hw5qI//sxphdiFlQiO0kI6ld9iK7
8fPXRsz8QC2phRoN/aoymgf3C1GyrVwDIkEDmwc20X1snYVcPcchISSQDf+A
MD8YCWNUks5DpWX4NZGZMMof9R8hflGcnU6GH2/DI3LYhIgqdq89t+/A4NK5
QUcjfAL74LHjxfQeHoSoqc78iQqB9QXv3O8kMliD0qNEcHkvvToMRooeBv+C
94l0NqIpD4SXy6v7pq0oGs36FibdSkAldiIBX5RpgFG5iIWIHKNyzptRpqO9
5gDjIYRLKSD/Xo1ap0CIi81Ilxt5pVzZ9vTRhioxs3R2rl3ekyrZ6byZxjUB
Ev3J0a0yiNSAjLc8PjHUWA3fq4LhOcoLMdaE/WGUNu1yaifYM5Z81vk+2BEQ
rHIg6kZfFWh1XetiFf96kBSVeynmFP/gt/qN5zMdjQedTeKMuK2SQ4+kT3oB
ORy0KGZs6Npayo6PGK974Xo3OxeceIjK9gvV1JD6UMsHmKotJODm+H2otDYh
mixxgBsdlKpSyYrFQwynv+FDawW9F9gAGDoDVgG2Td60yUhAZKHAIY2KEYs7
2Vyh/fsa+sSFszebT96Bk0iE+EOpNY/tEep7ZNZ2AnUofAUYCm0lvtYtLoS6
mRmvqIMFLKJdDxE/DoSryrtPUAxWcW5nhfj1gcq7NHlgvM9Bth06A5Z+A9qy
JIMXnypTTnGAbB9ZTHvjVCe2d6SYzJ6n1Mrt0joHGeK+RzyFDk+NaCA095wX
WAmzNrsHNQTWFs+XhGYdqpSjObGewY2FYFtL6ljuzR9UomOxorFRHRINUm43
1St+6/CHF+M30Xzt9A9nqsPjOHanMcro/dee8jOwqiHjzeQHGKi1dDRssldX
MBLakZHeSiSVL9Uvh8kdWuAmnG++jo0smgxkDP7eUA3u1K//STQjh2HRmTMa
pZIiFHF8Lm1dVm83aXD7OGtCL27stonMMhb932/ESEhIeLPPWn7YYF8DaC8D
IVVLobnFv6nKq1KMtmvisYsH1EZY/ib7RpJ038FS/dmYo4uNUNTHcw4f9bO8
faUX8V3sFEVkgvR8yuckOq5rP+Us2i6lIgHP4YYBDRm/US6zs4xvL8XBfrjd
S79CEoVMq0iJ4cbhROHDRK9MAxM/V9urfXsp3MPWUV5brOMG5a9pKaRyjwal
8TO71cB8alkuW4CgpqysiAAzFs0BFe+VN04IFi89+LOJG0vwHJjbpedIFYap
WExN3sGjhsfkzQSyb9I7wCID3iVM0DOgiBQLKPshHu9jUUU/Fb5tW3FYrOas
+KOHQ4KjMby3JldmPP/I65zFRzKmWbvXoZerKKdsI9xpwYoHpbSmT/jPv46S
Bm0wnQn1/xWSUtJiSzUxAQniMIYqZbazx4OAmhTT5BtDe20wz6Vyh6+qIAuF
IhUZ0M1WmWkrzhjiROzc1V/9PJbM5IF7b46V91zAeAMmJVILU545mAoJhrwb
VG+jAVVVOJHApx9ZVB4MoXSsD5Tc0hhq4z24h2/9jlFrrIZWsck7ch+ebeUY
m7w9/7o4tKIIyZxX9qXeKXHd38+8EJl/rUahPgVOANar+JQJy5+EkPUPFwBQ
VMhIuWgl70heDpRSnCE04HOh+02cJ16B8tknKRrIj6WZqpaFRcTFw4+taAwE
19Gi4tlUsRpw8TeyCk9XPXvWaC2xh0BM12QaFubD3UQU7eij6cKCRnHvIteo
pRgWRv0FAqiUCIBpK4mnxbq031YsMlohwXN/oIo0om/HufiOmJb1o7/zIGmR
x9nmHkSAp5vqNEOH68C1B56MAIBZBUetgAoUJxr793xxx5CzRG9t9yVUUI2X
UobWO/UOfaHU5pf8e5e0wPFr7Yvmgz2atXiF24YqcOXrljpXKz8jP/tU55zc
UwHJSRjI6G60Pken7oGrZNEXX1g5EP1D75cGVCBdiu6okMdE2LPfEq1lhXi3
Qe4Rn8h0EmFghkfjX5D2MDbh5vgl/NsjUvmDhljDg5jeYIWcXtkYYup524+o
OVTYhBtI6jwc0YpApZdRM8tqW2obg9pYrBnxZP3iIjylAUSIx11MZe5bLwJO
WLRWz3MiGF2zKXq4z688hl73TJ0nnWkcsLB/QIFcSkEuhEPUweqmb7r7j/NP
Dn0AlxzFl14Qu/mRBmjKgcr5PEo+yVbw27HZ/EJ2Pp5/2Yn07/khK6Nv6BM/
7M1h/h//N+T3xmckASRJihslWd6CzG6segdugww1BCSGf/9uM2a0HWPgeaAG
H7E3RNHDQDZl+9NMk3iRZdDAB7lwrhyy5l1Yg9ZL2qb7DMbFsod+KNXcmuSV
EfT95EOxm/wQkqUw95y2Ukgk7xrdXR2pZtbwTkXzeWFF+UJRtQHQxfIv+Ryg
wo8K4hpAUjbjVd0FcjbJzCm6srXItvYfyawfFtwVbJlRfcmKbSS9lJ39NyG0
PXeLdNSxTSnqfNuh9oS/V3kU+8v/jiDm3sGnrT1jAU3t/60s5Zb53VfE8llw
iRovQJKirU0oJPjes408Gsj4gP+eG9jR47odt+BiYxPewZ/XuFJV4pZU90xI
fqFCJ/6nZ/wMu6ChEj0XhhYJa9mk03iGxsm6VkeNGNyPCzodw19CCB+LJE6t
PTcxXKzJ+082u4mK0XVI1MAGUGyfuMcc102bs2P4t8lmU/w0dQEDF7LE/utJ
LIFJ+SQrF5wgipkThjGVvYOySBqcYB16uyKujf0M091kSGHc9C+gSUM3kLbg
8O+mVw1DVQoKirbigXjJbj3/mc/h0EJgiKE2jH4blHp9ZBcV5Joxf3wKi47Y
+0NT+fm8eXT1la8V7TOxs4QoCdxrE/Jjfe5G4yDyjP7ezhw86g/ifvdYo1Q7
N8t7m0GQhrPp2w2VhgE9IsadhQVIUoGvSOTExaIpPnShSzCH8+h0PSdMEvWt
fUlQkAqsmDs1mIMYmy2GEQcMZ/eWDULCjA1q0ppdy/MThY0YxdWtjQoWfT25
0XO8AJmx2hyulLor7j/DuKYkLqfsng/c7K8toRHHH4qkCxhMgews9bPsL/FR
1VD/GAGMTwwA4dFPAOVLMBRWYyqB8e+UQde33HaGWBeZAkf+vARvGJ+iexi3
ANSl3nbMenvVWrCRLTbOVQpEmTLfcPVhdQ87FKGqChZFWuT0x9sdXX4rmbxX
MDJWcGJD+PzNWP7z3omGIS/Quj7DPA4deiqnKgpxazvTC57Q6m7jTiVeDkt/
uJfCEYZXclFjIxTHvv7vZAHKStCMUdzeTRuxJwbm8lnNVU2JsAaJC8gOYW2s
W477L6PJEAtBVr5NrJw0E4Biyw1OeaX67HpvDlX6Ivf/IchjmmKu0Ui1qLj3
Td6Ak4dwCmeTeJZDctzKHJ3lAy5wb7VV30JIZzCFUlbPyMMozd5owt40ndCQ
DY/120xky/ZPki/OLcP37eXJpdm9rZo4RUrawamKBYMv7TE8LGcXbfFOgIxR
DYrfdP1WOLh0brU1x8qXRLbb1z/GSa4egKkJPtauFaqEVd5jlKqof9nLRUlI
6pYZg0MmjAqCbNe147+qLbVMHHi9BD9qEn6Y74/pzIfP+4rvsdqSTCrQHBT2
i1retUqklR+icBEe3ht/6X+E0eqqzG+pJTj+W2+mtSdqKnLPmQeTMJcXBT6j
dZjb75KdKpBZ4gjnRKw1sJrltwnidRtYcJu/yopWnnhsaoKF7LJbDDUMjYl1
5o6o2VoY4u6/JF0474HyHpA2WLKnl7+PYqZPfqcjFgakt23V/Mgko6PVsq3c
ZgZCXWCkJTUF/X+IXd6Bzc/0YbGdUoeJR8i6VB+VSivEDkYVFv8FRlfWMEHz
lXcj5XV9k3mDe6VePsQPg+6Q2vSyhx/zw07ahG4NHmICKari3RXFFXPsL8/t
1deAN9zpnSh5zeo82WunOJmD/14UL+5dmtmqKMuuGajyG7WvPjv1Bas0qJNL
cjPZuAttMAkRGp7y8Y/0UOJI5JVZ5L5t0hrE5Kw2XP6kRG6GFBMcxeYJrGbe
JBy5t0avqG0nJudIxFLf1BsycJfI1/AmhmJaahPr18/O969lwi+DuSXxkzdb
ZrDAc6IPtUJXzRT1RmeZmj3DoqRLvGe2oZ/fsF5h8EplbBLZyCUA65heOv5p
FlORkRG/iL7tpkEOq/EwCD2uYCaghMn0/c3h3OjTj9hpeP8XdtAsfORqyGaa
TSTzDydGpYPhDnjyWq+YOHmieUzuOBiGGma4fIuHeuJLsT/oSARTHl2nFj37
JWYUzuzg02J5lKFkxnYv4+1uMH/YkdX5tbVGkG/ebwiFfXzBKvT+UkNE4j3U
FxvdIxPvkAuQbyRTQWYcUpx9S7KrxlxWENwQ7foKkLdY7Hb8W+nQNdBAbRyg
QW38v1bGv8k1XMXgXn5efhWraPTNUJmTSQe7pmKdGtgeFHQ62JMQoMxUPYBv
qwRiwrjx0Mdhpf0kHm9AOSploKsMuNxNmMiDWr/gGxu45QO+fpKiVtynj8f4
h80RVJDz5s+1Wa1F1AVN5wGTMc/fCwvZ/Em9+SJerqY2UT87dvJa2BpZCQbc
5avNPWKC/eNFjZ94xrHBDOkdV5SRjfP1PqV3+XQwdnS4hHqCoTn9oNuYgsvR
U+j32k1mGq7X3FEvqsffzjZsRGGdTRPCkIyhp9dUTCX9/mUwq96Zf/9CXYGI
W5/nEBwElvGErOFLu1oobjKkbtZMT+EbLZr6XaCLwVeasVbzuKXwZjVYkTEO
141bNYgUfSUHqSZJR37Nbr9k8G82K84ek8Orw5b0U9CmO4b4i7QLU9eMpEcD
YKxekGIpOfRJAC6q9QkC/oksR8D2kC7jh4f7uzd67GHquCcLGbR6okn2LnJP
or9v3zTM1qrqgH4lwlkptBsm8LFJ6klsg3RuqrADBcJeCxsZ059oodWpeHq9
UpOnUF1JdIEGXMpOyECdyJpb1jrT8yJr0rHSd79vzdIN+t/dkBdT4sYzlDL3
Mq4IXblEWfkkdKlj7FboVh12Feqnl72j/NVnGCo1hJ18Pz9gTp/3dFvHG6oo
1cl0JpKgCE9Ms+D5xB7Rr9Moj+lAYdMbl+0uDqh7i3Bm5B0jUgZYMek/v3fK
gy1OrFUoVuE8oWJjqO9O+LE5ZZeNzOcOVUgqozQRHB+LZ6WUY4hsSu/5e2UU
u4yLDFuV3hit7qut0keZ2P3lSjUWWKDpZS//niYqVOHG2WenZjhh0T5Khy9x
fwu1DU4eU6v3oXGrMK0+ikPGaPO41qHhHTSWxk2S2DO0SJ08HxokyXgMKKmf
a0937+pDLX2nCdflwe0s8/Txh3fH4wQTUqHv5NCDXJW8BVAmlAh10eYztVWc
mMfBxvtVwPnC/zs2phrgwdDmYiJDLtkr7IYU9Fcm3++pPMtGVAQLU9A2ZkVz
04U3zFZzmp+khF5BzPlJ8nltzGPfocww9bPERuRK3+5sulA/DmGr/gEEU6wU
aAMXwDlP4lU6YWL5fWdBLOj3BQwaspS2FUEnFoydL4HfPY404KSMkYGBetww
p4Qr9yNsgq02qqECd2bWW438oCGQ5DFFzGUJ/S18FMM+vHws0PNlSF1LOpQA
LAAB893gPpOFO8unYCkCTQmUBTIVYqoR91l80WMFjc8WleSbQVVpl6c08WKC
mHFY0IrvFn3zPFdjzDPPS2glUxlt/4eO4/ilN/2gA52T6+3nYNyfutMGDzl/
n3R2TuryTvZ0al9O0lvG9b+kIGJV8M3DHCvV7FkxQKBU2o2W1YBlFgXqIGqf
lwD1bCOnXvSw5Z5pvzddcXcX7GKLGG62mE0gzMYxYwXC+jKFFNE5lltkRwe6
Om4+eQumna0kHCmHX5PmVcXAdcV0bm9pdocJT7icANfjwFXqM++s2Kp0RzNU
vH9HL9KFnZU2G/BZ91I9mgKUR2U5CibHC0yaOYstY/pvWuNgeauyv50Xyp8K
mPCDluM9paJr74whzjJcXLvv57TzyVS4sEKDCaxHGt3M/RYH2mcRbdUO1W6M
tvXPHnpRGw7o4ftbY2VLjx6EgNMcGzFdOBmY8lS4bQ0a6u5kiKAHTnQl42eK
1PuqR/vGVc1IKoVlX/nEtM4LZ9HG59fKL553W9Jou1sEb+2bvu1aVlPo9SY1
w/kxVkhFw/Ykhp+heGpr4oKAXntSbjIXCzvE1+xYMvRz6Dsa26E3nx6zCc1a
+CbmtTzKGxxNIexaIN8d9oQ4DuS2lNdGtxl/YwznJYgRFvALgEu8mu55OmRB
xDuyIJTG0rKFyfXuDvMC2YB5TiRhdHAYCNbaeeS4JeeXipKNZOgPk95umepe
vuRhWreK5brvs2M4TH2tqlBM5GdZNFB4SP5H6Wid0qtrXqaDhoFjVl+qjakj
N2ypDqNuzeE91M9biipx8eubPak10R6k7A/FndXUbo5zIrJumx5m9Jddj5ti
Y2gf+p0I4IWfV5UMKN9FMDzHuAiU6iPLXhxKs0j6CzRwiMU0k9S+Pwd2V8TL
sld3dmVkGgnIoj/MRvRPnOS8RJlbgVXC7ThePOVje69AzLviwPJPgsRzcDkn
SYNHqJlhqNS4LuDuSvtxXlTeSBZG9RE0Q4DWQA1Kh1ogBuhSrtLJkF5S2DOJ
ai+B4Cqq11nC02KX0cfnXN4tooLiPRkOnJI3biSbexb/t0y1tQGpYZ8HJZVv
R4LmhM36SPAzeK5YJT6oZycempd1j8Jaks46kmgxb63b0D8B0qoqEw2HadlS
NLWGmVthT6CYuv+nPWydRt8YLMlJM9JMM38SXfBb5uLPJczVdsKquV6idmVa
gSj/DJNoAg+vchVeu7gw/NuGhIbo6D1626b0kV2KcPIMEtquVnhOoOVrNKk1
WRcFBLPqKHluHoeKK0CDQ5yVh/JQO1r4LsxOnnKoyHnAkY+ypLQGblIUT9xn
rFP8tUUb+VrxG29vVQMADVYEWnJYTURzHywUKGPG7SKCAKKrcq6pL7hgOW/o
ecVpuhFOcO3ATGgAVADGLnvPDgrB6Kkd7oZvUBjbXj5FpeKMTDvHOZY5Chyz
B9TVAvaOflMhy8sUDKQkOKbDWEaVWnAsJIbaiAhJ8GuMBnhn+elv1tnUzocb
/yVQuNc8pjfSX7qp64E1rFJ7/yAj/3ovXJhQU+8fQ1cVwnn4fgkuDKwx63aJ
HIVeK34OvWXSyq64xXapRkk7bLmDZUOwWj6XZe+JwY60SUUFtTDFlsz4OJfq
N/p+UCj3s519C4oPBycHqiLel2UpZo0gw3HVRhInL+E0bIkdXIUkie3JkX8u
5qrIv0FJGfhHV1WFIYwGoX36brAOW7AF1VcjIH6+ho5+X7rVtm7I14XvgtwE
eBy/XRvl8NVwsMdNFN0036gsaUNDjTU8g7giilLpMnJkP9QFkLxzHyDHLECd
0eL2dLAZAaQs1IzTByr0c06dvSnHzOrWdbYoTDrS4Zh7uJRq8L3b0uknTYg9
C17en/U+heBXOv30mGXnjtO6KhjlbKqE1EwLVwRXNmL3Pmn3bz8k0gMVDFQf
Ku5pIohDQr0S5wzxqCCH+AhpEsH/te+F5ZtxlcIprMTM2zb0FnqMnDMVLxdL
PiYG6zDym9K2B6JS7IDW5ma+/s3hDD71MDUq9CqvXgVpKh9dQsPXbZvnjyBV
fR6r4JTrMebZ1JKJd9SKlAIAgE7fEmnxpndfu6tAVEH0m3pU0+smVbXamutj
wFCQY2yp7Lrs09S3vTHJtUli2ggdfvkGuAMTIPnZ0r0bi529TuW2HC2tYRiT
oi5GcyJ80aK32VkiokJzaGoV6CgvRTIcObeCidrbcDkbUUwjQ/lwMxnpHRP4
+/z6rk6SzIqIhlHPry8D7zYBRCHBgomic3l5iPsvHAKgG5bBUx6hBMgv+mIc
sWc6OedqRyMipRydgU/fDRnpbrIkEsgp37mf2UlWdsX5drCQkqf1rwvqsloL
BHMtOaGcBJNqkqNCvUWOccb42ST1EYV11vlPDxyGaUcuTfGtpUM1YWWBfMUf
WoUKHtc3E2lm+/Ids7YaEBem0ns4vh96IX46vmMSru6oDhYgMSQ1uyidqPnk
0M0RzI/oFu0yT88BnTVMGsUsA3dyGBz7QLPK3MVK+2YGwGeOOTgSTSL6pYRb
eOHpiDJ0MVzbyY2CIakeo6oUNoY+1sdjTdHqBhd13K5arIBZ4En9xByFHmDj
iuV9RykdYo9ozFWv1REtPTOQDl71TqkKPBNcIjAWnIvoLL/k1ussySnS7OMn
zLomSclJA8gGmeijJfRPQn5ZZSy0RdopmJAwAnEDOkkAh8hfWoYeJzAerM76
e/V2HeFUpqE2nYPcIyajvIKmQvJyt6HMSuWe0t2YKRSVE4gn36sLn6o8C1DM
FpWXGl2V8OevYrguaya3HnP4qBcYAID9Z1kMqGagsJEdF5nYwJpQ1hAWEKxh
ETGo8IQfJ53NCUNEGEtHBcpVgCeqtxbyBJ53PBd8FT4yt26HTlCzxoce/eB3
nZDYI3txc9bEpuHQpMY79aBMijvNl4lewD3aweKCIXPbwswyOMVsIO8RoWRF
R33wwqmO4NcaW4EzNGj+nC1oTAtwo48sINf3VHhl3+hECdN9JZBNvbkiPpCn
v8mtcwkab2PfUYT/5jDvRZ3LX1sGU3CWzIH6P5ZniqDiiQ1Dwjae9nf11DTM
DzZwKeUdIb+z220yGqzdbRXsxLDAmKEidWX0bIVDOtZGMwV/132ppYLjEhM4
8CFQhhD4YbtGbEgq8QmF5Ga6Eb2sTz3t77IxxXc3oNFdmKrfAiNtlmtY+8LL
FrR5uuaD7s3G3oSkRVXEPTmq9G+SkAdgTymyEDEU4Q9+sw5lfL+AOVh+3ENY
xY/LYlZochUGjgxYNU09aQ7pCsjTqBv5zTQi6Exr/BHql2eX0ZX8gNRJUzYN
TDfwQ0Yc5sTAWPzWLrJfUPZ+r8LI2ctSacPknGdwD4ImF6thydAViH7YsYN3
THTAcDnFY2f2/tMzwQVDdtuLwOdA8DL5HpiIHGjgibKxPGuHVuRFikQw83yB
GoDHHwDUNR6Wb7BCPh+rJA/3aI4L5ZNmwbM69kGfqiytXgx9tSOVh+Xqij5H
ArSWFLAzOUc4n0V+sljLvnlaxCsZYNnlxRWgDIMMN4Pc6G3/GXDw2jr3efQ/
tK21BZNnOQHPHiHnaPjQzxadGPxeC9XbxJJgVJnin2edv7CmOJR/pD3UC3Lq
CPpJoP/7RlFc/Gv3Jsj8RQX70UzG9bOAmF8Ynbb+47L4obXfQUf/rRwM+Yk5
SzbBKcAHRQTBKCTMjOxNL8q15nWmAIgNLp3o6OHC9aXj4kCCFSkmenU0tKni
PO012O57xB45N2ts2FN1JbW2Ocxr47deaMtt60TWv9MNs6X4aH0ydzy7Ecrv
QHlbizfn3pILpgC+hSdpSdjZEY+1n32jaPF4yF365YwlhpNxTE85OTq24DA5
uIdTc0Xt/tLav8V8I9ZzWhcZgAg78mTYQlJfFPnRO+RQT39Z7zVKOcAFAbTz
6brGche5sXbmbEo7b7RuJPA5if+33IUDdUcuj5VL8vNX0zEa13FuqQsHTHSU
SYCOME9qwNmyZGWxDB+zPjhvx3uUdBjuXOlgnJYmgMwgaMxmWVKekrdsZOoQ
l18HJSUPEXALxtv5bjh65SmfTKxvcwByaRM8OoMEhEZG1Q/FpVHJMyedjXFf
VMKxD+InGNZwgg09BmQ11DIZWFnmV2r4b+Rh0i22KdBUhm1KtLdQ8cfH5YxP
7PANDLH58JRQkodOhJEUZfNudJPZ3VH34+eYTsL5H6zb06UI4TC8X+EKHcD1
04V+R2EvNhLFc3TKBkLmTfPfaCqx4K/t1krXJl6LH5rQv5c+e7f9mBf0uY5H
P5Cf+y89nlufNlpXcBZEK/gGUIsln7mdAp1EiHcsGrm5WQek4RirTxozF+kO
ZxyiKP21tcme9FnmWE25OyKb2ZsZ1xZeKtoA3/vlUp4Y3k8h7FzhWwit50jz
mf4u0XEjMlUDcoc+slxYyFIGbwRoKhOferDVcEeXUjPL8TuRo7yCJoZBqng1
fkOgb+B7LJA5aclvRhLdXS6hi8bVPQXaR8+z/TPcgZawFfUTq4upZcwxO/2U
XB6uvYgrlt7+RCK36DlbXSVf3fm+Kb3IQs5y3Bdqfg10CUiZWU10JSuUfBwt
n3LDthQJgo/28Pfv+1ywXZHAYbzcwWMwrvN8Ol+Qtcun6TNiSSuTDIhRyG8a
fVoYFSdVaxR0y5wCRUXQz8jRsz0uv3mslRDy0CO6Se6sXucWgTT9eMMOrX8c
b0EZevCVCVD+/tt0XNQdZIougXl9hp3k9w6UkhsStRt8gIN6lrW4QZUYa8i2
3Y4ejGb+R/tzGLWSvnC1JDc60T3i94PsxfurcY6TByShr2OPcyabcXWVF3gc
tQfslbKJCDCB2s+mo+RVS1Hau4PAVK+8nECyRCvR5FCyyQecoZmjjMoCRK+K
Ml99YqEg0Zfj1Kk9WwXbGg7EnuKjXNxPeGfB4qmu6t16gGPQxf9WRFcFWQCp
aSiGSsgqLUcGQ88JtK+uG4nbr6Kqvym3GyOL57sfGEzcuqTouo3KeRyZYZSB
DLDAol06+joO3VQ2idBjWWdM3CVM1RO6emnXcLBpwow8azOVi/MOzw+WZDGr
jszQxdmcV0q2kb9F6oPvZrVGorR8muHTyb4bomRd9GIHXIrPUj2ofrfXUYr1
hyZ/G6bVvqAev5+eMS7cc9EO6JTP6MofIA2JDyAmcYfg1joFCRBTIoh2ydTm
Cw+bfG1/2dqLTfI6SdF9MKIGRoDa6si4GLMMUefxNETurZKKApO/z6KaF/ef
+IysIcZ126fsH0ENrBoxKxHwKhlXfCs9GCk2NBaqQoMHUqQnMfCOw6ClZklG
ofVqRuNIg2zduEoqNBiWNNSlFsoot8zJ/YvEforWPMGsaPYhtsDZx40YSFnH
6R47T+xiRUiw0JZjNl4KujFp9q6LBQb2u8aBf1/rCAarKxOPLQDn6aaAsJGe
ZUlbBMeQT33NlFk9LI4xHIXZpdwu5PlsGFRNle/qV5uPeMBmf2bGX0R99SVZ
lj5NU4Mpsyt33WyV96LjCbuwlKX4Ah+E/bRZYAr0CPpQqy/XzkNL8JUVsLm1
aVdpEAxoElKhxzpQKjZfxVlnDdy7dLTEpUSQYu7BGvlTleGEx4cbeCW6uoAf
RIp5x5zxcdoOUFuyg2bMxobiOUbOQu04gtLVjkIVMpYwCxBkAhnA6VDi/Odc
W5ySFfgetA+34l46/p7wgNe8kA8+vtAuLJPqjoe53L8Lwp91ETBxGNk8TfF5
3HHPgijI/gL9MBb7HUzs06C/U7iprw4wyBdYYw/9gYOXyW+gyn97VqU/oUVy
D/FhowA9yFP9xiuNEApksQ4c9sw5R7NIJy9O5n42ofQ5HumtCX2ErBrCdT7m
uGJEdj+RQ/jD5LLV2c5H4N+kmQpVpaYXWPMa7QsJNGN9fpd3zZPlHOVszTUD
YBHvjp2kVZzWJxwPMTWER2+hDTGaNqAum8pSc4Z2kHexQDV4JTFma1TTCRv+
BGRy9hoNzvVdV7AC6o8vmj3SdFSk0+i0md4C3Us2C+yrOfcDgzghdXMF7lKH
V5ekg1yNIAo2e7rqARm2uaBPIYujLMjXIKJFiayEk99SYXPnwxiu8wDBWssd
8kYDMKwzEvsBqh9t6mz5fLkIMgZsKo29CpGJbIDzP5bbIxohchh8wPHdB60m
oQ6yZVLBmF53NlXKmiYasabcMrVJxzu+SiqMmseJ+y5Hr8agAo8iXOrJho/M
GMRRMAgEZNV9D78+Tus6yFf52glW5hy1qrX/nJOi7l6se+DZveZxs1pZSJdr
nsDG4XstBoUnhYTll6cAuKf870796qYj28BD9You0LjqNw/tS8tBiLXETU91
Nhb643ghG8ldHdKeyFBcehL8MgjO3sRL3fPue+VBmtUWghRDkBpgm1yVBn+Q
StqD73mpWvgE98oQVG52bNQzTE9+64qHkBVDFn66zq/a4Llu2lsfnKbf+Ew3
oqFq4injKCOJCDBV4TCQYWyP9AN1ZHNNWDFOF6EBNYOtjqBZaRB5Y6gEEPVL
c4gcqRuRSS+1/2DOPhY/TKUX2wy0nElJD7gszAB15pRCP84NRCDyAY8wJHw4
5acR9itpAUl08ep4SVkFB6SAFBQXUdjI8+UOohLwKejwrmfrK2D7PTurFtTf
vPWNYz2Bx1CxzkVMTjfqrF0WucNZ+tRfevpGr/wK0WHRSzorb3hvr+5KtmhJ
CG2YH1npu1+0hk+SzxudwAuS/GchnMtzu08Bh/qS00zPKx3poWDEKe3j3RyF
p4HLLHcUmNBWNoJwORfhLsat+L1TWonVYOO/HPvDU6VTALPumJgdBayYEBV3
4F3s4GuwHVCSmPMjN+WZaAa5G9PP1RgILsh6gH1ZgR1OZCfAaI9HF6cigfYv
9fMFOSWN7kXZMEiQZVsqzeCcRobhk8WcZZ1t9IxTTboZ35mGycRglvsvWRBg
Txd403+vPPZed5B4dRa/1VbHH32c/s/2rhc2uUtRCqYU/8Ao67zyHPKq+Z4E
AJ8QhH3pY5IWi0yHD9N56uuF8BL8U9xyPvPu+0HwEZCR/Ej90qROus4BTWr8
HW6rjzVQF8geukGWADSNqTYP3sloVvz4TfDYkig/GBAXX54Uecmnoz/KWNU6
6lEFAs5oL6TmgyfeQgPozeHgPuXfqCQpQkRFpE88ADceAgN49uFLfXRtY4cK
H/uPgWIJ6th7J58VkTNiLOBB4Q5IvTN/6XoQxv2nX/2x1egaDii6ZCYszKUA
ElnzGG5183qigPusU9hQT/fdSyirDZfWk4g+DQ4KMVUsPtPBXMz/Tbig/LSN
KZQCOqrg32amSQQo59TQFREsA70ouTKGlyf2OkA5N3D/h94GHQaQxEIfhF5n
ymHF8mC6xYbVUZDoSCIOBMM+LsThrH9ddlWa601oDNKqLGhx2VnOhGivhMLh
Bc03s6VaViBC53frgf+JYYIT5azxnGYOkU7T02cS2oDbliblfIz3qtqRMyiI
jwLdVSrMquU9lW+oMfcNfhywQmK256nNdQ/7XWY9sWeVHm0A1kKTycqAhv0z
Mh/hY831BdvZ/YjrQ5cb0g0cfrWK/n/AYo9vyjhawhbrB6i4TqS30qQAoMe1
R2fXHRLBrLFYjlD29j9E5vR00ltLCF5taoTNJ7oR57jugCC+WBPLxNlsHRmW
X3ZgDhV4nTxbfipF8aaMAP7vVbjjhPAkIU5Jmppfl48+iFYyJkAAFcnb72/j
58kj/WDIG520BzmMNZMudTfMKwky6TmgjcuCx55U9dHaWTK6iMD2rgLnq+wY
Uvf7UJPCqbuLR1D/EO8CLgDuy4Lb0W/HgUNbszkGgkUGz5PjOTnxqPL90MuY
bio88AkI7O0uPXhRrYRKiU+qaU3IRRhRw6gGGtVhPZcFjLKF8KiHBrI8RksH
vDRMWdTXkA1N3TOnfZS9S1MtfxzS2jn6sIg5uXjvzs2KM9K5MYogTagXy/i1
iy005sAAjHkcQNNTPykNEl9/aQpofJ+rffHW02kiBliVTfHpKXUqk4Rx+S2a
FrNNHUHYwCF9jkVccmEqcF0somMnMzE0a2b/qd0vn7vRnQcXF7191QkM/8s8
T0cqSt4eJpCwAC1IdreE7+zFscL/rUOo6qpcoMQ5pVzyyt2+avf3ZFrVA0B6
6hDtmyjZcwwXn8Po8aEr706DnZ0VBh2fX4Rbl7Kb2Vr50OmhFGQMhQCqPX/9
68JuRXO13RxtfL5k7zMhb8KzYltTxmGcuAl6myGQhPzPa8qrITwlRWIPK4Oc
BjZ6WT2585gE+Zb8F7DuNuLbFidGrOwT4QwqixOCUS4CavFyvsKPRIThxY7V
LElZDBcSE2RBQhcgxs0GTu64ejSiroEypwaPKV3kBgreCwE+Orqerskogjb8
WrsuYMj6GRVMN8CQzkn7nKGf7IPKAiNfdXI9sAAPwaINWvd/bnF111wsKQwG
TmGjVFVJlTL/8X1Oltunto8X/bMU+f0Sx/53qgOwhuIQK5oa+OXKSSYFf5Va
CccnNrVMJNsk5ZdQ5WORC44mWzHJWrr9IsSq/TTFrhVfx4fkzsZeeFZvqstW
jEAZn7HFZx46F5wn2oZweyPc94fVWXC4nqIIDZu1a4ay/EVxoslFiAL7R8vr
C+4xc0XYzdmKPtrmKA6iiwTI2BLBmPj6PsQ5wIf2UN9J2Grf0dTiGgw/As9d
y+Q+EdxfP9cDxUm18nIcexs3wSMkGJwpcuwQ6P2qoKSZor11CdbE++5wusvQ
f2yV8zg5mL7jCQw2ZdaZuhDnNOl5JxvhaftV3fPnMhZea2Jd/5rdWExC0u8e
j8UsfM1KLZbhm0FuRxXwqmnoSjRiX0POmJ3sg2ICRE6a+5q0DO+uJ6DAA5bK
fMo2aztY1ZI7aPmJFGJUCBALbRUtj30cWF4yBjPbBBiU2PG9oB+8SWBjZD2B
mXPZ2AFEl56fP/5s41n41cdAdFXkwUnhgZ5uafMEYT3ixwBD19Y/8e7B74Iw
oVGgMX8vJcxL50YeWPT7uclGRfDMDx7VCR4Fecq5x590B1HdbYpPz/Hpulmd
uadDyISX2whmWNSS9B/LvR50shlW2Kqw19EMeVEMC6NEFUukEeZuh4g3sGeA
QebsfOJ9u1UTluNR6346WqKllqc+ZBcwb2hKcE++CeaZSOYxkFjhjdid0G5a
K8UuwdVr2dhvCV/OcDPuYZrUaquXAEzTnsnzROIlHSoNy3Kw1lBLzHPk+hUe
htCazHk8nrB01Nop8PMDAOC2b+274fg7r81sjaRIdgHyaPK/drtfyorMXZ+H
+90F+OrTjKzHkc7z1pXOK3MJ35w6j27gU49s7Xgl1kWsCYScLRvwA/u8F55k
eVHgIg+dkeWME7kDwe8uNswBi3OrGURDO2WuXyYdjQf4YM+bpISzjMxCwFyB
y3A3MrA3nQoYLVXl8/N02zj/5Okm+E/WqRzFZQ8CT5q+DVysRH54cJirS48n
iuWJh1+P0c3W2JeTiYSP5TmDbyhZ7yV1BTLu3G76P0DuG32errQnLIKUG7K4
Nk6blWx5rb7TMhCYdqKI9eCalXZjWMS4v4FHiuKaiPy40LK46f86TxPPakUD
0PGuOvesHJXjod75fBOX1ubbKyhjB3nRJzKr254t0usU4dwKskGem4G9pb0F
boraomWwnzHGMck+B5JDPGMPGdxdauLO5fKMvEt436FtRaNUqf20K855Jv9M
kzi/e8v0MkmBCuNU8TpYI8YbUBYPk5eEJBQYrPo6Qww5rEz5oXZ4w4ic/ZWt
QcZJwFiZB/9yUsZWZhm6cbRU5N0gHTEK5cq96jS2GGQl4RZ9jID2yFWvdDeT
8eW8WaQWH8slEDvWCaHH4kgqS5FGe0eHVWlRvOWS3QaKgq01yABLFgtdThZA
ex7W8c2BYw+dyvdY0hUp6HYpMf3W6YeplJt26AxL3Xb/yPsW8YIO7hRvWfWs
OV8YI80mtz4rZroXhehSXoDZuGLh0Vcgu/DpjxnsHvS8e0Zs2FNpT6BgYhDs
roR77U2WzPODWgy6gJkao6DeYzgI+YiGWkHi+75ONdOE30+iSRmxNHJFtc7e
0H1z0wnN5NH82IuFf8MJz57R35t+7YjzqUCcjzRPPV6DCJaVU+fJfwzBMcP1
osS3XGwe3i1fNgXzCsCIAV6KVB93wxNut62754NSuOXoaaz7NKhDWZQbpjxs
lKufy0lR3BtFsjRctXehRwQZKxJ2CFlf5I6gx5hRl9u5/p3s/ZfyBYQUvQHE
gEPNthAjoFOCnytLAy7jPVbgL3/e8j8DwO3qJ6r1oVorkgdjvrYM4ahvrETK
2LHBJVOHgOVW3lUjApNvdO2sFUG1qlD/B7+kpvngHeqE+eZ59XMY5E9Up+pj
hlm5J3YlrcZPE+KxQovbSnab0eMDrj/lib2SI5xOvbNhvph9YaeFKO2MopZp
VmCdM9dFUID1S5NwwZSoeXH8rIUkmy912LVDjHKcS81jd9CKG40ukGMMR3Y5
R0+2p88QH6RiVVIyOh9HuoRAeESoAwJKcXobyFm0EarJ22gPBuF5qjEF3WUM
qCsq+gOunVLduR9Fey1d1zA0LACk/JFiXrrXNhV0Nz87YpYk6vWty7I6RBMr
SK26cpaN0F7UnslcKlIgz9kMQGEnmkwl/4O/ZbdiCFFcFQN++RVu3DR4V7ac
+0tsB31mW+O+emdxofR5/0x+Zc7MYB4WJBeIZBESdtclRbMe1jFXxzVgsFwJ
lHXCRjsvJmiUd12L1UNHK8rR/nAbNp+SSYcwH4iim5BqrvX58mECplqg/zJa
vVIaQ4AebvtCikpioEhWcQqIDuVxPPShGwQibHpCXGFNHC3gZvjcBb93OGU9
jVky2NgYkssOz/cCvbo4vYfB4Lv6QfRuA7pOvW040dDVx+QgFML8Mh6QEPX5
zC8gDBmG5sPlUUnrWVYdDzCd1gJKEcileJrXk9LS4wGuII6fjoH6fDD9SZW3
7RZOCwzT1Xt0jrQHUbSna3UywbTO7LY6goN04FnnYQB4t6g2lMxEh/9v+mcv
LtdI+GyHfvyPYD381JzrDORVgVhTQkMMpcK5CkRFlmDaE1PALuDpUvmSzVqD
tGXAsfoQPjSw+g+p9hwviXGUasJbPw0/nOwx1BtQOHp9pDNqFxmDvhn2lWm0
jWH5fso0unOyjJ9Igop0aBK1GZeXM/TdH8gTZzI8NrSqdrLQ8pVRG74Qr9hg
lfjgoeNNhNjWlzckG8u2MGvY4P998eSjRMSOAa0WLw0OOR56ApGPjEAUa57L
Q+NvlTaGY9tQu8acBG8K2uCwFK3sZ+LiLx27UAgS4DhW9Bgg0XnSCe6hT5w1
HSGFGtT6xBI9sCyYaqOXHxMefOntYsHrjawKT65NUAOZtcf2Nlz0dFiUqSrv
yQ9lsfzOFCtKkXjYxOvN2YwQ7v48VdB6UBxQXDpnDNDcXmS7yv+cLbljbE7h
GdRJ7rhPOac/QlrW0Mlj7N1NuAWZTPraXWfshovyx29fUDjLiOVBvnXucvkR
977GZS0DIHlgHtPsdIF/FE3inmnscrMosnX25bGiyJ0hE2wqmmC9uQDJaCOJ
5f/wYWOAAtr1/TBOeP9X+F1JoElCLzAkXtNL0DvXBgFIu+mchYFoPWM2ITy9
+ssjS5kqSM/qxx9zwp46K9CmkxqG2Mx+cKbPR/RSfZLBAizymjshtY/rBZ8v
enXxrqwQGWs16siAFjoGHlkH9rPKgTT3nhrMMKCldxT+FgpT5F8G8cu2YRnd
ZdxzDrFRICX5MHEIwgDw0Na70pAO0lJt7XEH/mAnUHXy7eGRSqRG9ifxBpMs
YV8Cl2TAQK8q6yQ5ebaJZXLQFxPD3T1+9jCoV861fHZZx7ajFGEBRTOw1aDC
gpry3jXjgo9jpS/KT0Eh1GT16RI3BhnU1V/22iH11qhwR2KFTEaOf4NWUqZn
VRZL+CTB+8RQ7q+FL3wnbhzNYlj9D8LeW4N2MO2T/LvbuxrMyRuP8+r4f8sy
/KI9x6Y4iA8SKAS8ll9iJBRfu1FUpktzAhSu8URBTYSClNerg2DmuDi2NoC2
HOzEJ30x2vVab+HQUy8Qa0eJrFOUNqjXld2xzt1NRDX3IX5UsXIgfYMJ9mEX
CEkHP1Rdqm38qThaCtlgX5SOchk5OffvXmzSQaO2RosGmEAa9vtVWwe+eZsJ
An5S8EIT10W8HDeMgtH3HEle9db0ZapH3zLDYn3YSljkh34mSxUH1MByKbTq
VO/uwmrsH2Gm0Mm4kOepj9L/3/HdwYGT+t8oSLgT6DW93S3dUnK6jwn3akK+
4uauY9Klrw3ql5aNnsik1VxKHAfb5KPPmlMVc+dbXQv5HL3fRHs4xVqWw5vG
Hncr76Qh4UJ43BW6ae2VmMLelw7UdSva8jMspU4rjuRlRoCdy39ye/37eMlJ
FacuECUUAyxSFQQPbq/e747UveQn0he5HPjV98Jira+xU++WuOX4YbxTewFS
NMsgioC93NW9YxgQkoWBfjiF/6JMUrj6hmXecy7zMO7cq8DPFfzRPBrZqJ4T
JnXXhQvKxOK7Kk6dbGTdEgFzC2Q/XhTfpM9XdvReygvcdYueaYmYTKq+nJ4K
DokqBMacJWuDWSvAgQCllBURf9gKzcQXm+TW1JwS0zhlNesISxKZmItwkn4H
+h0Ts58U1w1osge3m/Sk38tUAvQFhRNIDRvjf14WNHUfD7uTTOqjcLaW/MmL
W8KtnrEDkLRi7yHfbY5w/yRaoBELURqLf5QibYSWIhapoJzWkuoS7Oinzcz9
vzlqFSLkZPvHIQtnHfqTzULnOm+qQbYS0DuKeCyUM+gZraTXicvkDiF32jGi
fS7sENtsOIExCHnVbZIAH0JtN+oLtlkUmfSB80J76m95WwYp5d8o9IUzEym7
AtnSn20mu1q8F/U1XUoHu68oDpaMNE4Y0RyT16Mmo7f0cNVKTZKDx3wavUHI
HEDqiE4Qx9iBWidJ2uHRjLRa6Vn947f02aqZR6RUmnEAQNM0LvVouhDTncxo
SPEZz2NqcBNwcGmxdK6aJhVz05BzZzb1zhqQBiIvoS9iCYHDbHVemGG+oAV8
RjzjAnD66sXI5gb3Tnn66pbCc7k/oxfO8SpW+1uzks5gVbJ+3+PXOSnPPpQl
v1lkmSUHUZXT/neViEO6VNvdm91m7xN3b971rTIydoBiD+bhnrvSzDNTui9p
Aw7rDHd/TQaDbarViaOq3Xh+qk12SdcmgRlWw0Tk6RbTKhyRGbKHXkZX4aUo
l2Ihl92SwE1CrVaXvrsSW/tSI0reErxN0vRonUyiuj7myZwPYfYgjtNGi/WR
iVVygLKi+xyAWEDJmoKBoTOtSXHbqlmBYUaNc2KiP8PlKDVgI/s3SJ90JlDu
L05pGkkQVYPejnT7CTKdOXZv7jFTPa0y0lA4XzzyO8wpHVGlrZwDM1Hbxewi
mQIHTuWmGQMv+MHu5vZRD9oJgh4DM/KbKGJehFGYEkKb+EE7wrdmdw4hOQXN
70tUaZ4143RqexbMpEFHp1lK+JxI+lNywaE2qHQh4CGfwhg2+zqVgsYCzxnt
fBrAls3h1J8tAxRtgVqeis8foYx+6EcFmYBCMC8D4BzRS32U7UscPYj/9dRI
mkPkNum08CUvpe+DpNDEy1iQ99gAQ3ql68O5vJt2a5FZuqWozA+RNd3GNrWC
6OgXRpz8DZf2/ncNW9Grq8Umf7oHS0+7pQOHeXv/9PgpiEbC4KKBxyHaSAfC
mu3nJ9bXZQPTJZnKEoOmJIIfoEZ4sZe3bbt6SpVcyugl/fEA5Zu72qig7VRf
syRsI5v0Xe1dlDWR/8cCCdJMdrVp6TSWGgEtJ9fdZabcFiiQlJgDa6bOdi11
sG9+x2Ge/4TW3EG25aZrsjZWW5D8MGeiYfolyf3wulMoVOycouNOy09Hhfh5
nSmoh+2uDJpSeZ8S1PhIsPbyJvoD0nqjjAc9yg8mZ5oxVl9jGL3WF664GNWO
1fOrMEwxnXVb8/UgoleCEXjXEKFbtenZ/d0dcN7H+/b7WsgX7apKYwQGXrqR
GC+0PieCAy0vG/FGKbihqf/cXmAutgrdupEE4AIqAvQAf109VfQvYHEozwoU
Akq7ze3yWVHJkdTKxhX8KijZADi10yJ2g00nQDCEofop7yCLBm/C6TcpWhY2
M+ZDlGTdoQXzOP/6CK+p0+AxEd6BqB1qUmmPP7GWNk/lUatlLPUVqTLs4rV3
PGjGB0AOG8xfM6nw85yzX07Xh9cozoPlFVDe83SPF03jiU8zl+A9G+O6+QNy
R1yCDH/qtTT/Pwpi03Hb6NZK6FkEcC0stwX9WOYzCMo1m+fDmlzOfIZed80O
N+fCLR9k/0hqouztH1WiU05mbbsUDd85utcUrjw4dmfygPhuxWpanXGc5cI3
cS9d+pUqyesBu2/ipNGWCwrMjbfbGf6NZ0XK3HS3RTDhHzpcCZRfX/KErhmH
5Zz8TPrtO48dO0V0ZzLf8lVkJb5oXW4Rvb7o5fXNiPeyqnBRdp4IDH/DqjYQ
eOmHykkGqEeXvtwHyzDwAq0m3t/8NV4dgPY9hopZVJ66O9/tXwj2isn5vMFr
374eIoa8j/Ly9OERCYFnnk839aNLVf7crPBY92thCWP+b0BUf1NF1FNRUDJ5
Zmtr74cDOHDRUm0lDJ3dO1o/HEjsOWZTnHxGzlOkqjpE0aPapr1g9cahPRT4
KQAlHFzoxgs9Nfy4/Mj+SgwOr18guR+C4e5GaR+gadmjX5+WBaNpbjIB2erP
xQzLYEmGRKKKciRre+SPQ1DB+sm49WmLcaexW0R5diRsi/xyLO7xzxFqOs0o
8fxhCGxKhTMi0zYsJbpNdzVAbGqDghCzs4R+9SuCkYb6mZEtGYF41YUlrmCq
rku8LOluKYdGA/RilUVMnzvV5yR4eOIG9x4OdFKut7JXVVtXTUj3ONS2eQG2
jigHHsvlqSU079V8uCCMtYPlIp2fdfCkeYFQa+xtd4kcNbDZ0AmnDsBXP4Kc
dsf0lSa7+GPCPOdx+hZLSym2YyIriylquHJJQBBHqCiAS8wU1myxdvUR76qK
MP1mhTg9B/GxcOxxNk+ICuBbWP3giMETkO489t3dSWHUwHHIc8vUiNc/bOm0
NWSN/Wg9BMvpZuITDhBHRfoJovYrgKhN2L6feAgMRz5apTkHeXrTkI945IOh
QxmzcMol8UY9ihCQlQhPeYLjy3oirgxKjdrt/ZtRRysTWV2YxVFVeN+bnJMz
xO8QjUj+QsImlqwwzEj3zQvNZa6B2/qc48CHGItPNgyrRptJgMESz2uyhCnm
hiNlfR+tGHgLQKSMQPpbObH+zqGUrjvQgXwObh1yHdz8Pq4xcOpVHKUi37XW
g7GbA77wGCSfWlpZGLdBVcFu2/Dx6fERS65RQZOEcfBlQ0kRKtGJTbfbCgkn
wkHgGLY9J6f9J1MirkmrnvhoxKkr8rdeIOv7Z0gbn8fqz/8ZXtuMXvcFwuO9
iKwvv4V5BkgnAW3ynyjK8TTEE8D8aGLA7+Bk+nJyaKrqh7vYfSt7soiZ5Rw0
UFxS7JivqYEWyCQ97Xy5YQThCo7KYYhkmrYw1EAMwI4cGXOHly2pOw8CBV3K
mWhUJMkHfOOx7rsOzRTu/syXuqEGtIU/le1TGT0jdGSfrwCq3Y4+FLE761Cj
IIvMi2t9tSCmD4iut4KujS3iS5RvJIUr0hRf73K9kiHacWALQGXwb5PMZ2vC
jpFO/sAx/vGfavFELGJbWFkpv9hxcBoKlTi9hpKIzer+u/hq3xr/0HHeTA4N
0aoWKO2q6syREtE1648WIaqe+4D9kIYilmR3Vwhr4UzJZcOyZK2Eb8QE4X+i
7W7Pt9J3NSeQLmqP+22apk6/hL5H+ZkuIsxjGTYkLBD0P3NA9WSYKciMgeJe
CkoZplwCXUt2+l5IFQgsS0Qz34hZ9EFJ5E2AkQEOI2/RyEVCTdj+ja+B4gCU
oKmvYSxolW6Pm0x1rDwi2pTXL4EH/346HSQj9LxmZx1UC9rgUYVjWE3JRKm1
bLQTSPbafEYxxnuhhiDn2wDCyNYy57C5Cp8bUb3wWo+U2jD6MgL+vc8j0vPe
fbcKop54N56WJyL7WyEkhqL/adfiPkaDXF2Q10rKGbJ1WfW1yoxrLqf6As71
cvb6cd5bClKGvfPA6dhV//RZL6qvLawG+8SapCeabOGt0NCW3LWcWpq23HsI
ygYDKn5T8sJ+yYjwpwFiQZ0ub7Wfr1pk6X+kX12gTMyCmx5/7CL9VhqeHj6Q
EvcaNuSBZ7qrGje4Bb0BXExofSEbtTU9kVQ/TkaWI36ZZ19vIIHU60O9Nlpu
UnQglrbk9CftqPvsyYDhulRMIT3mGMEuNFCngDBXDhfCeeIhklFAGFQwRkbk
VnhUzFZYktzPFF9mvIKt3F2xzcGSEWbP8k8Po1tj8hzlGD9nryFYyKhPXwd+
97OrpyS3YIAcQsukilaHDmBUe2w+2z3/yOyKY9KMks2AhJeGq8mKlGbDer1I
P2YgadLKIyRp799AZG5og4TasbRemVq8r4dVlPlf2Hj4iLe/5g7EU1pFDdiV
9HuTeeRhR8tifj8uacMng+U3ivG5BbWlcvEu49HHSZlaOlkgX0nL0Cf/JAeN
PKRzSvYlfIH9T0JZi9nVFfnW5cbAObBzV4ckBkFOFSWElH25jo0DUTHXa07F
MUzKmvip1LuAPwJeT1iF+7mgtn6/cAC+Wf2WviooYED4b8/J+syk4h4SBExk
Z6RA1BYUA/CGx4Aw1uHK0LCZCwTsXGPRR6WbJTbD7oNv3C5X3PLOFUr5eApu
196yCj5fwW4kVf1tJFxYpIPhWPfHLjGLlKGrdJ8EdjUkJYgCsnrWY5Ps7l5l
rLGP5GW6EcVh6DOMSEeWsUPs+C2KuIU2hzXaEpC5Rjc2JroNvVQbBTMTqLsc
mYIhS2LKJ3LA+EXqd5cmVK39JiUw1v9NaIDgnESPV6vyILy/M9ofWuMzB6uy
K7wByGR02F4OMalO8NUpofJwlzKEQBDi4Wlbl3aDo49rP2UcIt313z3462VI
ty59JjKkLYn3FNTsENgDbyCZhWRLobGOkO2CunW7QFB9YZbkhfA0xe3Bl8RX
9W6C2ho5bhm519gcaj8BDkg0Uz1UI8NiD2quEQn7Tlp0NCP5kLMcnZf+kp2w
3agZrngZcvMeAq+t+IKX12QzJqs7QcqqM7/FxmNn+SeB1kiS/bSD7sA2enks
PVXucgnYALbuNLr/hZfj4rNm3Z4IJMu/81StbdHzJHm1Dw1R7NBPSu/vofxS
j9rPJBSewjiXXkCmL59SGNNmpV54hTco/rosQPPrlKF8syNf8bMgnjI8eBCT
Y64YRho4gB2yU4DWvOipF3+g/wqAHO2meBq3a/QsyWUcRC5tzYPlw+puehx7
LfhUW7PPVv9Wn5rRKDObBzkreWGLlBx7NFwXPW173QxJu4wmPA/hsNQI2HY9
1ob6K5isRnlThG47xc7jbjEkIlIF8QFr1u8Exrq3sJVVQt7ayrLazFN3qtjW
Homi/mMGHqBdBY4PyJ/cdlNo+rfRqv7OcFRAlx/3iELzalti4BAsu98Nm7Py
IcbyVHNSUZnJzvySpLHozawwzu2ZqDvYTc1zEk663pqwpsyW/c9pnW15yWoV
Ar7pvbvLucdozGEFJvcqEzEsx8jlZio4ZefcxCzCnroGIJGBuweYM12S9W0K
XEdQknB0eoQYOYB/RGtcr4RdSF9O3A8E8AG0n4MeazuNqQhOijpYvMPsEBvw
ErGwD+34+jIYPJjAZmIBpCNN9NezfKFophhNnrx2kVEbuXpoV76daypEUHTX
9OrFL7D8WfU8FB+l0tsqKamdxBReVWOuWN/fOwTQ4Qa78Vw2V4szfLTXUCp7
2Qz663PFuN1ly2jBbr/vXBSIWuQonsWDvzkLprorP+eJqkJ7d8E0FjgD3m8t
HIIlfmKejEwtr8r5klHsqLtmHwhWyoMGA+WZit/LIUjf2v/eLmv9BEP3S9/g
ndiNWtMsJDucF1PhoWWCw24/TUbCiOauD9mlTSUlW863RAZeTZczUReZQoJB
M9LW3XROe/3Of8ZNiHw4ZnzJtN5biQbVqHwAwKGe0lLgJ4ze276IKe9Zwx54
4EqcUjUIdq+hIVBYG9HmrSDeAVcnWUcfhPFU2NnHLwUrO0Ga8Ph8zW5X/JQE
3z2iIz+WahMuol0olMjJdUzKJVAZ1RxoJjnGKV+ZSK5Di361C3AeD3nWrC+E
651Kq8mLSiq6TBzdQHkD0uHK/kg9onl2CwmX8AoiUMQyd49G/V8lP1KQa1uW
F1esUGSoeVY54KVi/5KCJH8pFgGne++UCtK1Y1lxjHgjdzpKlrHdcQSnBH1Q
u/KZs0GmusIprnjLXJ8+UBbMOPEAvp1B5CKnM2vULHtQZX9BIHTGX2IZNrpw
oqZg9wSiAXE5gkxt2CI7WsXf8MoztUrfb2bO/vXExK5fpawSTo7rCsFw9gjP
GcSxaHT0I2/0LP6fELtA4hPfyUT2cpiaNzRANW8cRSFhBNnoptmVx4hJGVem
DUN9wKgwkudg1Pw3ARgbw7Zu3SEwkvnuqXahxaPdxwfSQ2X1PukEB11wYsDt
L9LvMmeCNlwRqkFitpFKLeIUFAXUUZI2qcNS+Zojj/JuMiMVwnLCGf0QODyY
FdBv2QwjPZ4BMZaivqoJNmIC/FVM2BrkbmD+Fw2YtTt+r9nmmCXvWsuhOJW8
2T1DRCshgmwRbNxXkKv1Jsf5lzc/IWEMispsdVh2JKfPaZNeRFrluI9lnaba
t+ArVEH91iKMcoxKbYKItvpy9PwncSxXpXsH+ahnbKt+iSnqKXxzHXznEpFB
q6Z/7z7joOk27ddXxQ8RuCjQHtU4MzY4mcFipI150psuvThAVgKCEp55XqqC
v29RbeR+vKkpkctzKCokKANLnHCVszkrwTcQiitY/IFXllcR032t7baCN8cu
gHpJpgW2e+ax+8BQ7vMfS/2KzzGGqUWrTp1pK4EYc23GgREvMhCXb1+2XaEJ
3jtjlhkQSnxnRFMNqkA88qGJnIhmLlqtKwqZcmevRIDC5vJA0oV+2+ozsFlk
7OBJfYyJqPd01RdMQi1DFR19xDDk9JccWlNnpC/Tybdx3zxiX0M5m7QvGDGn
qWHQW3U8n185rM2ARZPQWgCos9LKCsqLuc1Z3t7wK4DwNCgHLb+/Na6QH1YW
HbMCIQW/t4WQvKiqJz/2qz0M4mg4rfaHqEzD0iW1WZxZsbY6yFCsWtbf5HXE
OOXzV+2h2J5TkMHjZJhLMhB/07v3LSmjI2Ip5qLHx0MLXhQ4Dv4LSOMA0/4d
W2DO4ISjiCGZjCu3LOrCa5/z2+w2Gt/P+wWvrxagGiDL5TxCvQ0vVEeZ37nB
1pkJr4LmAfHd4VMnm/M+YSIWr/6+qcQETYV8aTadlez2cyEsCojLF8LE0LWU
cT9ItDAE5sV46XmN1DnmIZFVamzDWI3FrbALjeKYCd04L7yRJX9jt3fycYDe
FkeDeiqYoUZIKNfW/TTjPMl7yVBEOzPkdNACvw9dtJq2NHeFtGrrBHIhEK5u
/QQF4E6TlcePDl0jDwZ5PR2dsGkVFcG+p0g9uop7YXRvEYqw3F1mw6xkZWLp
YNrFFJgtcWOIgFjNdlQZJ5qMLtZMpw1DtacnmAkgt0cKDPWoWKB5j9tYE523
nrB2N4NKIPyKXAyXwm/rdgoh6TvFgHs/Abx0DNJpNGGSZ/GcCqEm+EzHVySz
9AaIkvEpYhAFQWmJTNyno0lv/m7W0FZc1fWWtTRpoK+0lTpmZJxdpuzvVHIB
PomCb9YFLXsswnuYFsYWGvJWhSHZHp+3aoHNYSQb2LsKNUA2Ag35jm3jlSB1
UdCdz7yHsIEO0i3QmaH5vYgQlYAadMVtGSUapUeWI3qdp67x0pJXMUd5QAky
xpDqrCyCfMWJX358WK5VFO34R1CgBKFfem0L+k4bIpkRyd4fsuvDSY/Dq8yq
s1KQbutvUYPkoBLPJH1FOSr6e2v6yP5N7zGRAeDc3NgsvgK5j+x3fL7HWLrR
7sgwaV9yWvs4E1c34Va4qU/18cKWecKsE01QVPFI4lBm7B0Syz9c34l+gXfX
J4t5eSMjYUnCTWNgirja2Xy2G1R80OnXaPwAUIXFnFxJhUYcWFHP8mmvRG6r
eiE3e1GAZZ3xTa5P5glwIwxZWrdLZU0pTl5JjEiQS19ffX3WpIVnn9/HhOHe
pE0Z+hPOYAKaHqoGTuJKpeHrWUKVKQDxSgRDo0wl2I87aprpaYaE4aACqyxi
edF/j/ZTTqgIapli6Efv9C1iYMP1kZvk1vtxLTyv8vXqOi9ByrT6HnACByQF
Q00YHE3x3xxtQysmRDJkX35DrzoxW6KAsF50GvxGnxBTTUsPAC44hpcqVP9a
cJP7Sh20H8t/VCILhMYkeDCBByQhk1tiqbq8C60F7ako+DXoWrLiUeIZV4br
EThob5JQ0STTw0Kf/WHTiwpwqTRzZxuoM4DkFOATY/yxQTIC7sWVbVAqc54D
r9dZ0HJCh0SZdIDvNZLyBTgo1Ps+rsbt9k4p4T0IjPyQ/lY/XGQxpPeI7qv9
jiBZ0AwDkm2X3O4A6nC9PShL5cfRGH0f0bLuA/8TXIBCaWt8g6RNXeUnXRba
9VgoDC9BKHXbyzOUCgOiJ4kJ1ajfPtntvjJkwSY6vcTRcwPILfPzZcfAw6i2
cwEhGVETZ4K4B1/x6mCAD55+LqnwSxILER7L8LlmvXWUcXhHr/CWecywte+Q
uK/MbD+jRQqbvsaFG0WtyeDI0V86DxaBLn7BXooQv7PeDFjv8NpsktRZOaVo
ZltwfEWIXQgApRBa/B+k49BMTsfb042EvyCzmzf8J+WN4O9c7bsO516SDkSt
UTp8IZgmatS2637gRnFqLeF4MM0CRCYBhV8Fy3YdqjFqsZtr/hLJJqLAKAvy
LvUSah7GbT78nZtb7l8nlSYQFEMjILiBsI/Aaf6G8RQ3sStehU/uLg07RGtd
tZ+NuaSiN2MyCeEQdGpH+XqVPMD1iz/0rWTZN/uBbRGq++SYd3WHyw48SOj1
AY+H1shXJmKfrOXWCfaf8JxYBronmMSNrdOZNg+9wVE6skyjb+gs83vg1HZw
upcJXfEmRfsZ/gxt/bt0TMhA16BlsEuwKRDaFuhsfPL63LKSbEcGVCY1aCBF
vD4yT4e39CzHaZctjogd6/rZ2rBzdQ0SfHjRh33VdVDf85AhgkYCGo3c7C1N
SVcJg8Obl1+M6vFjA1S1KAP8y0U+pmIv0RjmFsUUTGeI2Z/00CS8jeBLylqI
M3phgjIy9ibksnAFIJ28JDYmoF3VVuoJgLUi2diVTQvii12PqwIOAiokhjsg
8UnwwVA+dQlr834b2fsW7afW9cA3DGivVQ6Pch3PRiJry9nMrL9untKCiBtk
woMVe+xl3wALG/tTn04s/KFndynFWlw1DCfYoITyctD1yyf9vj/MFCuicVUe
pR6g72cqp5BDPv6dV+OoXn5dwUC4Fug2lqyFrHo+nSWztaW1TDsFxqZPu+Wc
Y/f1OTfmx0w+nvP2eMkDh9J8yPVWVV9zOGbSUNzlVlbjjEEau3kVjpJvYQzM
cC4jQFuV4ZsZdFom7zW/E1hTL0fOeBB1PJvsV2fwVwzhO6iU+yCM6BLO8hmR
oLX5nme8jdwTOAjtBOoyPPrJUXw72fOLKyk3N1cgJPNGXUMQWt2OfOKvQ4YQ
S8kCAakiu0pBuc2myfCF2RjRCOB5QDbE6Urdo7m2iHkJeWkhqOR4E8MguDHU
12ArNxsP58Z1yRmBRDbTZUU9NDrd2iIiBsCVTS1kQPFy6P8HYsmZryVbSC93
QUTtNg4PSm2l2h+upiYG8aSrR3mPzUM0UTmFuc6cQoMtgw2GSp+c47tlA4HN
mEln+RZW/DjYExRS9UF/zHPUJRh50Zt4QVq5QDgykxWBsX2RynWhftsz9knH
ibEP1aXg3aDQbDgrr5I+ESlWKIS5IOiDmg9lh2ml+mY5lvrWpLsO8VAAmhbM
+9Jkw35mC4Ko9S3n2GFjUAOULIjB7UEMx6txrXX4aNfe7LvCSVWqt3OcdtUA
i7Pq0l6Gr7sdZ3X0RXFbjhvGIDMC6KB3xj7o7OOC3t1ySfXhIahtMnEVG+JI
egzkX1ZBf7gWNqIYvTHuRdA/EYqybfh5QYkzBZqNFxOGqHaXZskf5phCI6AT
FY+kOBm8pOH5dtE5bPWLQeWiOYk5b6XV/SThoYrnFoMk9FVzuMaloWTcUX/s
5OBKooa418NNe98C61l/LBdscpUhu0537dHFGhRUS7L15o06ghKVo4/6QHGQ
9zBkt0KxGudBf2/ywOMCojnR4EgHfKFSBbV4G0Wh6q6ID8UnXdf+ZA2Lj6lO
jeQvLblSa6x+gY8U5KDPCsXH00EVRWXEh0ug8G6HCMZolP24+jDRhZgqyQRu
1Av6F2TnFXzKBJDu6v1pgAnkimtHGT1fPSn0qM3TyKfthjQzgVQD5dzOoBOb
8nQBVQKnUnrLHGBPKq59317i424vyfPpP6caQ0tO7l9f4zPz+YEeUY32ebM2
VXPv7E6Ug1ofkkVMu+VruzkdG5Wi/wubH1JO/wvAWn/Kyd9BuGn0mOjRdq9c
X2MSTyksouqHqiiJafDQnnEH3PGZ82hPzLlws2/HbbESC0Y7OFVruytph688
9NGWAj8c4kkhgk26JcetC974leCIcTDDcRxKuZOfWjFAYiYowCyp55WTGAih
NMw3YpP1fLoKI5qdF+nofXl0Buqdi7xg3OBYJl9sZlrqUnhREhtowkti7J5D
2ZVJKBX5MR1PMH5zg9bNerQsFzqO/mZrO2xmb/WJDHuvlONONa0uSfbPoRQN
9WEZSszKUbbNjnukdGwV65ngVEKkG+80iyVLRff2ws801BEK4l2DsWnp3tns
FT8Y8NZLqZNpFgSxSxOnbD8BPuzdfCY0mm6459YLW1i4bHbQINWU+Hh3aLGn
DPl0TcKLI485ciDYl0sMGfg9yCA7tthagLrXJwK4Rzk2L6KKobzET3llfj+3
uFVayM2GJwS6KGpIpCTRvkoTzNihOcwIoS3UZ+B4e8dAuO+pxnCr0l5QacUe
/WoVIyooISrqISQ4cOPPRMvG7+c6h+1zC4npEqT6ByiJ6Ofx8sgZuLtZl2TO
6DeCEo+dRoF/frLQmxBA6Bi4hhbzfuo0QIP194gSnx7JeqnnFQxllsM9mZG0
xAHBKAyJliiFSmscjCVDS6GkIO9NqTv1KKjlM5/tZYB3MG4fSkVAYwA4FYhA
WXuOPAqHsPJU7qYUORE8rRtecHtfbPTu8r9lFKcSDZWRC4QWvYU9pXs5RPB8
n27EkSD2USyzX74XOYvy3kY4IeCih30XjPqQiIkEC08fpbPchjMgUN7l6q87
SHbc8i7uOMJfWTF9L995jynNoZMJqW2Jey39xnso5JWtthXHaz9n5sZV7z5Y
9KimNtzq6t7XEMBsYwly6tMV0bzLPZC+ko4O82KKTFWZoID7XZjCiw70MKG9
Fmue9fDdYu7g5aeoCc0RensrbBHmWPSGpgrSCje95FZhUol/cA7RSjGfgrDO
1VEch66wvN8/Ld0OM1UDL7CirfDPFGxozacEm/jTH5iLhkWqXc69XU+IUAtR
RucNlM/kgELQDM4uPUIhyiPPV06jZSUffbihP7LD1C7T4+lJpzFyWLWZPtIJ
GnBqLtMnW+UGd+uTn5Y5DjN1/diEsi1xTGPiw0nIijwgIFEHgkMZWZPzCeMC
2quClhPq1eQLnerY+bivjVDg7bLVMAO3PzPc0X5lgafGUiwfE35bpPUNAZ5a
nDgu0HyWuEm7/QbMaDCpXQKwvuTEz5tRzSgdy27Al8QQchpuD7WXlfw2Cke7
8XQG4XsrdKR1hizHrRmlJn+EfcGa2YW3YgKsXla4usIUdCXDQjdqpCj83WX7
DBFC5P/F4jNZTUm9AiImTbxc1l22P5NVzODM0rccc9pKZTK583MeZ2WTv5i8
JKXbyuNqbmqWyiHtGqfbTatMGtHIHZqtv7Nq8z+1fDxtTJuK6BzRcsmGO6UC
ec1dB0XcbJZbUNzT1pZ+70EEzzOsPMDclLXFOhfEZ95cdfQO6huvQqGuHn34
AxZdTCJv1n1Ktw4s1tNXiBqDi24vAKbIJW+Tp7um5M9gWq0GhFPC+yDsW6dU
Hew2WtX3QD4MDEXfRx6yfZ4bIL/vDGMNSG3cJTNEiyRB0xRCAYmaVoWnlV0G
3wXgp0kKRaKA1c5OSpIKbj/SEG5CPdDmRRyvEK+7GISmnVvFykHCcfil7eBn
/f8uwTLah85KfBJovA6EBE+dStv1ZG2fsJPhPE7FLG6IcNzJyFtKUYpnPNYe
YmI/NX/0WFSs1D+rxANer0xCDqXon2mvtiEuW3yv75QMupKqBizQX9J+PP7d
d1j5mZ/vRa+YUJoMhKbLHUSY6NVqt89veu388Apr43aY/7w4EoGbSKlqPahe
zNNpBqxKjz+Ik0FjzA7u08hFzhC+aVwT3DzUDxLYjX6PCNNXR9Ky7GGZlnMT
zaYw1ZRYSpJhW7lu1LVsKpauzbdonPXVrMZUje1nwcbxRY+SJkW1Di9QrcP/
Ij/q9RZty3luP9HRcGdmi8lBvPvTc7/+gzzbp/o7yYrW+x0n1e2zE/LS4CtN
gp9GaBItAmdud8Bad04K6j12VTYDQFkvV0U/Uxt+gh2WpaUuiZ6wFN2l7uRl
Tfh47Zl+jHh45uxG3Cc0fYD+ETLXYq6L4xFMJ+e/4jGyRkwkzP5Xe2th2n4U
+oeBvXmxYnPEqYdD+gfErvFyZyjaWQ1n4GYEEff/pqeLKxXKobL6z4zl85La
UOlehigehHP8KzF6UHzUzUpMQgFTdseKtVD1MTByGqRHRr4WfCEeGSGoQau8
w8nzsjeYt4ScedY2U1c2b4RgQj9To2YeL2I3tw6Re51sil4rUM0hFgO9aw7l
DP3v7oP1zk3GaFSRCO3UgKFOLjOZV6uBP7dhsWZGMur6cP9woaotXLkVXGk5
2IeWmrBWQCVKIn+R2iTxoL3e6LS4ElOydazVkM9xiRH4+/7TgiNb3wYwwoMG
CeDaa4GnM/VEoiD9Tl1aAMOJCNx37QaNqDvIbWFnEr3tiC3IjOpv8HgsOx7P
Auc43A2WqInuJd1FqQ9kH9i4akc2sYslJncJqVm2CWBwvRT2jWnc7vR24+d/
h2reHXOBXwuToj5viV7yoeFNI6duB5/iInPeOeJuAsl2V7hcrpW/b8lMbzUH
fcVF2yi1Z+UYMcUiXP3mM7YaTX8YVF4GVQ9I5j0KmJuJm9Qe7rXF9M/nd8R9
OO90jD3rvQuSiDg8vbQofxKRQH0Gfq6lhx7Fm5fpuc3gtTuqstmXfr76Q7wQ
dSNJw8ql+GySbeJWA9xeKZ6JifrsANl+4yr75rcoHHQb4vpAkcxVT2RGjoJF
gV+fWJ3SvJme0iMlna7iEx647kiu3LLPqWLTVm58uXnBRyfZiMD/WL4c+zOK
Qm+IPP3TxElBbZwrGWw0RsN3S+BLMqEgFz5ueycaW0/WhKFGlR1uNvkde4Ym
SGgGe/zoPgIW80SwulMbBPZH3AaZxlXgF18fupcWuBQa5j7HMqwtmS+sEk6+
tXQE5dpddz+EDCwUB0gn9VFSULpkJUT4hDfc0A3Qs1RXGH8heRj+2UNpgWem
AAh5vR1SAnjMqckdtQTlM3ViAY7ooTF7wZQmwFa0pTwfYQGb2aUnd4/iytbc
D3aiBkKY/QV5SdmpActAZEF23HDlwu/rs0/5bFRwaHDEcNsz8J66WIXt/kbX
hyQGNWF8NOAA3iEKvpvLO5JB/NZOXmDNcdWfXvpVnAEoiVvCVMuQ+avDfMhT
EtoNiaygtjQfCIW2sapmARgPlG/wMR9UuzIGpDcwRcKQMEuCUtk6suF5jMor
QR2oquH2LMOmHCEZnWLwUi/gAy+82g0PwSfb9l54lQOzunEDd+LQoqI9hKkh
9DlJBXyo8jL/36a8MqqU/n/SG0uZQ2vHGnU5YnTsMg+JCXELcsljSJpghUyF
q8jqla6v0CroeFj7XAbKIfl9FKJUxYp/FB6mj8tWWftIxk8u+gJnNfmh5qqB
CtsUtq00Zd9sAlFn0oBWfz7/yGdwkTWv+ERgy4v5dUnSoHju+W5xZT6Mtujq
Eycby1ZfDjYQnAjy2Svc+geJTgbyz7Jo4wPgj0YDREYlNZV1WvL8K9ls4YER
cZEIiTE0m8vqxU17k/VrdbBWEV7wLLtnVdLgd4Ul1/Llolou8QsSUMeWL54G
jBjyG1GB70HG4vOoXR7rfJDE9u7HHIlrMhUAjPSTyH7spn/jtXtAqRyuo2kE
3uKN8CckXESkX+iZB5BwEtl5XcDjQWBNcBTXSgfeFYOp05Au9givOFZoxc5C
B21aQIVKbXHneZutMN/c8zUioVmi2Uu0EW95oqT6zqqyA237Ap31WDH4liC7
NMN1CYEhvkLIBlHcbslBFHGCpmGpogvYCAzmG+XRP0kIR3QpwlkjBtNEm8IX
z3aTdOD5QbVu7OdcoIs7j1WRFuPitzO1Ha08Wv8xuRA7SdmPRAYJmWjHYLsw
yeYDVkoC4dAfYJaCN1AovKv2YlmLSHp4aimNdJxSMEkWbqCYnRPePP3gsbMy
JQopHQ2XEtZQoBRZyQNWSK7D5+uS0NVCV/LGDpjKK3NPjmcG+Ft1PrGxl1TI
pb9dyv5LFhXf7NAUVv+3XI3V4ztlIBvKobwxulXXGsEr/lH5oi6aSgkY3tif
5N2NkCh+P8gFHG96nlsXCwCZHjvwJKVI0k42d/39D2bFQ6tbk0FfJ8/N1kG7
2ehg/XFXxE3iBaYlaUMQjkUJmJcJTHWYYGQQt2V7r6VkYs/5SQ3fV5ynIrMS
rvAJJPE+QyV5G/W4bq/Lp6WjaHp22md9k1O2A7m4iy2fEeISu68fScoDtumg
O496btovniNFkqUky/gpBTXK0h+lEwFxAAXi4wnK8A2OyVSSBEqaM8rUStAK
sl3gbgUkrtwWLzRepozYWKLr7HHJRMH1LAdu+aRdmLPr9IYug9SqT+DoYI4H
PIQvWABopcPZwQRWB8nDK3NCSrJMK0ZnE6db5FdiipDnhr4HOEOYDWV2wIJB
SN4zhY7YytDxhwdlpl2FmA4EZRNWCOfM2a416RVF9k3Lfj2mQpil/7gLa36m
edRlAXdHtYN7mXymoLGF4d5k4Lf7McMX4scAFbB8CMWDv5LshDyIFhuhCZBO
vuYttPfs1LT/+aZN5ZxUHdt/jGwAnTpfdPmy7U+6Q4yDpphi1s78fA8Mbo1s
511jQnMCQIn30dXv7pT+kdEq2bjM9dStxVFdLv6jS0mWEf5bGqs20UcKMI6S
zGhWHndSvGdMcA8bT0bfSgwymoNtsCElX2RsY6194MMNVsjP2sgf9bx1opMt
RLcS1GsNsMv2eUD9LQSO9udRXBOi8vefaaR+EUQ06PuhEyTUBm1lnZ68tTG+
ajQJh1apLyrHzlpJJCH4MK6z99QyYToXRvANWJIWbKojRbWM593QavGhaV38
JK3xhhn8QFvPIshSvXUSvsTr37oVpAALD2r8ccN/pM240elVMvsclifs/I6R
Izkkt2BBPluhorOCj1yMGo1le6iRUywfQszPhUrJPyfeAcXYucL87EFNcf8P
99reZEGL0BbDYNgES3eWyNS3Km7HWVRwMN6vlh1bM9keWGA4KimGuMkeotd3
4DzKIizZQQrEYOPXNWKkvgFWhLVwW3mYyMtMFCpaeZZBKIMgJeAyQHaj5hzE
OJfCMUu0vl18gjcEbDaYlPIfwkeE2GJ+eg405XaWCND/7YGox0pdTAAPVIKl
5rcnXDOW16lIEUkxJyeXOe97MVqKNsS33j8oUEnl+qqjlPeVn8L7XXrxp6rW
Fl+9c875Z3FDG/VGT2vkALxJIemU39e7XTVVnu1WTk3kv+5n90c2tmhHq88A
+vF3ASCdcDDjNBt/rVrM9hNK3H85qgt8Elp1tFVF5Hx8KGFBG1ZohZUUggVh
dfY0HBjxS+txYbN1Hcv7KM+qeXngqdSX6yf7nxNgAAuXkAfKGVrRXtFgKu+u
WT1Gt2Gp479OBWzHpYwkWMPoDr763fvmC2gk6KTyFwdslQdFWuxq1vT2GcX4
jhzEzEDDgSYL1U9e/gw+FNa/fjXu4Txqj6htjyFrsOPpI9mNKhWtDfS6aHyw
7RI/ug7b6etzsvTSeFUsaAuqCG8JNKp4T7gHPqFi7w+UVuu/QJUwdchf80/N
12QYfK9GARe7D4hd6dgsRDnCOR9L+BSsiqLui0gCcv5EPSeMGCMHPldwdDUZ
7A8IQXNKYN69Eh83bIBaViHd5Yq7viktXKN0hMlyd9hEjkGXNNw0AC7rKjIy
MlO//UkVHBNkG12W/h27wi4FfdFGkspZl2mIxTh3kiRfQwjcB2g/ihvViPVN
bpVjx15NSDjTEEYsQTqPOmN9/TPptoe/uMOxFcjJDH90HSFkPlhO3zZcXItJ
yxO2XxsjikJ7wEXIYF/KEVEWM/jBBhKq6xAsdFdtd72Xk2xXFm889gSpMHxR
Xbw92Bg/NSZjYMp53hqmXfO7Dxmijcp7I+cX2yzY8GvzvIr619eqx9MnUP/2
UeTs04bBfgi+q2Nw8ryaQHQHuqltPfyWsA6PgTOY3rUta6PW6b1SDEzU8jmN
1Mk6oehReP3YEsUXdCaImTm+WI03UXzPIbU3CzXbGvmvKjprfG+yd7DZM6Gz
0fyxjd7ywgWSG+mi6n4GAUFaq9VK5PkPE9GB21rnIg+C0DZMpgWjwh/NvgC3
LvOJa1VHEbg42fBD3sQn4rfs2nj4K3ZdPcoKRzgpIfVxnC4rOJwAm5IzbkRW
9YqWV/o+iz5yNt+Iwk1f1vRp9+gDnca1afzFae+tCdI7BVGQbll2lECJkJwl
hiR4h0jpGebsgefDulXDxVzrM8usxEgPhetwX65NSpMB8C+YvwUPnnVXnXDD
sL4DOeKh67ABFrjbzJwjlmvKEyZoBBKigI3mQs7IO8eplTdhGoEFY/ov7I32
9WjE7j5Q9G4wv8ZI4Txf9+/Y5IgM2aLCTVHGE26/VhBG0P7dTgE44lbkrrnJ
ryXLoGDHVkwIuJCwCItMtPifTPV4nFqeSzJyWwEbI7B6za78fJAVKmBFGfN2
p1MA8HpKZXU8WV7MuSXcqSICtAq1HLHWlgnLJ/Jigk7dQ0XV30jt2QYdV6RG
IyzrGPnKa+UqatxuTGmGIJ3oO5zaMkUEYY+pjBeyArVRI6I4yDkViCufeBJ9
LIIxbfCLYX1oroP14NWksWUWkxAolcyBeCVpT8GpsqEN/Boe2jFO6GSD+7wc
aA1qXuwsqAQ19a8w1FBlb0MsuYR1Hlro2TLS8eALhp03xFliVLjst6fZftOk
JrosWfkCczm/fr5HaD5d86FVT9EFykFfqo9AOKSk6+/1ueJkVUUWvjqFtfri
jFQz4K0Nek4e/P2uZlRtLmQKCc3pSGoklOzwRMQZ72niGfvd1f0rOy7PJrQo
s6aDdgqBzAo56WFF69BZTrYAuoXqQXE4PQXPQPdB1HSis9hW8z642YHYvrq/
DTl7DrrJY8lzIvZctuCko1S4IQPpmOHl2ew8std7qBe5VBk73cfAgzHdk+PQ
t+YiL2uDU+nQVp/p+/Jz5EjqWmNxN42Kfsyq2QxeCoo5kQJ/PbZ9mF6HEDam
6JBPMcqAfyY4VDL+JgoC4s9KQUMgvk7/tzDGEeZjLGEn2SdNJX1x0DujYnZO
BkmDHVl/+tLY4Qxt6zCngqGuOyXcV75uz4GowMWQypfk+BYEYbDTHvN78pZ+
lM76GIEu2cIZeE2twRWHzFmRRz1bcbmGOt9o49UD4V++5rmXfwsi7WTEp2bH
KMSWy0fwAXzZ/mvX5zz+1MEeJ6f8EjA32kmq2oj+hAoabg86miZTEDBvruC0
EVAPWFWOPbJ8uYeVHVw12hi3DH08dHZs/6PJfI/V+5giPGy+9oLkpe1bk2mW
undT3aUJnIqkZHjXzEXXVbuB41i5kfnEg7h4uhcoLnCegC7pOwrwRIgPqaio
XuthVG+U6PVFFVO5Rd1Ziq1EGIPDBBbtU8B2U9m724DZPxluIPjwjvefFcz5
fwAgiQ9hRC4H7Bhexk14lRTfW4NGLGZ97SeHxmzq+pKbctS+JOLQFTuNh9So
m9gPbaeZQF50JrA9NJtqflnyulFy+LviltMAFpFXocA+/CxvAr5ayA941tuc
jv8DvZ9JXljL8BlgOyIarutKBJRh9kkg7/FT4nAziCuwkHKhNVnSwW+LbQ8f
X0r4TBmTToaDQA7T3uyGtZvPr6QnCZ/3YrVI+HICQ695wrtrjsRGrpKHfklD
KpswgkkHwoIjGFeLhgA9tqeiKCAkfKgDnJMPHHwHArGOTM17A+f6cRx5esB0
qSCmTNAfqo7H5Uy3TpjiIYPP+MyRncNWNTD+7cXMINhHAtgt2TTmVz0yKTU6
3haUi4U/0+5HyELDvQ8Nx8V7JbbqvE9A36qCN/9US2kH4zMx5ZrrneNbcYLV
TElppUmhIfRiKltM7GINdO+2fghmLwWIs0wPaeuVOXo0c1SZNu5pY/tWOoeG
4r8yKtU+oSiopcXmmRlCPZAnbkuruPzGnl0HBY/89lRM35RxE2ftIWKyVw4U
F1zzI3efZS0q8vNUIfMp45/8vPYoW4+MK/jksfWtkvN76nEoGU3K57R9HLRj
bofqeXV+L+k/IRLI+lqoWBb2Dq/3Bf4lvOLGRfu7Ad57ZHNV4XG5Pr+L+K2N
3CFiQztEJWq5jFYhdvn+gQRrQBD7e3QG0qFj/lkpYbwVAKF4IiUrf+Voc+sW
PA/uPRmtow1bVfgseEM0se2nof2c71SECVtTJp2FhhbowWcdGEQNeneXoCFE
Vp5ld3rRpARYMQXA0aYbVxXG0xohKEmqHlVBDju5JEQF8NGYjCI4R/lGW8Ni
NxCMaGMfJP93jSJgK5zrvzem27lxEItpqIbZ5gX8gsHK98M2/xHTUp5EgqSI
u4QYt0P+30oROTJvGrxmsIqcQ4W8+k08aEpa79Qf/KLE0UEv9m9M0oWRqmIA
9r3ftrtbo45xl24wa+IHog9MYzq74+iNhlkbMh5hPC0mfcKGOHNYXRo7Vr+p
7UCMqrYzBDdPqyu7JohHLTeXzyC1cP267c46Jo2ef204siv7tnb+RCTuirGY
IRmFIWkijQLt6M/CAzgdu/eDVk47IQFio9OmtSRhAT39WkjHiHZZwUZ7QK+j
o7n+MZu9XJNbTvYSbsNld2inhUlPmv8Y07aOpbYj3S2z+Ch+MSAPF4o0GUL/
ykVcps+IFv272ftqCCX8ReKQvK0r45K+l/N5G6KAYuYM0PptTchh4z7RkLwD
/5jA2+xbkLTW3WlogEqVtRfpiinAY1j2uvsjKwVgJLxO63baUG5ecucELgDP
LJTbMq8pBkcU2ff4CTGnGO8q9tt8pZ+h+i0sWhi4CJ6XmndPJQvFRLWXb5V8
felrNTMnipTHLp/VSANISdiZPQeKOQmUF6RMGdbgAApahctRg/fWj+HCVXOA
alcWqZ65ZxeqFqrWmNYigYawgqtYd4h/X5yiVmi2L10oiYVbm0/6geER8uPo
NbaXFGS9+XrDO+01SJjKn7nfyraE7Z7NhkjGrxMFCviW58ybzPoSK635wJXm
udGgGBqTgYX2KpUThsCDsbXUOqfdVtf9RcWRHjfqrUEQOa/9XXi2hAdYvP8H
G+q6t7SXj0awRjq+QEVYPbBeLnoJFIn4z0UyBPqy1C59bk5BjvlV/wzeHE90
zaXAzpB1aL+j8Vq8PyLq5076dgwPVh7MdBH3LDkTTo6xnH33QsEGKS1CGabU
6J/oWKzXJIxOSSZL1Z4UZf7TquGit1wVKBQKQLZCxodeS92X+Q+xfrv3jG9D
XgAbj5zBYkFJJ7ak0ZWlHJKV+UJeAvS6zrexBBLHk907R9Ss5x5o3ZkFSsmO
5fDMk8rHGsSKQ7mOJkho4e3e+6KkDr0KqnVqBGnsY/MKy5gEVNRKxoTlJeuq
Ov1hwayjTSI8L1ckDxFxyW68U9754T16xMwCjK4stBOkbQ+1wNnqDHAZjHtS
wM551KwOsO+2ro6ozJU6X/KYCQupo6+WWxsGLruCQvJXX5Z8A7CYkT7f9BsZ
hVEylZDNqUvzAe824zB0UewUYNS/L0o6tSO8ziNbwtdIRdlYancConJXb/q7
YTOuq+M62SgQk/EvTRFeZ7mIexy4qCKgjYYAAZa/yYwobCPT0L2iGueRTbI7
O5o0BM3ZpITdrepE1Ou2IIAVm67h8iws+NF2jU38vZlRCo+XXUx8fHtaQVEE
FG4lLY1CujfZwxzXOj/O4adXvCBPesQ497+zN8yNa1z3RUehj9ivI57dmmZ/
j1fY8sHtHeRGFq/z6l5z4F8oTudmWoMMqw1eouaZ5XKrfS6DhW0dG++Vr64F
73WVGGbWWPXXWwifD/cjZ6rN4F3zyylR9nTxlaciLZYjUldpk6+OWCXZ8iQc
NaRWuS59japnIdCddWYzxBdrxXamq2Nx1NVMCd+/iAslNvjiDBE49zCyQ7d9
1X/4sLsNeqqO018YwI7zXE4P7Vpj25JFJl3MhE8bu3GulsA3lCZiaN9wtxpz
lvImLD6BpKP/ZisaKedS4748Tt5whEDdEnI6afxaxtNZmAK9ke9WEKocaJKT
nXhBA+nPoKVYf/sryjWcBX3yIRJxxWXQCwzzLZLuv4gEUCBAqk0xVodEDYCe
WqznLmC4UV4gqJjuiNJC8FGA9LyiynZkro+yE9YtAxGZpt+8vpX3od0e1uLN
aioSDr2yy4YG9GnHixb2DFK97HgjhwI4saseBq0yvc5WthARtyYznQi3dD0Y
OCuysC6qYC7Nr6RCHXkT+cg41jleNUhF3t2UUAl401DMbRTxaD1bAd9dYLjG
IpDPCEBTz92/XSSplSP/qm2IvSRCu0ZD8R66vJfTRhybIj+ndNHD88MnLyqn
G/Dp+CD4E3CpJvCcnMp1WH8Qsf9FWuMm9Ggu/ZSBEu39rcxxX44QsJ04dRTa
LjJZT3FFmwvJgBDoXt0ui+iSSbd/djj+/ZMmSlrScY6UCUv8JtyylXr7kYZt
Ncgz5Uvc+arxJmmM6WtUc/QyDl0Fhhw0mhYvFGaVx7rfi2arYZPu74YkFYUf
mhrkH23fJSCVGN/LQ++rFeSp81qD7JYk8jtt1v+ZvP12/Sz8qQhdGQp/lq/r
p9ZkGnszxBhmOJoeKEfFMVia5LcAhPyTwMfsIVluB2jTVRffd77JrMsb6cHs
74C4JXY7cqaC3EEot69fc9MmWkHd7mtSLLPdceafNanGsQBqUKGNJRX2bpsM
VtmgYrw33no1Vt0fCKPxBaKZbz3gA3ioC+xGnlinElzanf8KFPYAq+I/Lmro
AxwiWX7oiJVU/w0ThMwB8N6MLFCL426sbEhh3TmChwmF8nlZyRarkDa2R1A9
C+rtF8+L3XLqW8xDnUjjiII/kI9z1ZpYRpHhtR/euX2YFXGunaMh4C+n3bOs
vTfwM7DptskTVe5pShE7qvojgQm1Y3boSLid5QA7AwJ0G/sDhSGOYukIY8QO
fCz+BqHrgMHPKvCecSjfoKpDKSq7wHqxMlCa48P0fsN3QLK9WzGzVF8i4evf
Vs69g8cRk8vikEM2SlrE2syDdNROoGus61onT/ZSDIAcjKA0UhoVvri52hc/
wwxHuG2lJ6flzfJMBcitNfs6P8aO2KxzqMJe8vr7G6uWT/gYzBBlz4INGvFQ
RHwdtxU7SLDgukVIZcQxRzimuJ0yPHTXuroEct7/IuiOIvYcKPgIIKkgq6sB
xBmXlb4jX1RRhjprCbVwDAWFYPbrthFbhN3sCvnZI3A+KVvyFYUSFSa9HUs3
xAde6jP1kHEX7ghCvSf+ij/XDhFxRdzOPRD2ySQpSsZso8/FPmdq/2YiMWub
SsY5lnP3ReCLSaIFG84bO+RCm+LdtSvPjQ57tU5XvuzhIidy9FWHdmqLLHr4
2hqcjEYGUzqsoR9cPxcsFELbWySJtEhV+QI5821sC7R/NjLetHUyGk3IW9wk
M2LsdEdKAB/52pbTgECKjg5JS+njzhMWEdSqacgJFPlT9lCGCSFl70PxkCLI
PpsjbcYyn5i/GF06Q7CzBO8zQhCxJhoLfi0Tp4I6nbvxatzFU8wPG5KqfwJj
ox/3GwnrgCz24IH1b8yUIgleWBUd5+fCSdm/FMg3GEf6eytswnkOLfpRasct
9iQGq402V8/p4V/3wpvtRvOoQrfjl/rpoZVpieklWimm4iXF1kaFPf/ub+Ay
8k2lF2EedGrg8iRyJOES3zcvbQis+7OTY49+mMZwsXCjDqIfnfaa3VtGHUhn
SkZjYRhK/ZevAnfnmn84oTMxqLOcU0ovL9BWf2KhTDYbeDSDC4rTysajnxA3
A+rQLFGBQO7tViyU1mIkNfUl+t1QddLdqWG96aQAKoE2R2VnL30D9q2nayth
F9YwDOwH2/dDrzryi6AyPIeFmOH0xVpH3cGeaw6sPDZ/cYIWZWVnknE0e79T
ZDoTpCd8cod7AuLEi17RKdZ3jHqh7pSE7OqMkR/QdaAqblvtqoVmxURqikz2
FWpyUpMXfh5F0E8i9rPc3ACPzqq1zDQji6U+zrzZIPtfhPF1I5LOM/3TOhUs
9IjoL+HhdI3xr4TJNka9EsrLZB1hhgIEoDVyV1XIk0yhyzXCqWEfACbi1h8f
xxkmtxUfkHhRwCtrjaoEuG/juXl+t7v4W6y+OC1+tlJ+ewUvC6sjnD0GxkpJ
wISqjVD9HiYLljsHYnPWscgRIiefKTTKm6TG/g52VmZjJomF7NsXRWB+8pFc
sS2jv3/OvUEXAVOV46hcr6jamM3JOUZhiswIAmPHwupXX2n4nl1tMwODdsBZ
yTTNp6HAdwR4AvE6pDK/YuTky942XQzymCSHle8DmoHzRMYx+5Za1JBAcnGc
u53RQaEK4MSMyo04JA8RhBo9+uqYozx/r3zfDCcyfRvRgH1iJmewWjtQ7IUF
LemYPikiO9fIEgmZJSWGcqcg6BXaux+Nq6lwj79sHToLTEQej/C9Oc64PtJJ
Mp6A55JlPMIFou6WMFvPrFc4vnsjyl3cZOI9MRLkxRrUvd0oGbnLx/rB2uBG
CbCrQh0/eTWmN1I+gEN557p9Df2y5O9bxTzpH/Gqx9a2Dc8FAijapNH9b8xX
UISIlbUmCmOW0ZhAFtQpQ4ZIwAMUqO6EMnaAIRJVAHiNmXFGahoAZxX1R98Z
Jxh4AEa0eFC5X1VgGs2zcr4vmBRPSMVW0tfFImRZoqMvflbrhRx4hjAyd766
Ujp9p1JW2FZ6vXNDiTNe2O/aAWgtqNYB2YW1TFlJyxWUSB7hwzheGbaooPqv
VHL6zHa3L5u4T5oVHVTazENfcZu4dZINEq1XEZ27B6MKbAthbNP28ZeBlJOz
pW7mcpEMWmGzSijZTULTYfztcnd0VAVPEIXX0Y4+sYEedpGoszjNHb8BDgPw
/Uwp4vS87eGrlELedkS5nH3aaBbdNNw73p81bQOel9s/OfkJ+8UrJV2ic40o
Ph+5EMdvokaNF6wT4akLq51uxV11nO3ZBfMTWhXGjiO6zv/j/0ig1y4kAwpi
U9IXfndDtD5ZcPSkL/vDxujG5JJgGQ6+TVtBSXQCR6Bo5awu9XpwqqnfwqhR
sxnTmF9szAYQVwnerKBaSW+hi0VvsRNeyW4YOdp5BpxCvj29lK514aOLB6tj
309Dch/55L07REg5Tn6t7LkGXv79JC9C8Utl8pJ2VtB+pqisbV3lhfe8diHB
BH/cOj3aotP5o3ipgyZMyZcTD3+8TE3bp/+ZY5JyA+kSGH6SNo4k1EBSb9+p
Am/EC48hUHgulXgqwOqXP6sO6UclahkHgDUEFGE0/f6MGTj+d51Nee+dTxHw
I4fd6Ty34GGegbQhHI2J1c72Q6LPAWZqXxYppfw0NsY2g0veTxqm1UMCuhhC
hy7rgDpaHQzibTRFxrj5r6syFiGqUVZRsH/11Lhtr9RIb1+biHGP1Ma8BOav
GuP5lCByznUCmfzGjX32g8O3qw+sh4OMpDpj9T910ZzrIRlaaaYoPlVflUzU
oxUpSnXjjQ/TbGBGc8UNKfIh18Z/L4vVp3l2kRoZmUP472bIX7SE3pXe34gW
um5Kz3bWB9FMts3Nfz+bRA3kIuBQWpavbvu57uSWNxRAb0hrJrYa6lWHjYdx
1w67KAbmKA5fuskd2IaOYsrFbHbpP0Ej+ERLaCDxzkKDr+uJ9PlFV+Kpd281
73v65/ull2X3c5a3RRdDZickkpocOZii7W1LMUfY8NWwLkdzx6wxiJtwMVwO
e3+PS2SSTr4jUlZ+Niyr0IjTtVSkkzQ/YQKSI4Ce+MxA6mlTiRN5OGOj7y5V
nnd8vbpUErSzbxJS3zoJt/97tzjQQsZb57VJeySCDMtgFMBZSjUrMOX3FsaD
HJPVDfu1DLIBcYcR8xvZ+ilzcNZnIKI91eqBLwuVPY2vnffEmYngRTErZN6e
EngivT6e+aWCVBlQvglM33OkH0qvm7djNg5bLEZz/nFvuO2BnsfnYOsLZAoa
D8s/wLPPbE/w8PhAZRocE9RSUB0KUZlrYQNMnRW8BNePept4BNrsgsVA+7MY
aybC5U9xiior7YH4hHvL9bPVhi7jkaOnEDxIiOh8NIg30MxKF+YBJETyYIDJ
FSvj8WABqtr2EDJhuFEXn29RX4bEj6bz4N3q456WvSmr6FP02f/pNW5nhOwR
wjvnj4Xryorlv6PYSEyN0tUseQ/tIyCRDWEvob1/Osqjtai4SPRBJf2XUMdH
EHKWPCRHhRI19AP9oR0Ty97k2rrZNM7/4sYLylTicfl0uCpczG7rLB2G4aSE
jXlhhoV32AKHYC9eVfrhysVTz35pxNLzHSQrsThbRiSTko6+z6/yAikYlMOe
i5E6IYQdxuwKBvtfz+++o1hLl2g7E5mlSR8a4Mlnz2YVKObLKcsmDq1P0akx
ChSItHN4ueqEAdQANZtQKgNJMvsEovmVLezuEXI8X91nAKk10CkGpeqFoDsx
yY5dMzhwBzY5fU88cQ+kggUyUr0C4YPAKVniRK/Thk6sk7sOOFFN66C7ePvb
L8fUBYdLUKOkob0POkbBrpeniOc/bjdHhqGyPTG6Gdyly9VLP333801DqYyD
46D/leFtLs5eMOW9xYFKCeJm+BHTZ0P34oEU9y2jtyTivZ1W7LG1wbzmgy5R
k2dP9eLVJqlIda3Yqw4lyi/Bf7gNnIWb9uAdhoEtC/vmFvK+08qd7sAt78yZ
RzA64yR/9zhaJNZY9MbzRo9z9rnxQ9xW8wt/XSSF4yB9ukIT1LjwKMbyev7l
1ikwxL+wDb8+rSJB7XYUFVJX38vWu1gOlOHS2dVz69twWzgGbnKmIMUrjBLj
dameaCVnCzYvJz0Xvp/fHHScrKOKFvRXqkVTBDKIu/2xu6l54ozRDL3rUexR
boz1A02Fbya0P56PdrOuhyzFZauYXjMcniScxdvF924qSaoa3FvoK5C+ndFd
qIzKRq0HfbbyXobQwB+QLXto6t+CmIaeN6fRnUrnkDv4sn3/igiZ8v9Qxusg
jDDL3qtHfV84z+m+Aptax3KW5isEt9H6vCPB+Mn0x5ZQLLZw2crIk7wISSRi
wfBlxd4A7DXPS3Eoq8v7acZAAbjNBPJK0p2VFshBoS2s2B584gexN/BVRfFp
uMozboKRKhu0kju3ldUCaZRVZLNyVWxNNXzH4ZvGEIW689ZFzRJKVUvMhoGg
n97AJSij46r4mjN6vQLgM+i4UcdflZaMU7WQ92Hdu58+Us4jxbDv8yXCe2KI
SUVGo4XHSYqsj0FwInoZcN6jSw77Ig1jSyRlSExtqPDQsLKm8cbzw4kiYs3a
ZpbO8VzUGZMC679NGziDH1k4M7UTMj/wu3mPiWaMki3Zd3S97XBvQVsnjN0G
3sFW

`pragma protect end_protected
