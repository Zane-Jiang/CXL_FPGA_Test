// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cAcZzoZceTSyAwGFppcjGOFMGge8zRHThThnbRHua9KekMSV4mtoYUFNSUc1
FHrqlJoCWHgEcyXuRecymBusOkwzUAIZbEzINZy+SNuwsvbkSvu/d9Y3AaeC
WIFdfys4SHkC5k3AE+xrJ8h9C6FD+0d4JgCz8uPGBSl7edWFm52AA7ZzPWab
JxnVr1t3hEbp7iyuIOy5QkMQ+B++fX23snTm7sgPestHWmxwk6TeSBsQubMW
2X54nukCqykGdivuo+80bIC6+GI2ilDDF0iKptXSOigwd98IwyN1ZzPrQ6wP
2zBR7V3O48TkI0BSB2HxIJiZ2D8DR1YvoclIHrE0OA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
e8J8MzOcU4d68BwiJ50/b4gs3joB6RDZS+48uqgkydzrmUb0KpVxqI2rzz9Y
pJwVjsATLbB27gnQCzbrqXm75RNWXJs4PvdI5tVXNL57/CSpmgNJfjbw9ibc
KbHo8kbBE29jJo+WMkMAKL11bSswgHmJ205m0v4EHCM+iBQODO/No3t0Fxrc
WM0H683yCDFWvmUxaWBVnWF7Z8lKzB6WQzWS1GWv694rlfR0hn/edt4FUZmg
rJ7M2+GWJMNDReDBUH5CG93XbXL27dGReMBiN7R3cltNg80gaovgpure3u2E
+g9I2e6H+T0iMcg9XEloV8gsJHJoNu5fNFvFyBTPNg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NUJV79U/lmDnvD8En/6WcVpMWvmOOFk/tp/sSM9fVoBeBYBZWBZy3JBE6L9u
8eJ4+V3txbHRzF04qELn3UnsQljlxdZd7eYChooudc3J5bnv3pQ1pcUIO9RW
FppJ5GuvI9bE5xNfKulP/ZJUKIUpBNWf4/Mtr33DHHl3lvfak62rQTdKS0Rw
bRVbSu4kwOcs+ILwM/eGqipSlgJB4vLVTFW1Mb6BXfMoD1z5cJ/vst4WiqeX
MvuNKdS7ZpM/KsS8f7wPXk/ign2zQFMFdU7Rg/Z8H+EaDM7cOOZwofViDfzY
n2Vdg3STwRTF2qpwj/smGQQ8fgW24CiSyhh9jOUlGQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
naUu+L07mp3iIIfDAqDDr1cLmYHu9IwdYjfle4NjlNAUTcuIxtNj7dCl1ytL
ZiAiCrvSIPjoYXB7T85g9sIAEpUYT1nS5E7cNILGQTn1tyR+JjkWZFUPxUto
/GEZDF/5mcfeC2B+P096wHKPAzWapRQo4CwXL+P4A9ryV9txkPA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
X/MC3H61pUTSBCxAO0wqK7PXIas4XGbiu7WON0aQ7md6tJQJf3fTN/7m0wCl
PiYTAn/CDLFX9OXclNx7sryOqv6KVQYMYswB0bj2gd01hvJ1hWZTbCtjpDhj
4OTf6tLyDAgp9HCJJQdaTHVlStdNH3SQ2QWmHj7X3BgZ5sEXcRmPfkz6ZHXi
5BSeYSw0VDLvtDoeiDivp/z4bWUBPI+MbCHAQdHa+daaiYZyTnP9O5/o13fq
NSTBwxQUYL0TSfI1FzW1iGhaUG59G6d//miTT3zmEcNsm3q/BRg3h2EjCRXB
Lhv43LC38mFBn/1/8o4UhrvPSQ7h2JYAkWUm/vU2rGund4RCrdVqOT1sVBTY
llkzBwxMcmxmhFT7VC4G7eKQKlSdBx/GwNVvxwVgEGKYvfeIVqfSzbYg/QFz
K25wp6fieusXPUnkLy6QijmlhONg2KF+m+pqpzGs4kEjNSKJegYGrcM7Txrw
/nexkTmZA0fecdQa/2Wa3V8/ld6+o+CG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iKuvq41uHLvdntGPwgQ7KJvijBSkCc1IekkztqKQt0V4Q2Y5Dnbdpn7vrnXI
m0gzFzDlI2pn7BWwxyltFum7uQC0NGzLL9869gn8NqIZ7G1Cn5DLU99R9m7s
8HsWpmdKUnwv61ENapI54GhtKycNnHxTxkf0MeoJQuMUnNAISOM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n+fc0fpoK7nTCka046zVZbQbLzjknLso3XXzbk59wY/Yhl0gTr/XdliUwOoK
gPrzudodyPT6v52/6wOaEjm/TeAPjNQCVZJoB5Hit1Uikm5/EXT+pm3fAvAv
nPl+FZKY70skg3JXqtnTnJI6H9WvY8sGdefi8TbHmIUqs8BTcYk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 17440)
`pragma protect data_block
fnAK/nv1EmVihrt+cJftmMxX9I5ZGPFeC8ZIBXfrvuWyKJxLqlRttGBC+OzR
lfQPIqHShMxqLXQbWFiBHydg/invG3dI2kqbwsSKmp52iPdTTx+cJByW0MPy
5682ucfZq4D/L1ciJen1zqyTc5WroSHyS+3816wKd+lh8IzUbX6QQtr/+DjJ
0Q0z89AtVX5mGx3pnIc9wa3kIngun8l5Z9tULoU7Np4xF6r96tx1I4vA/vM8
gka/OXFnUtcMuSWxkGn9C4XEMTlmde/bt4YeNDx9RVOQeSqpOSopiNmCqUPC
EDJDQQwSbD4jWH/4SLhH4s89rEENgBsQxlNfDJ2yuY0pq86+rHFQ+VIEj4dr
2+udi0W6MR15vEWc5tEMuE9W1+vjDGcrnW80GWO49gqHQe4jOHCU9TL5gbU5
0+qcmO2vpeDDbL0Prn/5pHqm094TI5QCORlTaMvNEs7a85c9/2gSmc2O4iH4
hiZrnDTLRfqDDMnv7tng/LL8AJcvhi+1rM3Ro1eA3Y0uKvkunAS2XdpXQJvV
YPXGwQV6V4UArMEQdy/V9zJZfub9NiJWEzeJliq59yNWI6+pVEVwVzfktQxw
U6SekDDld3NJ0Dby8A2vgAA86OnPAvY4R6P9QIHN/XtifarEYewjoOyrcFuf
h04OUo7wptzkg/lCCYQNmiUSQyxqes7OJatfwd6Q/E0Yl8eaGgkBENeF/Sfg
ZZpMBSF246vGWoCa97J5CfDu9jdSMf/+6NiuO7kiT6abrO8MUnYK3HU6Jyep
yM2wTKOPvIHHm+4GGFtiXO+7lQdbzcgXGRU34gCuc/1BvbtQjnLDpFvHSlRV
l0SMWXIWcSJf6uzxMCVedQ0Lc+svq1FQ8IjyUcu8VWtdqgOLMt6S9UIgoqTu
IgRatWyQut5IdrWXBDSwnbPMtx9qBDX8ZgA/QLeU6FwbByML+uDmzzTEesmu
Q2AcbHBJMdw+15LdNpNeFV5CtANI8ySP91afAD0cDbU2pl1HJ26eBLem1GUg
1MUw66iAY+z7QQqknECKksfPtc1YKo0WqWsM5mZRCf9oIKVrNaXd4L+UbJfD
z7Ez+Vw1TWftIUkIuVF8STT5GgLY10UOmKS6BaFI0DqLBTcQmGrI+douUlik
plZNnZPIZjmW4qa6PQK1vUdhIdzOsABgMkIonLQBSO6/XtKaZrWUcgDeGSPC
NJ8D+RX/mUBQgCsbjtacmE9+ST0DkI4V6k8RGa9Q+FICdeARilEPA9DgY0wc
Apn0tIfOj2dIHVcffAdqyniDQYE6q0NN/72AfcBYfMSGfy5J1qFfQtiQlO/S
MMU3mUcMxXR8Zk7gmJDRRyz+xI7cKXTOZeJuGmvshKWWCclo/PtdFaw/ZijO
UlYdPq05txUFb0yyTclTw+6nCn8/VWXu8w9pwF0PELAwjDqQHZ67Ax2uzb40
4Qs7A2R5ObnMvpptboUpxURZO6IzwIHxWfDu9VTtwRufZZxSF4iLMfwAXzyS
hkLeqIXTtu7S0pabjq3W3rKBCXqC9jf273+iDHtCqVjxHdK0gdQsqAoTI/rZ
mfaJluGM7xDya14T82lLS6bK/sBsphMclGzVoWLHiqRt2kuo0zu8WtdK+i8J
z3YOq/bwWiWX4RyAbCegt2b7ULBtvPafDZygbZBVGVTVzej9ZObRgP0cCm9r
Zf9e+4zOVpUJCX9zI0RAYr0Sexh8W8/ntDlOLS4c4jN2BPvNtVA3ZUdhg62R
V49UxuX2mWKkXye7FN7iMhlhYv7sCKulnUXsRk5Toa3M4ZuzgUYtooWgc9u+
SuO8zj1jgJKDuj9M686ppeZFuopR2TCL+93MvLqwOq5REbAuGBAyftUTWa/y
Urj02zyWhRwu716z7Zh7s+nX/gyButTUWaDiI4dEnTnHaFEFzB8s515FIH7t
AGYpQXWUROd557syK0800NxShZvENEdY+LH/HMi3AhXqjD9IsVys6WqyhHFN
MZGzPVLqFCZj3U5v56wmuoGxxhLT8IyV/2leAi59bHrMpLNQJv5Jenx68U0d
rACQqhUkoRkEjm8iguVToLizNjZwEp5IuLm4gpCcnyRJnf89+7gyl8+hutRy
6JaFTKw+sH87f1Dgou1jNwg1wOyBSaWeJY7+W2fWWaZfizuaVzw74VjdNCH4
XWdPKwZKm5MDo/J1Bsb5a4kBSIyLZG6fOWk+hz49Ru0CYIB3uDsz1cEdylrd
iG3qu/DHXtdXPSuihHOZx24Q0zQudmuub6ycfAbxdPf4m102IUWzx91gRnEv
2OZbqAddwwIK4h6/U8yASbPLTIsK24/2kKKPzGpaH76VeHyyao9H9WA0S0Gd
odxSKYH71i002Ot46VTWxGGLzoNdyQLefWn77OiT4dEe2zp8ibxPhZofLv1X
8L+vRTLza4wVnmDeS/WwyjOgu1Vpnmqa1/jliGWRBG0nJG3iO5tJ13Dc8gD2
DTdAwxbs11w9XJAGb3PXf7zTUZQVdxoVV9W4yvwF4/Tqrg2RnftM+xm8zxAL
E4aI/MiaKLSVEzbKF8Hf0Occkb0S9bfcx9gS9FAi/+w8GPJDu9F4L2JoM9xn
4GdeRXJ7E2H//d9oacsKJnHaDvXg8VibAC54fNB176K+yHT7kSSmBTNw3LLD
JB4jkzE4+JvKx2Z5eYt3r/M9jSzzr3mJ2S3ekoJA/kTDgkW+uDcgxK1M6mvr
Tixj+ikhfkz2Z0mq/oGKH+iOU37wuRhZiQGu/+sPBx1oqzPFa3P3Fx1inO4U
Md0VSBqVvSgzbh/K/w9zafP88xynON9heFvVwb9dIBcnY1Dg9cOwwo05KPdA
SA2KciID3IqsDOkgWn6ePEIvA3mDLprGJu/HdpiSTG9CukgTwaIXnaANIQnm
kcNA/egxS+wnae6r0bjyii2s2b3PA7bTxubwwvxI1csf+sVwBcA7n+8J2iQW
PI02Z8V1KOwdhGsijGrVoDikgOOZe9agtM9URNtQcINGVfKzfKMQewxw+9Dz
D2QVdfqhtkb6tN9ztmGYvYBwqXeLtvO6MKsNMyiApG44nSJ42oeQzbtDPxV/
nCM5tQ42cZIfgm4rnyjqkvHZ8J2DbZOZQXHz4NTuelam8bxRA30VgWBX9QVo
g/fv3WaxoxyKXRCFCnGYNrocRd9juzg2hBRonHHLAjxsrb6cQIyfgl/bnJbB
wAUS+mxwSsoZSZ0+u9nOmrckYZbc3rKfzN5Uchkkvxsck92Pgr4wv/mUT/MW
pWpg1Y68cg8xjLACCICLwIojRjk1qJS0o1Ptw/gVxdA/RP4YmgYgP9G9U0Tm
Iae7/BUSRNVW9N13v65QnaY9aCFzw0oHRD3kU2eWTYUH5DWjav688K79Poj8
8gxk4hUVoBn7eiSqGasFJFKk0+gm0B0RAznTObN6YAJAOpS34cgr0NMxTFPF
xTJbewWMjstaNcKTzPOIDlrcxpG4VJnDxgOed3KyuVUnnAMt6W2SemEdrdL6
7V/90zSDJYYyyeUiVTfdkn9Hgs3UUFmtgGUkwXeVBMav8bwChqJZpHhU+cWC
X2qip5orUuWp9cp5tVLEbt2y7an+3rGqvebXcWLjK7+iW7H5QSbPcdrT8vNq
b3NQmt2Q2YWRGBJciWNllRQoPccird5dAUoKL2DKzkG5SNctaAcZLX48qw9H
rkhD46sgKewLiYQatCTyNvTsibCtqxotnauwv77UW+pOvS4Kx2BVBXpxS0D7
Af0Vr6hFrHp617FysU92NA3ftvyu4ulqNWgTBbYsfBHmjPkeKeE9a4FwTj2c
dRBErRk/dKYRml/j2e/USppzsDv6GRLkh4LH13W8aSNlZtKc1I1kXwK9hh/s
TaLKNYgQYXGEcOJYiOIA4IuBFKVyrHVv3MjYVHD7i+h5QOE0aQl/I/GIbJIo
/El5x8mfdwp01LWXWidBQId8kN6WI5r05j2GiLy/7S5FWLjp7gJUJ/g6Nxjq
RsW6yNUg9J+J4t2mRAQsHrZUImyjFFskksIC5fEKvzzcBYSFc3Nv5dEFA0md
TrWl/MPBCC3nLtC47+qOUnqETDbYTRxqLbHILE67NPi9qK+721I1/Cxdvx/G
RcaEqopgE4xKwc3vWARYZhtnS114epcdPIDvzQHvI0R58scR6wEoLeryC+ut
a38z9wHg4kdKhFSnH55dHrqksheh6EUAxyze1ZMxM9KSWVVRr7/u21l3XlF5
oiqO1jqDKizNnV+Xb3rGgi8wNC39GBy/0cMzeAJZgFLDWUCWdKi2jJaZJhpG
+7qzWBzJpWXhXCMp5OMyjj1YGgkGDMWhqe4g2FXIKOPl6LGL9ot0MfvPjR0U
u24LUkLD4NkAhc0j9tJeZU98LC/xAEOhBY7uFXjI+yruSbe90s0EC2I2z4C1
LpFBM390LtNIC0lnPpvmAjg9sxj5TxHZ96CMN7N9ae+PU6RciutoFBZkXbUQ
hBfmxx75PEwgr9QVj0oJ+vBnT4ULwmoORLZpN0R0cN9iGfiIOgzVfnRl87EG
Vu8mgffFI+WDFlqU2I0Fu5vcNEdUZllkD0PMGb+f4HRAmt16cpxZcxFuwm2L
ETQ6XDuPyFZ0u+lVJLYNvmtF5bajnzrVmZQDuQoy9fLBhfgnbVydRn4qkPFe
3BaOOE2Tzd0gnR0zhwklmK+Rn9dmOrAHbsjdsQqZdiSXuO9eMm8n3krSiBuX
P4/u0gUu0BLWVy77r2VjmVmsDMwMGbOA0cKN/hBdgyz6ZFFe6NZo7/XBBKpP
05r1xh+KPjQDjsSlXb2ljlJGT2IuG5hLDdZuMmoV29P6EmNJPwxicUMSvsaA
f4+HQMyAUDRVZ1iPxqDZl14TjHMHsI5sjXtEUA1yZqZA0oAqeWKlaycsDhq0
zMblcRppocf5vlrjA20YxyE4k+4ImeOT1PVuy/V7tO5FwFvbGPQw1B8d6ggM
F6Fd6LFCFcL8Fp109Ie48Zz7sxurdS53PeWZhgooiYapxiSmWSaUamgvESxx
oyFjE9J3KAL/677Ips6sJX+3u49ZBo3SoqBiVvfHgIkRtAVemMeI1vIMU7GY
EzbZ5WW5vgAjwZPDocK69CZK0SU/puqScCwlucLoQrWeDI50SeODG/Cknybx
hKCH3jgVHTJGEgZ3MVd9h/OfNo3dsX5c16AxRCRmgnQaFLLfh/sw0pXYziEk
i2s+fHgAcAy2jgNah1TNbw7OnaYvG1qTRrtEGKPUHithrW/IV+LoGF9UmFfF
YXFDSBTPjJ0BNtAeAQhtStNs7CCk/6ui2VEFrwwlhUgtU+cqV64cOGdcQ2cz
73P+mu/wK7KgdXEGeEM/yXNwfv26xAa5CCVmcWfPcHmhczbhhFfZ6mVYkzZ6
Svm3FW/ChR3rOc5IuTmTXImFAC8gB6uBicsE7NLxRgjMdubASYTo4foaWyOK
pghxKb7iIj+VUOwQ9uq+nZkR7n+hGOrcU9lfe9IzBkoJfOW2FzjFcdfqLZxp
lb4VV9lqtOUi+b7TPyW1gotKZCZ1LAnBn98oqq+1IBL+PwafkMCqh/HsyH/v
LNloQ2njZ5yxo/1zyBVK1pSTYFXkByq2+tK291+U/BV5HOQIWZAx3bhADWHg
2FlY4M73F2es1cVxOaGTIg5ysClTieNKtTMB4VU8E6gJcqgJ7OaqH023FaOd
jjO3vo/QlBt1PWlpqcuTZbmRMB60Ib0/YrNcQvbahEz7HGcAKzyEQGZuRM6a
mCqJOQRyjw/w9ZUNoLcUEv8EYysR0vm9nvcq3FMW/++l6K+cqFXL86ZMijCf
Vjy1kNPXbiQr3OYTAyKdlom0oyP6KusKx3HhFV+XPzAYf6YrLmyFBZ3oUb39
k1QHBYMzVuH+vn11sXqFc2qS6JEt2KZC3J33F6+B0fJl94J5tEYBive8qvaV
qT8dF1VDf8jUiAAnK1J3N+MkFYjLoyXxCiWsPXB6UQhp0TlqbcC08iSqElEf
2p7HhJ1S+3oPGLzDXrFlV/byLr3TscBhA2eGayI+u1uWp6fMijWYPGQzUpPI
zEEYo7RtuZNkrm/bFs7wwsrPuv9FHd3ugQMag6YZH3LfRxOZCLmVF/AZ5m8h
A3GPKBt/MfqzQY6UC/Uh+USAehStaKQthMmOHngxPaLJdLhAyb6EQSADTfnT
UBBqZ9O1kt3uQdQKewDN4UVAjs/E1siSANpWbDZh4toui9P+FO6b4/cucGhp
uWSncpnrV1Kk2XxXXsxBXTQV9S0DJLDsr28o+lD8EqZE1kmiaIGKvRKMHNaS
LfyA4v8i+mmW3qg5N35lbsFGMVZUCnvRJ7+n4z8/eQaYuewTUE8pbnzj06VG
O/U1M38nzU5p6PnhVU/JaNiWCcv0pjkiWQg6KsTLpiTs4Gw21+ooJq+IZ8Mc
ZB4cF50Ew0j2JbPJEnGeWYOeO5vH5eui/6EMU07x+Xd2qJ41D/gtFxgFNeFP
W9qaLKpNlcX+c9QlaPAJjx/74/Vw7K5MsiooZCVURVlVRwU0zSIXEsaV42E/
5yi+SMseEou3PhZ6j0UPW6xgnR/6HH1nDfRlQBUUFFpBNw+qZm5lgh/Yh+4B
ufa+7CbIT8WSkbgqW0mm8idysASyTGseJHd0BCHbW0uDsY1d6V4bG+DaL7Jn
mfmAODQb3Y4CDiiVCD8k64DrQM1TNhNJLcZqwtQHgkDBwltJwQ7+CQwPAN4s
IT4ifwpaFxCjGNBZmAGOqr4KlnF9Rm4As5HJG/uClva6IJ7NmnNfz1aebYMG
FCJiEW0ehgri018xECZXvVkSuQrLlwLmNW35n01HBpvSV0LA8iQnvfYJ6vy9
iUd8PvsjPYtERIlaotzxX0EkhMkxBiqgbZtVtpv5/2G1+LMt0HNR6jloRJJ3
jWG0iVwaOqonGpYj8hfRWu5khpYFz3PdQhE77H0vVqnN3g5F5TqCpcrLUk0t
mWf8fANh8enevMvw7odVCUoDLxAYW62yRZ15hfqLtWAv5IUBQwnN4qKHcu0l
qrF2UAOBtfMFh9kjD6trqtNefFgB+5zteqY4psH/kgWqA3OeswsTKVXCiBK0
zM1yzsY8Au0gqhmvrpWIyZqE7JTnkVSdZbkc1hBlzlCkIWfiVaQTq+8KGxEt
s6MRu7r3P7pOIsS80STdUHe8L7kBKEwgjJShyX1ul5HCRgjgAAskwyEUheG6
10rhCCPIugzVvYdcRh2QG/Tk7BKXQrMvhtTudZpANoaQoI0XYh67TV5tq1rn
PSws9Sx7vUVy4bqj6LQTxyDD2qynQYG6WdQXTEUfHSm/haxfHYNazMg2zlyw
e8ZX3IJGvTzB/3l2JBOCfyfEO/9XpUtTOS6SQEgkYrrTwHCp+epIB04TTXGb
9i8QsFDXhntUwCXiFug9f+rs9WYxk4WTJ3vxoEQAti/jdkBAl4hu3Ol5wfCD
oQ0s/JdOqG2eQg82jNuZhB7t/QSRvR+faizo1ZhDtsl3BUj3vpLBPczkVbzT
B9g4KCe/8Xy6uhtye9h/JSx9tTPDG503hKUZDFOcwAginJAiUw15I/hIft9Y
GNafZL3frsHvOwId8JzSFtQnYCSzViqz9UhfZTsu9s5EQdf3VUXUhqZbXWmv
zJbe1eRSqsm4UlF6vwFSHsRB2SgEH/7ZDhVhlarkSF38JzYGPDYGIN66y8Ma
WemJoStj9NiM0YFVipx1MhtRDrP/Vir5ClAvt3eDb3rB0+YQGfKwTSLpAycg
fliQ/iOCuze34SorI6x8fJcNttYdYH/8RpvAfkFhX1hyTgoEiipoezy0FyY9
JigJwdwPZ4RPDzs+OL+3IMNuAWhDoteEJBLBSY8HNIz1EBxox+VUPUQEQdiJ
M0b8F1q+0zA8MCHnZKzvShbB7ZNJWajNxJXmH2J3v9qUCucpE3PkQg9czqf6
tzJPZW0sP3JVn7cjTNYNabEmcK0P7CoMD2xh9Me86GgNhYB/jlhFftgmhFsW
I4WffyYAbhHz3q88RQ3KlaCNdG89wuOLmT7blISlJuTzgjoDOaxS4pmLrac9
KbtfY51zU2J0buOJr+FHcQkBy/18/t1IZ/sRPVzCiUCoMOyizaX0M/i/zthm
SPjonL6/phEGhZ8iAinYEHbHsf0cHWWasKMya2GnZ3e/Hyksy4GHkgxcZ6sd
apTy2lqsPi/2OvPKodpsSgsC8fixPVhI6LXYcWVehu+TUOsQoe94goeS4mYA
pG95LIuvyR9UfBtP5RVTM0Bd0CuN0a0d6I2jl+iYG6B+DBmrJpABjKsTEtv5
lcGRuvM2nduk0UHd/pXPTc+GJVGe43i3IxCo/RmqsnEB00ixz0uXNW/uzUR7
qrpRHSMeXyB9RpEAca4j68CC4ZyfBAlD9jcUX6chr+/EOT1GSFy59bM8HupP
5fmuNbVvpGvko26KG9kLgY+AJc60dsFA+bdJ+LsOvRCREVywbMHVSW2S5iHg
ilkFttg4K3Y4pj/RYfuB//PawpF1R1HgBtJ2EX2eLWYjs7to4jciQ/4CtT5h
xvyJn1764H3sIectW9ubkw/kPaHrrVngyt0CaeOrPZE5IW3KDR9bD2xuHPxp
Ip5Q9iz/rlmVetYzclM2kUdmFApfHjtxETQgbJtXjtfqhuM62GQ98jcsJehv
GY/RnnjOxs/rRW/jbxgoSd/pXu5xLWC2AoDtp1BRt5gEyXJqOlCfUcYBHVaj
ha4hLiAH5vjxG1cZUUwRAcbMV6xzVaVMzOj13iPPl76jyXiiT82wxswGoISK
xwo9or2Tim4gIcZfzm4yhDcx8kqTqTLWp6HUdVuo/m3+i0GvTxWFbyvvOEZ9
pgN8ryPv2c3+yml8I5kjzj+hAeYg0BaZ/W74nEHtUN5Qf/mcP1r6iovsy+KL
vbndWL48iu1GqWhPmMzoAu5ib9zFz3SHfFFxiGtQD/8i80294Eh9YhQ77yHV
MFybG+64WQ+KhGSPSzrH0SzgiepJAmIMm2D5qoND9tqjn1N1D9ik+m0IGU2I
HKeg6eL1gl8HgmK6ipa/7hJnrBcg7dZumJNgvf4eT47uyK0XpgOAhnPqmGbp
VsKarDN8zsnjWvpUrtmagRcwETy+7FxDTkQbVr7M+rvs76sDgCsfCfOcyJen
oMUsabXtfZrxAoAZECBRJI6sZziiw8S/c83fxiVGxnU71/Ywy9i35Yzaoqrn
dxpKfLldW4MokVPFlh7VLaHtXQ2KOKgRsQXjbXtvz6xF/2RI5+H2gk3mSqxu
qK8EozemUezNx9xanY8V8pb5a6LmM9+8a6PyfGg5g59dlq/DNJ51s9YbdOMf
CGKjMTZ3qWCvy8h5iHER7DtIgs/J6Ng5Ly/sbGCheiUXkrQ9UK/Kb8wTfIAr
jpGyNwmSmuDa1z8gCwBvY1nNV37xtAHf38i7zzG5oiITskMClj6q9OzW86B/
pm51mjPhub2oxh/GZ5r1t01iW3wjtw8ufyYHkekuDItKQo722XMPG1wfb3x3
dbW825IXkkY8uJZWL8wUart3CVoy5Y4JcydlVq2UwGF//QMeiuQV4/96q3f0
te5ugktCWWYzC8pBPTKEN2lCoAmpb1s2+cf4cQJO5+wUL8TGtJr8B5vsl4kg
UkNS1+RoHKZyVKT+pa+qqRseswrrknaqkzCVmaVO3z68ZlxEw1wydGm8UoqH
fVVZJ0sYsUt1xGNcKu+6/hMRLQ34zrdTO4uR6e7A2UBh7soxpCM43Rq4iJy/
s63W8Da9v6Ng38f6UzHbYNStFrzhgTPC42zjmzgfRSrRNWatWUXin929dI2/
4AkjI+quX7N0aWT09MPFcW/u0Bs3ZrCBlzRqrHfDaa3CkDNHmdLoYLJILJGW
Q7ru4+MdaTeq16Fmrt/juZwur9eCUIZDUztlA08ySYmRo6nBV6L0eU/fOdee
DoffY3FLdoIBV39SnFqrD6rwLdkHXkOFzS13zRlC9hREdUpI7o6yd34FWhBZ
ucmjazoPfEkocFAUM6ckNBsXxq0cwoIPqTQ90SlpugZQkNftuiyOcry97RVE
PHfN05kLYqPXNUCndPnOVlp8E+WedrSBx05f4ftg387SsvVT89l9AuADC1Sb
Ee6ErYVxkQRq0QbMdJTENtBGkaRyiGx8oVeP+vVfqcv3yb+v0fN0c+Uuhes2
3NNHp0yhnhMPCDE6w7LY38c7wCOAs+J+UcTbuFOurenCEJE2vgSiN0r7Smn7
c/f3ZrB/CkNlN248mfXt6D4GB7QWipaaxzP0c/qHS5fmUEiCtMjsOogHqqrV
ebHgFo14D6mJr1Mp7infS6tVNaUxEybGG8QRHes3a7H7iUb/Bx5D3MQURnye
Q8IdWVLCdx4eszWulvvq/H0QBVVj2HwstlBvnzYbI8Dg0gEIKQFYXrLRn7r1
t7dBv9WwDqk2y1IK7/MgCPYoc5jaQkIWNvXFRgC3JvnmrgK+FNKawX9MLtPu
BVxIpjWIwwzH9P0r4dj2G9/Jg0RPMm+zX3lVO7I0yJNP9ToqIbyKfKcBhjqr
tssIB8By5uQwViz6dpPJKw6Te8S9TOrAsDY3gS1uMujc9oCp5aKragyl7nkg
u9RrV8lAd4grGaGlWuSCk2anH1KY2hiSa5AEBXOEFX82kh08WG6OkW+p+Kbm
vZgFAJAre/WejJW0Oi3vGwnu7/Coh4/6Yf+Y18Z5jAUsmVvS7P1h7Q0ng728
hPxWubwNPUtFZxVjobNRddZosAKGmqtYb3MNMXJWpC9POmSbigznQYsN5Ygp
/TPsBwSAp6q+GR1jOUY64ByW7IscF/nDY0QIo62YZCI6vgk87dE5SgpQVhtn
4dfjFGVwQpIfCEANa1BEcDoCmAkTTfgzHmpI+u5+oSmGvG9kP/yWeLqM88Lk
o3do5Fp2m+VURwBKAKR8kbONDWy0iZOVjBievq8z8+G6mftyuE8xMc8fN+IC
bVnET/HydQ0U/cTs5kHkVj8yMiXyS8Prvnz9rD7S1Xzgxe+4ptAxttmcY9Dj
1VQDmztGnkoRbCuB9/kUfL8b/qgeELDip/OCwj+WH0FAhZybq1I4m2m3kvye
OrGx6H3WyZ7rfvxU6QXZs9OYSQFMi1kM32R6Ug8AHJ99iloaijr0pPeCzVOW
d3LY11wbr3z5Xz9CK2TMcYoNuM5VAW0Nhry1QnrLtQZswmGvvKhbOizoC/P6
ISn21aA198Iq8f+aB3JxROy83b5TO6rZ0wQlPTY0jCHk6yo7fVNuuLJlSP2P
FAkZHzFkh3VyqXyVzvQ5lb00Rerp4/V+/zTe4l6E4wGGC/pOdIz+TMYs5VAa
aojUqvWcX1OTica/H/1rL/fNy9VZt5zpSL1J/htV9j6UousZNU/hso/x2ePk
xdt9rrOYF6csFxFsWXXa7jyCJn4JusiimtFYAyhffWYikSBPuHI6vCp1ItRN
sZPy7Er5oP1cUZmnoN7pBxoLO9liZEjH/yzrJnDfA+TiQz63CrLZ9ExyvP6X
mJ1/U6m+WwAxUELTyve0T53KHrTMvSZgi4/gW+Saj65VdsUuAjhJtJ6s1DYK
vxjHDZcUPBM5mmVBGAnSgitqmDyvHJBSzEmfIf66muwlaMEQtkB7iIlojPeR
P6AUO4tBgYBvA2J2lsvKuzLqYcMRQ7lOZ+v9ROdBVXyDPpjTcvSDQ4M9KysK
UYBegSGM0Ol246yDqB3SJskRXGsf2bE3n6DAvRt8T6yoyfdcBCLYJ6Umi6yZ
ajvWTd3/+PiToAt7y2XcC0HPzZ/XTq7RT1WDodHpx8N3gQq0yTdWUr4hlDwX
TuDj7h5uLOyVbPOZm9sdJimnBgNIOUumMPLl9JuN5fGgOha1zIZVPGtlBW9x
hAVLV4BFs+tRXNUrlNYYaUA8cE6xk6UTUVHBfz2ihAHGX7eO10fsTfATJWGw
kKEDezAz/QFuoyK35FkJkTA4O3sRY/Kxuqngap10fY+oaPWNWcYxBVUo90q/
wnmmlF8SUab1/o8SzReugvL4tPNsH8uhPIhJFsFqaQEyPFJBNhr3E0yeOjKx
j0VIk3ZrIvWwxBHz99nNooZaEiQhkp1E6VMsCVs8Ld1Gx1TqFvo42k2yDMBH
jK37gz8WLvOQyYWGnv+tVfeaVsKc0TVEtRsi7Mg1xOuBW9gH8flYcWpBsX5Y
C3vNkcWFrPT9tp8FL4VGJXfpNEthvR3WNZJV4GQgFIHxaXvSccH9BMrPAVY5
7qr/8+TFQyJZAycKEH1IK9rLSX7MfNdS+16S1T8lqvRfJ37oVDMzlCAJLFQX
gdOE0TjANl+mAT/N8o3fqi9c4XRRXrraZqWDi5vS0+WI2kEuUF/uzJz7mlDf
rTgtRz9FHh1HZuzzLj7nbmdPeaN38q1yBFCEc3tgdqvao4mIvDcdy6jFLzyv
8IjpStjdhxzW/XomI9+CMQJDOlmCqzR3AedG67BK+n9nAzZSPIFDyCF9D6o1
qeUfX5k31aeXLSW22FmUfyRzG7+yG5h2s/wW5B2Kyzjm9H4TrN+BeIndfPSE
Sho9QSWi/+SK+kh2S0qV0G4jZs4R4g1pKdX2HuOJoD/vCP9VzTIssmppBOht
cNYsOv3v1hx6aHdVOGog68XIcSGWrCqhRj9ltgESDL/hVMLqE/hDVxMiCpc9
KW+JaHl2y1IywZbodQ/ceLak6gXOhdmIeQm7w5MMq1WhEYMHpqwigZ14akLQ
wIs6fO4YSWT07felJaJe6qs9XeBJ0NB3zEC5LZstNoSwja9rDiGgYkVIvQsh
o3c02SeeRmC9xmDaplXprO5RQ3PZ5z0trUKYkrKCwuK+6aWaFVJbCmb3GT+y
x+GrZb1Bg10b0Ltz3RJk9yztVfgBGAyxTgtkCco7QjtKCDSX7RJfWDaH3DgC
0qcqntnK0lggrgFtOGSZZF5kOW7q71hm5IOiSCIYf9a89dpInrg8aesRFTQS
7M/JV7wO81jRLQq0Gev6gvEZIb3HuXbTq4CH1hoBMzBYSVXdS6nVXVYAWVOb
jbXtou8noCqpyIY3Na6iFBcDU9bcAKxDRvSw69rgEw19kGtdg8ypUoNK+XFm
421AykDA1qnQai+IlX1TdT+Dtcvo6S9a1f39Bw+VbSDrZ2fvO605sLvsPNjk
QMl2mX7hm+XvYzKWzPBOMureU0XBaoH3GokeyfOyIc5WRFY/Hn0TaONrbNis
4tCVz91aIgcRMVmoR0kXIN9B+TQnoLutvYOuhwCcXnNOh2nmke5ZzlMTHoC6
ZM5DWdy05dp8FFcdEkn8PZ8MZ141P6MzFmreBHXIAT1WUf841/rh9iAZTYQo
kuxQ3Rhe0QUsuR/gkjwitt3zZFwm6jjiLom4Ek2XjD5viPAML05ZtjE2RzAt
KVQZaHWfFE3HuCSWqiiWWURntazKXVa0ngE0P22JAlebClkBNH6GSarxjYs5
g8hfPjoFMsv62iNlcDlLeo5Xl7SalDmx28rr21tEAexXPGNjqTcw97KdIcgb
5OpWCxiO4ISuUXQTprkf7QhMiptBrsY7wabKf1fiyyfv25P19ZZt7WXtMQF9
2+ryuVjU10Psz9ChfZTzeV4a0335Znd+ysWxl4kh93VjgRouzR3FzShVcLwv
iPD1WbpIvzj2zr6guS7dh2Othhj9byAqSsAkbOEPZyYnIUgSzSvtCrsQ+Gxc
YODWALUJV8a7bcRJApxRyEkX1otemnoFoW8ZHeUZ5JyzHp/vhK1VWb5M5zJY
BWjqljNvgVnKHJegxkHSbR4M1MRx0ZKFcfYXT1CMi1pESGaA5pKOs1DtZSTj
aTf+VDLQK/nn66AZsIfGQTugxFtIK9iRBEhJl4MdaXR/aFkk+8fj/0vGA6BB
CWvpLO+dqO1ETCEBV9qhFUgYUFjm4RZasAOq5/cp4FMRg92JjpDO97g9u+AY
K5O6XKY1V8zc1FQlKW7ZIE+pEjcEgMwIX3q4AnAqSz+tI/D4xs1YWKSYlGGj
i6ebmytRbjqMGtECuNdfsMrkcBeYFum6+JBPIlBle/iF6HEnN/L0V0m4SfKi
4/QJAJxrijSUB4PGEIpy/3ZayjvtupJEDtlwdm5pBFM/hTFrIJ8zkwzNC4Ih
1vCbQr/xDlBWbPk6qJa9toOJd5Ww+FEzJPgcVE+3khG8E+HB1k0sm5iLNu0M
gEVagMr3uOQSJWRolmtp8HWFQGFr4cHPNlADCQTC+fGz0oOqfMTVXD2V34q3
dWwN5m/Ys3oOZzQ9rx4gFg3z/WNsWsM84RdpyJlV6ciwpBn48vWesztJ5Z/5
hnTCKm43c7S0L/z3bJBZk8PhUtpMdvtUyi1ivf4Rq1dkDuU+wUi8O443AoG4
JsLJqchJsGCJPPXphkn7cOhqtuFCW4CZFnsAuLPtVZjFyZ8aNTK91OBy1jpP
KA1nUEeyvDfNmbEuwKfh1HC7A44kDJmutCSDvegD0vOupV7ZTJXYM+upQJiB
cmQuiDyoNWTz9Xbw3kGYnew/wtpvWFSHgKMKb+py5gRfaFqqmIYeOxykROP9
QiY7yKwCskJJxL8W04ah8D0QTrgGCXYpaMoeeW6W/kQYKWVZzX7U8ruhdu31
XyNkus+DMoBSfFOHjolb8iLovcX+omaxO+hSi6MEfcR7an8vnZcszlNRk+5O
YmyP84YcJVvb0NkktPNy8azLQT36+DlSPk6tePdcKIGKqCtEXXtWQc0Zrwqn
d58vrQ1CEUFlZ08UFRXQzzWrnKX6jvzoleCSD8zNww95Yvbtrd5kY0iiDhin
F4N5IWYRmI+FE4Ogya0+A8k4etzfjjQWOSh/b/PP3EtoRsV0e0nK/uKr2OVS
SEzoTAA2lfkgpQai+38E+JG4qcHZghsCnDtnKQ38aH7b++1zq/RlZ6CC/agI
qgvyj8stZVtB/3ciadcPxvIJEwwddFA8eIrj5BSqG2gr/F61NZlj/E8wvzuB
Ti0gyd1dEI9sIIS4vv++58syPDwWP96uQSJi7yC404c+3W/FGCskwj3Qdsy8
SOlFoPS+nUfTs3pzBALmd0ZVrGGxMmkPCuXCLPR3SOymRd/1SkCG8ANls4qh
8r+OMmuDTzgUa1q65MkYAEwIgukPuYKSureZfQuSitLfxdBtd+MhInDgYP4z
rxZWbMjitMKqLn8c87AyCAhG/93B0xnTNsb/5coCbuZXyeRjKLc/le4kjV30
ss7hT1sVBIv+xrGRCX8l2o/kaXmq7eOWTkW6emQmxzavjjpgbb4pu88QJxLu
aHa24MWKqjBUoIN8ll9IWM+uwq9n7GFA+ywGuwZzg/Sv2qzTPWitn9B9qftj
q5hKVrplkfJy2rfOd9tW1SnC0ToSuVSvB0YtacTFOJGENWWvUJhKK71vZcyI
uhjuaZdH38WAEPUOKouCsoGsyDGSWJ6ObYPovzQEua1uStOuxi6cwt0dIGPy
IKLHnCqTxZOaY0L2fy/vn2vJBae2WbqAgBMKi37OU0tMFYNe9r2qkxNhdBvV
cTosy44kkSGoeJ4JW4GKy2EZ9qmNqHpnocx+MpFEXFDHJq8R+yizTZYYmsEp
DM4ZluhlPloehhlO0zQjXsnEj8v+Sx6u72cm25e56ntKGpq4sjhvu7Ez3RdK
2A/3LOCmxpWLAOYt+5Yj7qOVXiy56u0UcKc5pGHbTknBohz+RFtkYiE6L7oV
cABhJSf8hVop0KzhO2hQAgd+2QKT+VHZP94UjEPgzgZPG3tWx1y+f7teE76U
VZ8kzFAxrLhAB1vOgo84O7n4JwmM3aBPknxZ5gwlFCRJUoOqfAMR/Rs4vHlr
7iFOPuDGDQqIU/fl4vFpubzdD+BkKDdqLHB+8JKwg5aIOZMujd0vJRDD1Rd0
k0x+mHk35gq8aDIU2rxez6m7NYshjzdBFxusTPEhJxAEts719P7jRD3N6kAN
IbN2is/N7Uiq4PiRLpp5Dnbnqqj7i9HrGSPHCcPVmAEDFKLXmxQ5Pq+9KvMx
Whe9jxxkSk+dVZNAzb0u0J0fdwMqn9ANFOydlp7L/TZkP9cZIVZ6pKTxh6IL
4Ed7cgfdabP4v0in+gq1A85YqvY+Z+KKASH4zuIc89x9CZBRXSYHdX59FQcv
mSrKcdkylpGw8OZSbL3KkHlDkCCq+zWoRbHrbqd6gBZUiVUvAcFHY355SKBL
2vZZy6g8E5/mpX1knComzA5qw/YAXYp5caQcFp9Ddnh5ulo89QzdLx3GHXUx
8H4542OusIsugXYQ4fvX83mzKopgVD773+dFzuBNRiEF83EDzq9/GJlr7uTm
Pa0xuvsrgpfHnuIAtc+Sj3htINegNvbmU4xt21BeYVt4PC1TTXyQ5sMuLkOA
gBGWru6W072NTJ72Iq+B2qmBvbi7gawoxsBKedzl49eVTi6J4CK0YuyxeZfC
Wwwf1cuucVaT8aqVFUrP1O5Bm1lp7+tt9mN2ikopB3Y+S/1Cpztw+hKPIO3v
AVWpwAiJikA+74p54SLLoZEcfrbVRLILdCfem3TBAmV6i5PAUwaPKgAp+s9N
s48Sfu/etU76lU9XQi9pKZz4/gUT13jPM/5mfWfVHhI2DWu0iHtuHuBEBbsC
XTrG2hmdP7MNclwTqwoOL/206VDbmYoFajrIaxZUB08erihnxglNTrNoPr0b
zXC48+Q+1akDj42seknL2BaDFxV0CkzgOULtz+IdHwC/4U9t8oV7ZplANRs3
mXBHl9EYJPcGCYS4D3VzM8QCQokwxxnZL7jvzoJdj7gj2uWENcOzoXeOZiTn
bMYAVQamUr9NEQ0h6weuS9VXQwnsrdKnyXYUKFq+7UiCr4/f/1W7Y2wu7N4u
mw3x1oOM44+U2QeiXTfsnJAAzuVUcIDgyhVzetCJqY2ogYoDefSwWHtDOQbh
UR/3aSFV0+npGj56iQTG6hDkOjVRXnTm1nt452ZPsgBZVJ/dI2cY5tMldYOE
aNLGgQUtfCW3t9V+swEBlqxQhMo6sdKVLuOyWnQVn9YQ04YI/7+OFAHpP324
AjaNx1FVMb+fGkaKmzKguu7WXPQHmjpPKxkwQunLZV3+WdvT5mCFxqdx9Sha
zB2fki4o23g+IWsRbTJcQPaeJ+nlPhGGvUJTq+sONUXid3N/6sPL+cOERbHd
EGm7ZqcJomEs0/LwjbUqGj4QZ0YfBXXN3l6yovzJmJlJX/tzUCL7IQWrzxj2
UrSHSjY3rZvKRq8LTPSjKGK+ixSf8IemwfFOZd3IaaqPNHKPgwcV0czGiPEL
VEuBQxjOkvn8cN5MIN2nVzyIs2frYb7mBz0tc2qgh3E8ioMDGIl5uDpJ/oJv
vYceIjXpvsW1XYWrVpMh/VhQjVKzDOwe0euWC0ZpU+wFQ4X00RIyWa+Xb1nN
W1936VP2iFgc3uK3Pgl8g+n97Sc5BhyizBD5X507V5XNKMx2Y46fv97BXJkO
FIH33ZQJzWJEFpFIJNEa1VpigfXned9pKrNoayLcHxgacpIb0Z0RVueiIgZQ
9sdnvBub7nGeoHIS7+HgZhENEsZHP+zpCvP+iF6o99uB00omHDUyrW6Tg1Bo
08oRCqWxaHbwvx0HBfBSOZ4rfDzgu0H11wFjJUPZuSE9LyK4nwUCBOOvFpok
4+EBbMsPkuDsibwbbh39ZmRHJwbnEWmhti7Nmb+MionJ/1BnbjpAReYZjnD5
WEedOPnDa6U23fJLwww4x5RBHCLvEF4i9mZJjSOlwm50OmzToaA2FLhVQUje
waocS4eHdP/+vDAE9aXGt+MuWOIU+X3moudxfWMv2wpX48jIOeaoxQAQZ9Hs
skcPJISXP65ggxfCVtZJr61vBf61qk+bDY/P6wqcE4V2o7iNTS45XbTRrjpm
rtUQBs/c0nKmpFmKTEWM9ibBXJclmo4teeJ/7sBwPztHdanbEE0FlmP42mdt
2sblYnFT3BMGBPoP9wN6nmWQCOAVmzHnB0W0VQnO2PpPg8yyciAW2V1Ulz1r
hPc+bNae1q+VljRIiIeqnmob2wj9Q54i7P0wBl5Gyeh993mIYcepX3qzlKEk
qoZYTsB7lD/y1tfclhOEROZQeNMiNo6y2XCEFZPjAk4NaA0my7HT7MEx+MiX
V/dd2ueMUH3QILeKY2x57bshKU4oYqwR62jSfmMwVA/SrPcgtrzLy1aUnzZv
VpJhdKxHwCQdGCzMtWkxnG+V5AdY/fhStVF+UQb2T38VK655Mm+bhQfQsivg
sVfyLpODEV7w2/gG99aKEvGpChJ1UtI7rhkEQGzvgcuEd92IxHMxeqrDLUDa
t4x+NhFAQmJCeX8bIeDFt8fhqphyHWu3pAtc5NljjD+itGzeakgPiff6cyRk
Wox7rxPWPSALjydGYks90IF6I0CxuqUBAgkXvX6SJCPcgA5Sqe8nZdHJYzyY
TIxCBH6FWtsgh557+INzKTBev/nl3vaqDBHbxqrEzNMiCefnYUa2BhL4cn4N
vDOApAnBL1S5t/PiOq6G8lQJQvZwkyIRr1wqUndT+eNta+RuBJwDqp/G7yJM
ie0G40zDK4neh1ebOUzkTpNXJFTAGHwy4cFJnbG0xggR9PXG5UUtAvcC+/XF
0Kr8pp+PTnHqzV3K0OOyuBXEbbckztmmXAA0EJZyBP/uIsASm4SmA3JDzWMo
tuRm1XizVlYP+SJTrS3D04FzPmpRrcpxXuY05S2XcX+5nxKfWqFkBGH7XNea
JZSKJ3fhHaX0RLFTbYlk1EZh/lgsFmCGGMqNieHwW7BMv+ySILJi5GC5589L
6yxgX9Rr0X1EzpSj6ii0iWb67rFnGN91fNKt8ia4YQZCFP/2QoRiVfsv7qC9
lyTUy2j7z3Jj3x/u0azDgtObQHLzdxJdwyYqMp0IMhhydKcFKQ8rLQFg447v
e9s+IsLhI53I5Kx45N+aLrgqtg/Fxdg8pQwyqkW+eHd++575LrAVEMcp938j
aFQFZg9bG0tO2fdeKUJwuLaHiCVoRXy/IFt7iunL/pfK368FVc8Fx6b3NDKf
IdySH6ywxncqbB+oQaITxjUkq88/Qtzz99YMgTWjunGLGU9YstNqHXFEZw03
6Pn/7Nd3RZr3oGaggFXTZPk5cJE3+kHEqsk2EX+ywciRhkAj++KIXUz9FBeX
8v9SGXTatHhV4vY/9NXfe0DEralcJ3YKHxS2digqcRu6ZXIsWH+eu5FQ7A0w
bDWCfu+WVk2GnIeQJE4fx2tu4kBWRVLIrn81BWR3gfyY6RFWxoTaHR6n9vLb
JRqxG8lz/lKjSrskTqy9dbD+Jg22Si7PrH5yEfYj65wt/c0M9s16Ih7T1ues
IvxuoLrKdzsAXqXhkpfq8P0YHJ6Iof8KD+EmDqkcpvRSSt7Cq95vuXHuVoY/
7zCQD2GHiKcQhA7/05etCF14V4J7YQ8FO6iRa8BbX4r3TKqtOkCG70EmZ56R
nbIoa65eXYG4zj2BZSkA3aI2AL/1dDcK6QU+6BBU95Rkx/idVkqfecxHsQiV
Tfdai6JYmMqctLo+cKS6s5CSjWP2TeHTZRqsYQPvANaoYNNWAuLeEu1eRZfq
XfkXl5yrqMaPJsyPFIRJcWKc9PQ3Ki4y0ZYjIGJNHxDtc8C3SARcQtVzavEY
OuiYDyzF1nrQaxfKTAX4JQ3mS9IjVt9Dkuzh99R2LenG3J3EqOgfjCNtuVHK
9r/MIfMUxz2AtM7jrgrxJwQAdUqL0n9PovIUrC6HOzXkv5fi4CbNjmT1Zb49
JaDzmdhGKBvhe/wR0vbjyQKUqpbrUTdyoWSzONYFiog9Qh9AwZ8juQzsnXEW
sp2xuOYaDZrvo9mScGW5AkRAT3q25PiJ/1l9Bd208c72jdUZc8+KOooQzH/1
SYgK6pUgfRK0CYPklg/cMckJdHy9UyIP5WBl9zC3p+gyY28/KrQJwliYtpmn
UaU69T+i97gBCDuP0gWj+mhN5Vt9CSD9TFdW1IZFRqS3MMgrGrmn9ruJu7lO
U8TulYNWkiQ8Pdq39YR1+2M9Ur+IhWjW4usgYiX41mOusEKxZERZjWfcxZvz
p2pJQDmLymA4SchQneZqNsD5E4VMidLyMHSSbQ7jRww0VQzp8b36fTTjxGlp
kOvvi0RYYCotMLTy5R4ib7vcl8TM92e5I5nNiBmnS0kgHgXzw1J93e05pJLh
t13zYOjz+OmicMVEuJnm8AYJTsDNanU4BT6+T6w0X9PFyk2qZCehiB2WRWXS
hytzggfs664KNHEI5kcBKR5N5evwQfSzrIzO3BSsWc99XS98Vq10F5igSfW8
aUJn+GMwG1OFnWQ8fzrLCuzWiXG9RXWXKxi6OtjY1Y/lc+52fmxZgnPo/3G+
lJEFwqFq4JjdH1yilDf02XCVmyK4yKWWbVE1l/XqySaJGxGmnz22kzHbkSOp
3sGX4/cBc1nu0Va975NW2ezbAHS8N7ECtO9CLKl5d8QY9DA1Cf0W7uEXstDV
bYuwX5tWdrIUPITT27//KkjkUUbjLD3Aji77uAXpu/4jyxQkdqkxGBSEdRtM
0N9GiLDDBTfIkv4Fa4T7H1w5hE53bUqwTIZSyzk19vxWfSTePCzgYLVNLqMk
/nYzsvfTi/NOhDpL5kAN2jueASaTE8Lms9n25nA01oH3EIQd+NG8ER0f78Ye
HjHVmOFx4562T14v/vbu8PQeHhmA8sfymhbGiWJ4JoFwZ0Q8hvLSXIpis1UP
R67htzD+talt64JVOEqDqxG16KVjqwJ5zgAdSQU2ex4miFF+qqLWxDp1HE8H
kSa6YyRiuY0EzCPdUCwRoCMPFRR2pQ32aIEF3kA3VZg5iSsRsAewZLaGW4CD
78jHGkpBjhzG88v8ZMPyQM2lrlI8QGZAXt5HtCx4vzxCLIiF7ZnOpf58GNtW
qfbZOGpBeoJpSHXVQ84xQ0BkKKSLE0xjV6pDT/jmJu7IRKzTRNNJOip3zLcr
KvLG4FzkaXLxtTJfIFKXs8c6yyfgn5K/royPjLNX1k/UvsR1jjKs18mwELAP
a/NUhN24CD7ctp6oGiLqf9ItZ8nCBsgsiY65O63tcA1Z5PxfGuAQahJubnwo
y2ocQN7/Y7jZ822rouRrjMyHLj3N+XVJMQ2RU2Ct1yEAxI5Nq9Itwg+D3KpK
mWSKqwMbBZ0UL3laPFVcvjTIYlYjB4o1eBxrxMHfkN6CWd6A0ml+wfXmMCMq
3ot+1CkDjY74gpcCgG/lStE8QPZAvzC4kTGO2GvxdQF9VirJo4Hq7sJMOcNV
0uIj4I5s0GaFpCfo7ZCwK+87bNspraM3/Xavq9ypLwTC7dWrwRaGElWMTVxw
qYyTV8FFYJpa7X7HbDNAmBPhT0A+7DP4t5d5R9+Y4HmlsBGYFZ/OFmiXDkqT
ka+XTO5AlY6M7rjinONfCg8SKTB0PDc/rZSZxhW7aSMXCGOf/iTkJ1F9AJ6Z
u0pSKRxlbX3DFFbt05XgYr1hAISX5lHtNmhkduK4EwmZCyhgSU4tF4rh6KJx
RTmWBqLS33ot7+jcmeAZuU0F6UqH8EhWgorbC0S9fMY3s4zlV3gx4ieBYj7K
wPvTJ6Vchynb6LaBCUI4Im/27B4XkljjJdX8T7lAK1TEo8un9Exo1gIRxGCM
bMSVWdqwVjXU9FFMgGWxdxZY4Q0rJDoT5QhUXPm7O88q8PZ7rk2rVUXRHg3j
OiShUhrOXyrLjOqInxE4bY+PBhdg6h114wyV7wi7e8SID7qsnv9I4ayzwnGN
fqSUR3MNNhcAyZK1ORTG07MdNjfUQnGmrfO3ImB/JAFy4n9h8RpHf90gaisv
bHjrqC2MqY5hsKum29PdH7YFfqSEZBsj2uDmkh58XtRzMIkUSTIi6C6V62Hp
qNKKqNB62uHBKvurubtu/HgLuBXikQvpPaOyNsCF7HY3cvgd5WLkoQBeFdrW
86VUoeEYIFgPzforFSeTPRs8iU55fsqPCrzlrAQY8/dSvUdzpbA0tS2iJwpS
sSswqX4cVA/5wOgxWLfKs0g5Evc8lMgsTkBvoPS2tHTeyw7wHio5UrWz6d8L
L0IJokVxRvPikfwMGyeqA8DFqjffOLk+jgiotCEBEs4s1mwRAXQiUAZb7f1V
RwaGtq5bEamscbkovRd6c10ATCdxtfVVW36GgjNvkWz1Uhg0y71qwEfIgV3o
maCv3cg7eInVihenxO9OqETN3REFsSCaSFCVBh/iDnNoNlU7yzYLikLbkNt1
x2GGmVA7cx1L7+o1mX/YECPH3vUFfWYqQXDcOnkcs4CqG8nVj/gz/Fg2gJnv
6xVdmgoSMmclTVIR5RGrL0PuhIcZCmcLeDbhajaVZEEY8EOTiV0CKocZ6MSk
71alKgwbMc03vJUKedEoWsCuOdIFoGcwf9i1mgc4uTYPCfKkpsDOCivwJgT/
zvlXGoEYTOgCb4WWQai5Vi1QJ7lNMkooX8moydrf34wwa6ZWKeQnIEg56SHW
V2V0OIE43aue7r5vSBzk9UJIGIYbWpxhzmBAJPalTsNw6cMT4aBXWzozDVqT
XLElJKJozeUBqAlZxgdw71EHXVWlB4cT/39JQWwVKou3jXo3yM6hCQtH23Tf
5Xk/N5FVtFD9YiirCK+RBOBGrCQV66pmdGUIJ13SRkgw1L5HGEBxQ67Ec2W3
M9tYbLT8AIiz51iHrK8qkymyp1moT4Uiy70Ko5p2AtXmAd6zSzKZzmFqdA38
sERr1f8cc8o7zLBTx1wS2uq1DT2KrzgOheNnY8G784t7oNIk0qCg97wPN4Cm
sez324nDSZso0P7Acv5/MLtKbAYTljPbbkLJf3it4qEHlOm0/b0qKhUaTLQb
QczM0bG6DKxQTzdzfpk6qa/bQrdgdCaVVEvpsyEJjv/CC7NUBm2Nd6LJRxOF
1pvbVsTNeTB4SjYHtlK07ITeRqpriHIASqB2f7QLGs72AixBOcPlVEKFUK3p
KlM2JCJkV+mm7cGOOvziTph3BBh7o5kUiz3jq4RuRshD45ns23hieVV52z62
PfwF1Cn1ePHw1BdrIFUm3Ixkv2D7z+OTpordLtIAEKAanLyao8dxaElj87Cc
5+GXmWCbr4Z7qc1g2DzvyPcfiVWMp4rbY0mW00W2xi33Gv91fLteQb6tJftJ
aPHGUqimMfeyV2Te5aEDESxrpKOMKU+6ql/+7x7iTmJKGg7v44aHFzyr2I0p
32J1JWnHcFBdAqNWxu0b8Qpl6r79lc4bdOVMfWmCJe+UeWdmOxFjSnKFVpzQ
yFjqfSor5jIHaVDvtZLBSHAHE2T+yM7AL7+Q9bfGkJ5JdOd+unXMIIKhxYc8
RJnr7+XUahJrVG7vOn6wop5o4XDFWb5DvDLp71iV1FEGo7nqu6HkpwA+jeYs
HvH86Avj7gHHmOTu5h7ZgHrWXEed8vg0jkGf+nW9NDw1GjploX8UnspEMVqv
7Oa3CE7nTkebMSD7PncIobR2HBIwDqPvVA==

`pragma protect end_protected
