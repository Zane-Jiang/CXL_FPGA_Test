// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aT3G5idBjoxgF2U4qYjpHlQBfbgU5AV8jX+CSRLSodCQOUSOPrTl/wd86wff
gMpwheQmbHmUTZJFOF5gA1Pxcuzejj76u6IgcuvtSua81LhjF0gRM+pUpVI5
/IcMV1sbLku/G8q9TdCOsDn10GDO0RJAiffBf28PE28csRCaTyWDcJ090N/5
AA0h/MVNmEiZwiw+vxFBEljDLyGBFI4snLMHuHKHmJXXdSiIrZlDa2RbXgKL
wlnOqGz5FmG0Tlg11u7akUd63FxpUW2Z9yc6vMdxw54mxvq/kkv0UFD1DfUd
K+xZmhPwsMhrjLk0CnrHzMb0Jha2d79DECXgjMA10w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gVNUTOKaZsPwp1BtU/hmGuv/9BkHjcuwW9BAcPxuaLUh6RRCZ9dopf1mhydI
YC9u76uYYkXdhuWF4TQhvbs7O3EPksuj5PFJ7Jevi9XnZXIrysj+Iiz37u1R
wh1RP4eyvo60oXaFPv4QfdCfneHC0CHaZEpkHRm500Yl0lvj29hCP26Oo63f
kC1KUYSNN3dg87/pOWZy9juykKf8ok1qz7NQBixdhGtdB8H5wDpeLJwaAG1e
YPMurkvD7XIIzS/+BLelVS0/qmD2Mqj8DadeN0SZ1QVfh0fxOgzpjY9RzHmV
SkjF0bVk4c0HIgqGuJN+kCLijpGW5Sgi+pux1+JLKw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BVxNyO2OzHC3a7KJu1qI8J5hS/zrhb3SnaxNwEkHbbHKnxxydQmWsDhnYtxS
oaqZQIi3kMBzxwD4hZM2+b9QnpWtKSwrFt/oki/B+NrcOiKMr2P9vWjRqm5x
+qb2h94n56c+OnQyLARKz/YIZYJYNQF2F7qt7UgZ4DmCX/fFGx6SRJ4qM1EX
CeQeh2DL3wv4WvG6SHb8mrDc72xPKtax/6K/Db1PleQ6lVbJg/dSBkhaMGQO
yZD0c4B/KJ914iEDmY/MdDZfbXBEgbRbJu1zHzN5isoufdbZneumHyXAWk0N
+tBJs2e5dPhEE9e7drOcdmzZIQrZsZ3CKotP+VTDTw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WPc7/oje2NNf8XFkozvrlbWGs/rdxR6zKJ40I5pna9DXWvtIU1Kbu6XbOit3
IlLOzYhdqKFe2suAYt5xLNG6mJKPsubHz4w4YJJbwElFkM0WjGwUE8OGNrM2
AIZzHXfBVr7E9zrqXPVdXhBTcFb/DFqkiRdOmU3hlrPHOSN3gR0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Fvh8cMAMNajCRqsEOgUyk4z0UvcX5aVlx+czCUtB3NBHt5TjLt141LQwHVjX
3msCMlDzrkKDnO/jAkHL5d5hAfkjYuTyeuc/oV/uhT44FwlCirA+jo346wzo
I7sj/PoZs9G8topZDYDtPXQrlolW4zOieCF72ky3EoHv49eYMs2TDZvAFMEI
OoEhnzz6lSY0sH6vMn7rxJreGVxErxMxpBPaniPNpcnliyzEGtuQD+12GG33
8NEpLRe9qWnGkcbToNp6Utu3tfJwMrXdO241fFbzKvktWz7eky6Gxv/tgEyy
sc+bazkO/1Y6ajM60iZtifBa7qkdzgGAk3xnRtkb80DF5DFnqgw5RZC3SHOY
u53Tx3Xvr6IL8NJEGrS0O/TyghrR4EswzxV66uoDRV7LEoq69pNXENqFbAoU
bnIrYAwrgy4pi8w81zAExu5m9FZasEkJCTfF5sO9ack7lvb5ab/kXmFBpndh
sEUScaPcP5jqynXhh5vrN3krzDQumkct


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gsvJs1dQzkXLyeNK0ieHtJTRdwmTQYGW2Q8SUogVPmkVB/EmapgNu6eQ7nM5
jaAuktiRfgHlYN4vxqVoJXhxYA6QumqxXjEc8kubKQhVO2Yiq10dpscllaHs
3AHGqgt3GkBMXvh89Dyc3r0S9KUKQkweyM3pSmGRWA6TpjMvQNs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tJewd/bJnRcXmPsdTXbBhimVm6uw5y+eBJAfyLFdqFuudpPydMNq17XreqA+
ir3Tn+Vsem6Jcx6PcCI+jn6LCx3VV8BUb8m24IUXXBsrhKdwIKMtSXXwgCbY
wQKsWG6dqA1xcDAl3f7iscB/gf7mORoL7CCYt6TQLg3GHOFu/ME=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2784)
`pragma protect data_block
pRl+/FWZeWnktYrLuo+q2nkEoS6sAtZk+o+1kEpMZBfGvzq6phI/TP0gRKEy
1Xo4wcCNQJr2Zw03LMj1R86FGBfsjMwKnpLQ3Yw2hp77rYFE0J6ici7DzCbZ
lKH9QTa+MhYBTg8qIA22hdCwR3qS+ES9bDhdyl0rlTI1aQwOdmFrC9HWBiX4
BiAW3QKM5QYqci+KIK4sR5rOCEwf16QDjGKLnIfWKIl9wN1LYd/Mbt6OdY+n
uWaHz6xsXqOfe7/HfTv8OJ3wm483NcmCGzXw2roSSw7HJ3ogSutBRB2zHocu
f9+/or7sUTQZxtbsavlMxFrWJ6G/zxB+E2dgBq+ERwxmMc5SWN2rKvya6flq
6B4iuIqBlh0Jp6AnxsZ8wiI1cVG6F8JQVnLNPP6k5+O82lESyk2A2OATozFg
HsVUtuvG3an7wZPIRPYf6irCmsOtxzzBXAUCrsgRo4wGCv8OW4tbt0q2i7vR
FCxoIyq/ZQD8M80hP7KEGVFmYSGGZtPOvwUtBkxyuY8SNA5MGvNfRZ205h0O
WyBbhfx6pTdRy6uIDaiQkKWHQQSVakd4/H/waIHTPdKXqfqS9XI7lQJFWxly
26Jzr7CRCE2qLq7hgWufnN6WPH/N/c16W7OPZnaRJ5YZu5bWYujUKbRl3OKf
RRk37vL+CKq/Oi/bYZp9GO5vLhGxhWDTx5nHXZAM1JgbunjIkEpDQH48F/Uo
sGztJmDtgZIjeU2MiW0Y3SDETUpeFQvXu3aheQI8VRf2ozOJDicvlAwsnIJI
rHl3WcMwiamFDukAo2YfFoRp5PTatMTrQm6mdK4PH8mVF7VtoIHKYXZ84lAC
QTapYA0WPvBrZCrZYnI6Hn/HMCWL+1F8aqVm9klfg7v8IWEqyaCWhaAbia1V
CpoygkXDbPctL99aOvnGwZNCQ1TPFMmCZj0CnREAnE3DiU/6wqbrksb/Imf7
DDKFiO2eLNQr22sqMfdC75zwzEUMsH0fjev1zuF2L7PYqMh8g0dQrLC9h8s3
fAP994oa/cKyinoRVJWjmwahI9ib/mckGLZM3KaGdIfF1RJZiLW/OE1MWjId
yc8c6uPHmNWlsXUI6nlNXhw7BxT2xGkdu+n6Wt/JPziRp7d+/3NWwGKW5R6Y
QfSxm41xQ/BTfuOp/b9I9m9GADvpbaWjCV8jErXfK7UxnShIZp2o/9K8Hqy8
I0KYBtxD7BL8ntL0jXuusi2+3ZIMn0oYmiEoqsLemYplpDNrWbK7UlYp+py8
myRuamYiBZVKZph40Lb3HyqTwtAfd4TOkazWrLZBUiju3PshbH6GAwUHpq/o
Bpagz0MGXUymIHeXY6aZ4gq9SPYdR/aHqPnhi8trGZb7bpi4yFPI3/dUqzHX
VTivEFi6UuyH8NI63SRjJrh8ZQJMRlIZo/6yQFSvuFFMTfrBc4CwPs/1BPrw
YTeY0/7ur1a/Fgzly8lkj2JkHVPJMvU7FXpqkDwMG10WmSQAvpjWzMWwzboX
lHibEIHMvhYeI+9vnXnjVFoscpbACzo6JOd7n7eJf+CPNLG/q+tO8QeYlC1j
8jtizq9oFUXFThYTI1fcMsX4lFTAq+SbBFtZ3IGh0DWBieSyjIu+rx4r4cDV
frjMDqSFjmM49OSZ49XEnIEJnuxXXkI3+prGLWtKfeMtWdV7Kpkk8/peTNec
TUhdjGYYuP3A4dQcnFhojmRcyaLA5KbCZmUxtN2kY5vHO32nQrr14iG96w9b
AvapqaSOiQmNUYgU1zUR/TLsDzs4iy9IXEQRPrlN97/WkzxOtWXDsRX9oSaF
PrnkHNMlb2rPBJH51hyDE2a5M13jFYJSuNuPoKbdG5KF/B118DwBpCRe5Set
P5eYBiecmvDmzQ41r4J1ziPyXn/LuGQfMs4ouqaHT47J8PYCUo9Qw37fV6MO
RXImQpIWNIU4tYh4w/eiMai8eOtmwBRN6T7ABMb1vbEkbGf+w67SeeF7q4LD
ACUAHx/id1+u2Pu5xRoRs5JHPiAEXsMCFrL9U6NGUGnkIbYzDZj2CWulESac
H+vFLk2NBpttJ9OP/BoVSlasdRjzFVm4wWoem408V9avs6bzNFRDSKbHbneb
VAZRuukqUM2DjU+57r1L65QdEYir7BTPPHDVWyknj+BIAbeoZzLgTy7dzlIR
Lw01IoYA2wpCsjPXD48moy71sCyCtxRmkO113Az9BM9H1pMClr7M94b/1Vte
I7aj7Xopm3z9qOzlX85byK8LRSOZIcXAovmT5RNxmG1jalvRvuPtqbgJa5Hc
PGhQMJmgS0DhhUJ0X8685QdgfbVJAOezGklJM/JKNj7g3tr0PAHrQpCjqVwo
bmjHqeHR1gI6DrE3sCRIqO/PiaIvzBMinGKd3tDO5hd+gJv6nz2oVIHo4U51
R3bTuabdkqstvTSAN5htKWNbt8r9AL92VVwwd37On/tbM1n7+8o6prlZxKjF
KwpFOk8VY3WRR8lDvosbC75mHt6H3JakKdX3GGIWPbGVbBKVuVncK6mSOZ7Q
4oaLXxk2nqPvhHwU/9R8S3BGv/dhpSSE9bFE9WDamEdVS8pyBCchPtOUMzhf
Oph+1eGSpS9MkcYSM4q2otVs4VZZp2HDJ335LP6pm4Bv0UnGp3TrN28Klwn4
9OdC+6smDLOjsQ2ui22gDXfk8PcfzUxD2YE6nnLxNTzS9tZXJxORp5/9kcLM
gbD36zKW5Ha3awhJAAFJXiC24Xlu/fVH0dblQEAurpz+qRr7O8VVC20owwAV
fxUoc5eQ/txKS8q3H9sYNty4TU3ndRr8Oq1DFUXyf2+rpGQLJiE8NXK8gjrN
bFtzlCKXsYqGLe0JsmStGWLTKNEP+vR27GjardYDhJf7+f6IP+cOgu+oD2j/
TrGkloBYIONAkY0/Jj0+cuKRMfOSzstLAAy/yvnEopXk9PchELrzMf/WmuIv
hJDhn19yBr6N+ibsgWvEWU70+1MmPa39oSKOMwU5CpBs8/HFxrpWgSbN2LwF
rG3JOjV5BL3qxz+af1CLTbeFP0jzQFOlaoWR0BC2BT6njTMzcW3S1wUMMMzM
CTzbk4R/m7QBj24AEZvs1cpR1kfLM7/zRuuTaHGnEyRvflkVvKZOh3KuDeC6
+45OITFVWKmMWHYPjBNJbzNs83bnLdBJDYGuIyV7mTpByKVwOfcv3njSPRfS
qjgRBRlqsVJdHxTbQdPqjbzo79LfPnW/uXgxn3invUM/jVaRUNtb6SMYzH2z
IiMWBw3o5gFSUthQ83lGmyiyeUo63yvfUNJ4BBZgAysEk3xh8BryY+i5c4VX
nptVmzRh2ar5cNVE7i91l0GQhzyo1616VptHqH+sx7iyFbIPdQZgoBj1ufdV
sxQdb9NzoVmsvzBMVQBagrWijM486CSuW3W7koNwbg3toeNepPvm5aYZRsxL
zUjELJSepbGYwI8b0xOON78uhyCdnL99ZH1GGTgNYOY8eXXN/4hBBvRNVzZH
i7sU5qvyxwaqkF78hrxHhWgBmsHJNhXc05ZG8w/MG4Qeax8OGpKmBV7pGOET
VChRlINbERUuwnOZ0uTCNbFt5zUe1uPh+vljnhrrfmUTAfhxNV4tN2VKak59
FlYAkxMAsIHlQFIjdLvZRZ1MIrCa9gBD/BO45ZccF2X2dyhsfqiMKeskoxQC
khvNtNN8AZcCg3xo2VJhkkteuTvwt9BpilrHicX7SQepExibODqv

`pragma protect end_protected
