`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
OQBJPRHAzvkhAlMv0AaPc48jFBL6h2hcdhg27jdzAtWgsYAdd761LUaxom+I7D8L
+QdUptETEVFDIc75BWQC83v7TjUImYGv3SYqaOyS66x79daShAmIOS7VFnOa0Y8e
uDEHSw8lIYOXYmJ0KvqTB/oGtf0x43RXUdGWxQfVoG8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 50288), data_block
zs2c1i4GFwD1oVNcr9RWvmDVO/tTdhtX90vzPH/I5U08X9bd+h0pCob6VNi7oqfC
wqcC7xDaPBudcWcr5D6aKqbHcF07r+bZKBTWkyNGkwpsAjGa0wLqsL5AtL3JT5Bc
7Xh8hA/DKHM4vuIlgrIbVLoupaurTIlACxoaW6a3sTSZX1Fjw0XzdwNnYzkhKK4Q
tPkrFLdyo318TB3fzmgB34Wn70+VZqTF+i/M6yoAnWQwLfK8fdXdPobv3aNhoXf7
WFTR5JPrL9jWULl9NogyMyg2MEzqyKEf9l+PlJ0GyHFNrjPQ6c43hQRUenQeTxws
2sqZ1X4ZuiL7qxwmFBEgxDMXrX6OEcyWNRO3IgRsP7s1D/m6G3OBjiCWLqBGER3f
R5aZHav18K5DnFYwkiKAvAnFtmey6qz0tONUJXleKWnBvma7aeHwYbi40eMdK3pC
rFDSI+4N8jm30GC9QdD3N4E1z+82mRntUhilLCjTrSavNsU1tmgxW7PSD9Wu4CaV
v+zKCStmRGEWWz0fB12TsWiNgsRt5+XMcRJI1MAfbFuJE+FJae8jvfRgMDToQfiK
TEiOG7EN4Oqltt+tgqRBvf0/jbZ/AumwsS7boq/V58pkYIuRXYqDpZeh72OttPgk
GKrk4H+DImHQwtEvqKECCj3VkCojOmlWuLfbPlxXzQw6LKmitq9dx7pqmqlrat3D
rK0VlPnh4YT/EDlJQIRac2FTrdGreT3Z6l2hfU0aZ71AuwPNYn3jCF+AsS0xH3/D
HndFQ0F/bGMoI6IszRkz88Ww6eH8OSYJVI5bDyx3QnaEMG1hcJKGtEbG+2O8iZYN
OambUx9sclNeOr+/OrzWJAf4l1NrPbYU5Z1o3GCASXB2xsSW/H05yxwtAdMrryh1
cj4ptLVpuF2ivYFbblkJkl3GgRg6/9gdD1/fyii/waJH6WWBEmFEwhYeJJFHctch
wBCmRw7WTRreAaSA0ramXIpOy1n4JHDG12XZ1E7S3Vx+obLcJwpr74xuV0x1e05m
20/b57YBZl8gCrSk/YTJuvBckiAI8/3rplKPhnKaBCdqcfpmuIxOPvG7IhYYMK16
1KRXOn8b0LVnMfYkCcO/r/Rg4nLHG162DLIBPX4hg3EgTMjR5CF6aoUkPgUoXcwg
DZQg7IFizeHTC9lBKf8h1bDbGaAf9q3TtNKtYjI4460uleOeOE6OTbK79Jd2+cgW
y3umlVS/u8R2yCFQcwUW7KVlItVaeOd4Oi2weMpkA/TJ57jXzmB0QFrPD+l9E87L
89sOv4K5jlQTTvTm2ZcrRUMJtis51yfNXo9Zx+F0fs1WXiXWilzJHSgPUZkBiIQW
VaZmUcMBtTx1HumcGGU6yTTADnFlmWUQcrjaU46ca7T0bVmMHPcIQ9OGlAUDLAy8
JTM3BYqcXGTH+SBp24nmKGNDipvkqSVf4NZqoKzUkk1X2MryERJIw21gZtz9bLsD
ZUxVMWugui9Ap1c6uFhM/29G5oxwkHTbzWSv7VHtvNtmFZEoQLfE9PLAcVIdh3Fw
T35NZt3F2KuR0mLkcg6lgyJqsviFGhkohA0LJ58B+UXt1btsKEz/KyK3ziB96cGm
4xXbEllH+xaZh8Dv7+ECjdC/BhDx7yPtGC5v/H8F5mAQun/8A7pcKoaj4xjG8XzK
8WBHJDIAQ2Ss4QWmqFl1H4BmBXxisOdupB83rq1i+GdxvRbEaB/U2e0LuVz50t+/
mxfFuNfGO+VJE+3eBNSU8NFg4UVwUs8jxm6kk3Ap77EvansWlgyivnlSCOT7SgWl
o3zwA884F9UDUG0AIiTdm09Lf7FLFdUa/xKjX6ouayKdpavow2r2AV4J3jHhCHeI
nKS2J85lZgEnc1wBknOKEeF8HemS6oUKXpu+zdh3QQBOrSmcl1vSmzfjHzgrTjoB
XmQHc+gI06seX8Ia6lzuiBqTzIc2yjaAVRKEsivSdv1r5kYkqBK3ms/OqNgjIoSx
CHq0VzTuxcgZGY32ZdR9+L3V59Yvs7iVo8e7DHKMmHiSAps07l2d+TXW20nOcoVj
6kqJWDzw79wv9Z6XYjLNzPg3buYTBpX5iWyrfskjAQDRrHVYfc2ooiiOK87mgLyA
Lg6tOGuwzC1sjRUSMgUQxafIykofKOUTuOLEuXDjMxPMDso5AAG5MsF4MI2ofPRI
54+POFbpp21muYarWmGbwZO2YHI56UKGXAMFbiMe2Uw+VrdPto5rMvgRfP9KhpNe
fb6gOWm/IEC327/u6re/H2WbyY2UtU6nV2EFdlMIYE1kyOin787uaG/V43gF0Mpt
TgaqY1eD+Y/xAb51FALsQLvEOdMmQcp8XXludPUqPB1dZs/nkmlRrU7ffHo1KHM4
KpM9Cg1AIC+YYVsnf8twjqJo7d45C4fvfQ77bDXpADB5igZjJJjcTdH8uXLl3Jw/
0X3nf0KMryVLfMUIXGn5bcQ8sKx7bwQCOYXqH/kd56rpNEULNDqNeuNUr6wQwEzW
hX/x3lImDOXVeUFJIt5t7intzwxAGHRiUi+HjldMa3NfcV66Gy6DOu8cjfsGHpl5
82UGYCUZXOO+cpZxbsAChHxXnN4QmC8pLm4T7tvycjdtym/uXw459BLXZjo3wfzm
OB23ZwBh9irMK1ccvf6rEuwD2ePzQRrR+aSV5EAHEccQfVGynO98V3wd6/hflEk6
C7yRgCSngchLNQN51S9caR6q91PdVSk0kjwi7ZMcaOwCt1wyZrDfXns3DknPn3Qr
VQSZbX663vXI8SHkU38YmdcaO9ZM4AqyT//8zjH5FbgUvxh1lfCusolU5RfkFagC
09vszwC6rxUrZsAXiYAn7X3sXDwUbCcOTOOW0A4+MboQlY2N40U37UmLWrdeXvYW
0/Jkmr75dj2hj/FMPDp34qmg07sOBJwtZcWXj4kfMX9eLM51FIjZE+eV4D1ej9ph
C9W7YMVW6zo3eXeznbw5NzYBSdRfs11D1WSHqMxy8ems7//SNRFW6liJaA3LuNpD
+sGlvcy+whMKmvgw1VyZt/QL2p00g16/C+cTdJdSLncmGmhxaDnw2boh9RVwS4Qq
rDvYboAhrlo2C9D9+v9bdWWJLrRFrHNA5T6OXqZSgrf9Y41sSM3L/8rHdfECcQlS
xj6NZE+HxxcKTcA41EeqJd+xkeA6O2QP6mizO+L+zVF43HIynx++YxN1rTJxiQZP
5Q9ctZukmH1o1NvWKXyi3QfxRpfyjKuAjaNwiblQuiw//KF+Q0V37T7VAuU+dDRa
iBtCdkS0mnXSh6W1RCHXwUZATj9kF5h/OmqRsZ7TYgauVn3Upd4VLQo2YV++1pbs
nQvL+VF2QX/m7XcsbQlv7LzJ3fTNeyRzL2vSDJrD5/Y9TlKpxlD+YG3rV4ioLKs+
brevoKNekm8Deuk8QWM34eiCSqaWaKiGeXSjmn5tJNwZOKHRlTTdgF5uScFggPLf
e8YekyDvs7OsTLISM6CCMmDAcAlQ9ozvtwRUHlLca5959q4rKybd8Huz5uVA5LUR
/s2tayqNoJ7UJK64VqTKM9z35LqZ6BB8bFtr4dZuoaPiSeJdSAzi0Xp6xzFbCrgw
dq8LxD0qoAGNy+q0jAIQGZEawHhemskpsuv/hWffqNlCEAcpy0wAFUCc7VcdWRou
k2SUTRS7y9KY1OgueZsdghktO4d8+8TPPj9wIFtDC1TlWu+RE6fHePBK5FGrLs9K
WjlBrZkeVyRGpxytKGu9j+kvC3Btdxc8ndy1GrIlHMxpuka3W0WaCjmJORRxQvLN
OtmK6gsDLkcYTKomk6ZRRnqwzK9t71eoHZBsKCc3apiL9BgsshkcF+6yFxxYqqJ4
MAfoXfAF3igCQUxaxOyqL8tBMwTY6DM4npQUOoBY4H+lvelL6a+X0MpPoohzxvKX
TtH7/gziFup9wolq0dBPYCYm5mv9Hjil9DKZSe3c3Zs8Yw51JFdtAwakEguHfiXJ
AKWkEo+DioWL5yOa4pga7f+wlO+uAka6lHlLi6P7/6n5gyPwdoFtCSAJycIMWPvU
QjHMQCN9vmGOUy9h+YX3Ou4AWro2GmiN3FbTCQkw1VMZIPzcoy8iv3GieCjE04hQ
CMX4X8gfXhYGf54402+D4evOrYuMNcFjGBSxOIgNshxFg9yGdpwpKYmhlejg+mIj
I9lMZrcmYKOhI6usCeP/ciXU++eIo6mnibphqwgHYf/HcdVg6YuA9iAxyN5EjPIR
GqcPSD9O3RG/qxaJlyCd3btld1V4wyD2kDU7KPMHXfmlUhJVCyn4W5inkF+1mxT2
wO+58iQqgGvbcMgUnDc0Lb0KHe55x0drqjIcBetcfppfEVuaLLZKW9kog+fc3wsl
fw/Y4G4pIZyidkm9bwujsp76yPQJUfeKOptTJI5UNYreTJ8+m60TfpcQ1WOX/Q3P
q/+bwfBWSr8qdL36B9sLKmPZ+K4z1zLksURfGzMCxP6hcHbjIvo/yQlbcqXJr27y
n4/F1RK5C3h/DnJHpJVffd38KkOcZac61dHL9Rnw6ZdnnWMXrFS5YgTfGsVBjkXa
R7yZc1FBmiFCWHO1wHPcU5V3JEu0QLTeTEgj6lS6F82OTsPG+ipTulIg1dOIVbu0
htHpLVpdkUvyY6q2Yj7cU/Qua7LEeTnyF1tThOHJS8I92NBGX5ZG2pJWnMLmU/jK
7id4oago6MY31/jR+t2g5/Evt25KBRKsh8iILDPEzt9LkO0FD7C4/3Zv4L9pEfhM
7LTgWtDTd6Afbfa8Wayt8G1KBtcvHFt7BM/UZyYJv3EhlwirMIjSK0YB7GOVe56R
on7ICDu5itfI8HReqz0ZaX6w1unwDklVZ/8YLauu9jTCQ99rzuB643bNZwYrcU9D
bcGWgOJajxDUC1eJgJJjLzxjqDmMOExUToa+QfBxoRsqE3axQShhqQZHAl8a6lXp
z6i42XPAPC3n1hSHmMMA8dYW0gowHjKOwkJwH2JfKxga96YJHZEQHHGcCWUnkxJ4
RgFiF5Sw0odtr4zKitnBxjAwiXHKZNefcYgRkiDv5z5Q6OZzR3Udm0/GWYnByUyL
0kZfg/oxKsfH7nnsr1PUfV4Ybt249afcOK6WL+FeSxkTKVsjxGacJy1y4K7kpIbq
PWOR2XR2t8nIUyGWXvM/I6EJhMhxpy2hqfJfVwcDSb4zglo+2zFF9OU24DGjOkKK
Vv9I1ofWwYRs0IsPdYRMRke1qWZv484PlrOcM9W8412wXBM21pyPNofkiamiPwmS
BNluyBx9GEENZPTPg89Zu3FbdCUML9vxbbaX83+3g0dmfJ17FBeAdXdnCdAh2Zw5
AjEvrM4S0WaWRcchVc6JHVF2/lypVQdSyLMv/Ed+zV9f3G7eKK7pYadjZfIhA2nC
dEOdd3SToSJj7JYD1qgvexvtjig6kNVUpw5X7KO4gC5uXLpY70RlweD6zqh9nVjD
l0FArg5iosb4InxfLQaB9681J2oA0A43BooBP15qjo7M/ovC9a8bfF37NBDntraT
2hUpttqegyw5VPHxUL91Jvz/tdmDgYpFQs566JE92mOMy8CmPwqrJHJ5jCuUXOgI
4xa2txVsBLABE0yf9pirkjkC3X4f2Gn7Tlay1RhR5PugX+K9z/UnokOyLOvMi79i
gRHv6ypRn4ZiL3iRcHA7FavPvRM9bZB7Yeweccef7k/oeOIC3FXcBUumboeYP4Or
95xVLd7gE8HGIL4QB722RNi7BSV7Bb0mOoO85QFuZq9Pswf1HRThb2OaD+2N1Nxb
7FjJIJOf2+gYoAaaB/kadwb9OsUue5aWShgmOs2Pk9CEv4zL8ljU8F27XzyS06Ym
PshBiBg3mNdgc3eBo6IosA5VE5W8O+vyjtyBEAjvAwxiF2rZqfN3l4d0toFmRSQ6
QjglNQksAMIOCx9ytqi4P5Q3MUJBukldFhJFnZZi8TTCMxJLBPB9VHSaZBrPtTi5
+0+CaU9OI/pY80bXiYJWDVPYzQfy4vZCxDiRjerE7IKgh1zczFzIRhNAvHIj3mym
tSHJAULFXI5TdH/gBAZH8+wDkXTI9oOqEfN5eFHUo77vIkpYyszp7jB9o5xOpAS7
TDhhMaqsj6oi9fJi2uF0c9cec9zOW1zOBmYEZ/mlSv2Xk4IXx6xFzpBJRk5D15D0
Kza5u3KUkw3pV5RTkdavqU+ZhaNjYB8p3yZPV0FphokCU1cVg1YBP5OVBu2IQBcQ
FZffUKUk0kZMkcZuF83HYbehVXoQfrmLW/3ync9vQSjhoBSe5yQ2mSJANkrx0IfK
8TgIB8tsuPOnFCV0aedUp3Hhv5W378FMV7BIKDQ9mlDbMNpfRSAHZi3t6rutKcsQ
X6TfJLY3v481ExF/n51keKFFDZkCtCjHq4hs8FKCvtwjbcEcjL/+o31LCRrw9KS7
BgUMtbS1t+gBLlkWvMwUNqoPgmIOeHwrEPaQt1UrwL2KPfsfgB8xxEFZJBsbCIgp
GNj8EkBgR8lYPtJ2pdHhzVDQxBOEAKlb3HQB6b+oLfPTu6dsayosSZqkES5U9HAj
X575G8zPJLRj7T3c4IiWplDr+GVgd3iQ/la47U9GColI+NYHl84wXNuYndgbAD4/
HCqdG2SnHI1QtZpBc19mkLn4tA+Jo26YoldIoDZhsFCl4bDvE1tvf9cWPfwygRmp
nF7Dt94BN0Tprdgym1FKOM/5M1QMEOE2zXqjwxt9urBWN59IojpRhwMFQE767dQL
jG0S92GxFRCHEoPZddcMOS1uysyGbxeHtifG/OFe2xErq+7OnKLdGHzEOtXUa0Mh
cOzpF6QzcOhc+RakFT/kIIDg+s5k2XS0KwoXrpwb/DITwFQgfCGXcjZ4cuOUYTXl
PLUH2KiL7yqLkmJo5RwQGWNWoiDsYieUw+np94O3L/OZzMwoLkmxkaLF9qO7vZRQ
dJsXdeRtKjQSfv9BVxulHo/Ft2DBCDWdP1kNXBIkFvhmuNUcLIR0G+kuIp3z/lQT
Iwpr6p3Ogxoca2VOxfYbAeifd4x61By38Vkn65ubZQUp6s1D5yu3jB1JycglTcNS
8WeRB1t9ioxitbtXHKblxrgPp+dprV8KlgwYvVjIVtlmh8FTsRol7hYI8HSRvXmC
b226ONFVsBZC+iaJbcxBtIkRzQbEn++BCwc9O6v1g7cTHrQQPWMb4QHXwf/YdfqE
QmclkQ8tSdnlVxJPjYge8FYtg+TO0pakL429WI4Xaj7Ty8h6m4fXvJV+LZTS0qU5
rH/gK9jo3l3/5b0QEBi7oHbaUTkoPUpD2RxBgRAqurWU4Tlm3wJt+7RokbCw1VBg
/xeVGVQJx3kaUG2Nl1PSO+LWacEe4a51cZCdHJy2++5iQgfCghKQYntPFj0DoZLj
TlGD4PuGhAWkyZbO3RybYBtwemw93vVc45/frRBZ7QLksk+um3EbKSJLQ7Elx//K
FCqaF5CXZ+f8b+rHFKPC1oSZwJq/x9JfITEDZEgwxERTXgCsK0QlE65hCza9p+wj
xi4Vk/3uV203iB5yMyJjNJ6q759MlCWeP1g6uzquTGh2eOU6ptn8QAPH2s1aD0xy
paiUH+VQdFbHPzMUL5Zi72f+XudjCf+aUajx+s3voP0F+2O3RueBDTuWAAE35Qpd
zGJYhmKp9HVxP1qk/l0/gTEL8i52QYqR6LRPXyHTssTe8MOte04gaBjrl0ny0P7m
GKCoYsMrdlRyAjVD6RtAN4czB8NaU5IvQuMBHZJ9Lj0euXc/UltCOX+kHzvEpddo
TXprrOHXaz6/C4KNoSs4PBXaIE7/dL+HaRtQ4eDGcTFhdecjb66rMBfYgQ0PJ1/h
1xXP7JKWVTJmotLenmn8GvLwsKk8DpJFuQiWjJF9Sus1kTlJyBAoQcuhqLUiXsFg
+GTzJSS0y0C8AEVozmTkhyuRwEFYOgwcy0FvPf8U/THxbIXF7tVXoSuGXTRCs1BY
64egkngwfkbuhl3fpMy6WvcSk0gf0o/4Jz7Axbw9zICOx9g5oOBK2Bhy/Q8sU6il
IN82E6i3TxtFWpYG+iLg0XTzOT7Ebv0Sc8slu/IASDSGuTiqCPZ2imdjU5R/nJao
mPXqsfb4esXwnsMUfR9ifpnIv2HCXnToqohvioT4NK0M58A/ash7mcuI0UR2368r
p8LLX33usx8t0c6eT/lcIS7HXm5sAekYihEyUlad510FFNZtRsljTannVDNDtXf7
qdmPbGMqBsuyaFEMkYtVe7KtN75AOC0C3gRVx09tpN/k1RRfztINNf7nSDTBIltc
Ioqbh80Cc3G63PTRDEWOspn6dO2fJywoSVheBAsphhBqL5gRhl2oJ/nq8iqDVY3N
hkKkqsy7NyOGVq7DJn+l18cuuDECadgO0b9QHyhwQAbuxOPAJBDRnCugvvbur7MJ
r5U4qkpUbFnIn/7WjYwrldmIp12myHoqhwMYYA9L/i9z1PZ3ReqJrxjd5xovE+/J
loZvpnu/05BXtJBrNVnWyKWfquP64nz0wg/bIehsaaxePM/U17A2KRbGFQ11gF7K
T316XbawC0rLmxDGEV6pdeWQxgsdiHOAU6bamN1C0GMNWnyKLlVnc0OaOrCi9Bmo
iDDdoicVejxOYGgDad5TQWjTtMw2Z7TpDgG1N04t8wz9LNl+yDOcH6/eWxtEfBHd
wQ86cTmdw0Y6GEo7FNggGFU3RckIYpoGvIHiGxlN+jbAsjPCkPd3RTt1tHNFX/Hj
ehkDiO9EiYmwM4GFwQaSvZMjVyVqM3zlNHls3tqvBRKySJgwvAqIyHP9tlcckXq2
Qi+3xiMijWfFQRMqXJRM9woe46kyS9ASZ1KAFvlTiqG22d2n+QzrawbQNzYxFuYD
eRDcDe0vRH1qed3guTJ8LK9qOE93RkA1V1+5YI/NdT1mIc+YbVVqeXJnL/53LwtJ
KFoeDOvD5+F7UbFkglAq+ZF0HrEY4PlghkraEEKfO9q1s1/0+L2Yjby8ocfe9Unm
e6kY053y3n9RUOp5+oeqQgTVU5Nk499aUCaZZ5gyZ+8GufhaGAe2Tio6gWYf17K8
fLevK939/DvAjsdlBYZvuILF+2BjZ+ZHZ5AjFPCoHeXg4T+bDI06mLgN2TB/0Y8w
AnO1R4+6ZGHQCsHTpi0zYaINvXOB5hfRaKpkm3Mgxdun6/SHZUY7uONckC4PRIdj
O72zLrdJywYP68WO4v9vGbml4QMprZ3M7taaOoz/gT7plVghZ12JFPTpUETOotUP
OvB8TXeuJfHzc2UcbK6oSxQQB8+hyX5Vua/NSzJrWG5RpNSTghsCpQW/T/CqsxLM
/OW9JgE38EAZTJdx4p5Ind/W6qZWlNkH5UL+8Nx4UlMMgVmdr8t5nVzvgKvWePoR
GoIoXP5E5LVWxhNhfNWKYOT2gST6hGw6m2q9YzqsgnWrCNo4fC3xin/i36enhpkr
+RG8+QEkynHGgdWD8jVyRDc65R77jG1DwAaC/ADwZmpLM3gl+Bwcg2FYkg3i4nZv
nDoPKuPU9TzybO2f8E2wa5vCrPJDgYpIWugrxeaSSgw7S9QULR6qG1sbJRp3vo/1
hhmjS9zHGbCADeuQvAZb5NzpdzkMEDNqh8nEK1hoP0sESYs5672Htf7JPXgR6sYM
+R0mgMotMnTBYOQaS8wQqeikJK6augxT9C0YhaBfZMwpqFRy+PPYvCv0M3uDz7GP
MogUnO8Gt5IxMVKqG4+sxlbV6J7MmkxYa4i74RepBVrkyVkWlvX1WZE2V0XUKy1P
QGarBsTNQuaofLNQwT2wINJFAaAeHRWORDBi7qADSjZj2clJOF68cga/Ccm/3jY5
eUoA3Xy6nmDAgwdacqAiy4xtPW+efC6IJ+IvKhdygAmbpsS5h6Y0UkIlWj7pQ94A
hE9mzw6WCvMhJRpqZdJWzJd+XF9OIIpvNAXzujOw7iZPPcZ0PckOrvAx/pfN9QfS
JhEmhs/DgiTBClzXkZ15/mqQOjQg9cbfb3tvPlf7qrLOZ8ZrftEykQW7la65JRku
rGU5f7kqHGb/a41H/Sl8fauXUUriW44Jkp6D+heFCKpOvf21H1WSDCT7ICqwnNh2
BnghIve0Y7kIOJd8qVCCdA0pWKV5FiJs83cmJSVLEg6rwSlFQqq9F1PDgoduqjDy
ByuckmImdjdJ/+6M93uGB4lV/7QThGRSzDeZegkEXl5S/7dWnWYMaHCeUQqOZl12
yOdXCGLmGRg5ebTuQfBnLl2LZE+pOztT8IlgCu0zR+rD94zus6qXLq/Nos9GMnrg
bDO0bheBiRmed0oEYTb4C8f0GJJflSvvx1D2BIDW2vR8jlwzdwA/MHBwmNmfQxlb
7fwlPDbt9Ys6m9K7uiReDaSbskpDmyPAeCYN9/Y5Gh/vcKHpzy9rNDPX2QS6gBKU
e6I5L9Hw4k9sFO30tJcZer6N7mUG3bdNACzwWpDX9OfHSyo51Y1AxTNCK0+AP4s8
JYNhO27w+yrlpyX/tF9WYMYCzUhge2svkPXsbWHZKSsFO5XgsQ2Utgvltwqf8U+V
CSDsepUalS0V8kT24qZYZgsi3bASOkKCZuxRCIagzbcQ/l5ZqsavCiB/08/AAQAK
JhCzko/j5WT2CpkotJpdJp43CPnEa0+7g2Jncy1KvQBlV+vgvG2GVie37sGJukLJ
eRgpnDbN8vu8bOuJDRvIqt/Vf8AmV1MG5Vf7XV1BB+OVQdDBHSq+JvcJkA4nCPdX
oZRu42mFuF1qzNwWt/aCtiuKwK4M3SxgdY5+6jmYLSj5911nxdN3tI8vwMiMIUB8
YSZONrywhwioh/VnVRnrDcah6pULFvUn4X9x333k/zGDpi0Mi1+1ZAfLiP5ZsYiw
pd0PmibfsdQk77xgpbKpGM5OWPNbEtBXqWAYbIG8Nhz1uI91640Fbqd7WVe/0hce
7AMgWi3efKPLezuwZkD4NJMl3LTQfFoGoVsh+WEF8fjtgEGZTUXlpRE+U2HWdiql
rm7CuXvf2g1BxliHvF+Ef2KM4bTlWD6rS2yE4OgpKLTQnzyMwp4nxIRQFCxCbqzE
qJZH1FHbmIsw6ytNnLJG6OCky/xS7WO5eB/NaKiqyQOJnhzddxXn+6FvM39PSk+r
ggfY6pJCFtgrfNjPz7VTd/o2Bujryffz2bHEp5CBWuYoJmxvwpSkRoSoSEzDEkvO
pyTDxb6H7NpnpipsC2+i4itlYH6ZT5PeWTdDFTknGYSzUV1nwqba96IGvzjibiNp
koaZlYZfnWyr3I197HwJ5ptMM6pH0JoehYizFyCz5fJ/HPR14MApokKyBPu5H95f
OyclHundQ8qSRZ0JU5/GGgVZ/AcagdyHslGgg9qGPMSq39NHMmcNv7wVlxs1kB3m
rbSy0isqk1B7qD9hOSFJ3cCvz9upBTs5gU6EiSvh3r2rvK//l2ovgKQy13sw/30/
dSw98lgwZHi0g1CVpp+5iku0p5vj/zta61J+u3P317AgfxLvCUk4odaaCseb8izu
ncO9NYExB9yodLEyfmw78u5u/t7w2Fgu4B+uh9ibQ9KGRzxKSWOZCLrpeCGqfLYl
Ai5FyOapEo4D3M/AwSK7xObeTi9kLyJEYubXkH0jx/jehmFWlpWI65bXrlLkEOG3
Fv8qN2dl7THAUlp82e4vpEOpQQIo+/oFpY2ycjoDHsVxl1xfH0hon4wmZZ1QERki
GRWVeEWRSFWo7atqOyLn3m6qx4xOWPHcq6rfEmDqK3UVKW7I/QU3ZkcjSute9H6N
Ultn8qk7aNDDWFVJ/bL5LU6wZv3AfpL5M9/kOgsX4XAsTmJb0t+OfiViWrA4Sv1L
SZ5OlfIU4RQBgrm+HDMiy2TDn2VKunu1gwhvVtsEiS1z7bqJatdt8u8KvgOH2wLv
rXyZ+IGl9FX3IeZSwYCYLR5xaYW/LxiVMLHxj7iKWlRim0UMGQf9Ie32hvhCPV3n
8fD8DNg6tmF0/bP6cEnw1zCf00QCTunwW5ICkzh8MpOIJ825ylC7AQNQhody/0Yx
UZ4X4NqGfkJ0DjDpZgJ4aIqPcrXV2+7NskXaQhaH1GkXOg7H7rOhoYB059ZybT80
BFuE++urpXuDj0b3dL7JdEbXXhUMchhZ+zfgYQIjsxqr3twhsiV/CQulVkn9NJUW
RQVy+klUBAcdFd5vQV+7umNHrbYtc75VPoOWcWlKJ0dRWin/tIoi7Ehl0vEEV9bT
YxwaMnGj2htZJDANOnGkWtOaTR1eddEPsITYn1zh2T3B/eT5PxmBoooNLeznOQPp
ZE7/HvRKGsdHrxvwY829ymcjQm3/qm5tCcPdurkBCYWARcnc/4V45SzzXeeAis5i
BDa4xH7ECsHmYpf+Px9CeH2m/8AWu4H5JyMtLOnDmKEL0ld4Fz/vrPTZn77wPiru
2qjV4wZGM7vE7JDvgpevumDdlE2nCbgWlk6vyf3ftxcJUuGYibtJGe/b5ICfS+rc
f8E2aDfzW39AcD4iwERQMYcr0IqMS/ZGFg79ckMdaZ2R1E2odQZBHCVr8rNNvrmc
5l8awPL8eoCGMnlPXyXM8rc8PZipkyKEOL1PInHzwqFOnhKgtvCGXuNPzwnTzG6V
sRycQKzm8PFaSeRJOlg5VyLpqiY7GZddjcEmd7FDGzIoU76nL/8XOoPGiQFCQgQ8
Mv748NL/N/4DN+0QaS+NwvmDvrZXtkWEZF1lchFGBOo5d6gb41AWiXnOv9V3Js8L
1r6BMQ/fmkUUZEnT3zDg94DH3QGMkhXcwoIFM2yiji4MF85ZqUFw8snYFZzYM+QH
wbwszXtuwfpj5ATcQJILBxzszVZa6VyFnyW2hwgWCUO+sskTvtGHc/hA7KW9Say+
Q+32agech5D3miLpRJUvuOxH5Yy8LzP/oEiSbu1JDcZK7flP9gCgtxqzvZaDJJVh
YnJiggsaH8oppDkczmLSbmcXuR4Y6Tlj/odlxvBYDgK3DH5LERjwivjTMifa/Woe
j/ol7R9SH8muf+9alZEfijxc6m2uNvJMmtVe8gOpmTCKSaNZ5hTCc5RzqmWrsNEi
8IEyOsfFijt2DSqsFyIKEWBQptrNR7XwumhFnlDIq/iUfu/pmrd3uMjzHTq4mvQO
oR+eraOevVWGVlmXXbVZJoMAay+aCWP/YdLXXYNImit6qoBIKJxefd3zTIqsW+iN
9+3G6JgMy6n+ivGIGb2eYo9RZd3jy4vsDs2wfK1j7UX0hT50MDdYri348hPQGDa2
ORgY2OrpWshXnIJYW50Gwh7KBSs4IN9kd2hX7BMhlU4LFhz9r3ww/xPgzNQ7aARU
htLhfjEnwS+lyJDUjGQB/qUKbZZ976f/fcPzJnX/m/6lGBLnEgFxY/1DqM3C3cpU
UZ3/zfAC1MZH3ip8lPpYZOqyU4z+62V5hwVQseWqDKTI/NTIi+S8FTAXv6ExKlrK
L2OQkUduP1NmjlFj9IhlCzze+0U2syoGtb6kTeRzngrzsrXib/LV7c6Z+uSfYW4y
kWlGYpCNWe52rSwwkTPZwH2bHczs9RUIiqz5zOSLP5yc7JoWLwhD+S5A8uBFGcLT
RC2agLEONNNce9aU+ROvPbhwNwAYV+p8beDTwb2bcaVdflmhs6DPuZm9P40QvAeA
9l/xwGdn2L3yFVK9Nblb/QMLfaeKC2nCl+f5CTKoFxJB97pMnx7b1C7Lm94RnJU2
5ye2qmzdMA1EcK/wTmH8CrjzbkcyOsFta2DDn9ldx8kEEEKq3DVcTA5Z22J4K2g8
suWGZ2fiEnZ+nvDLNFWHw+qFpCTE0Ym9+7aRjRtlcb5N36cW62ORQ3nq5u+qD1Ie
4DG+17sVmr8H3H5Gbv/fx4C7QQEOzxuV/qv6hPLkQA7CsbEN321BcYA9rgZSap5e
pSmQbtfd64AFz8LpbOxHg6GU7iLQlKhI/lGAxDzSn4u3eBV5XYXQ5w+xRHo/U+kn
tsVZtKA7ubaJFyiWKlziJys7GUJeqx3wvNqKB7tQ4tKPf3CYLH8O6xoMYWvGEg1m
ELoY6UdNd4KXL3sKmnoa6tLKmZEsIWV+mIeqxzxRBhLr9l6U+D4mBprJPckT0WhY
uZ/+/k7tx8BVHbIuH84Z7FS9YlDJfIbQsVL8r/nQfei8c1KxJsSQXJ1Kv3c6f6BG
H9p9bolnhCOZf9RqoRLQt2UQ9DDgu+js5+sCjtXEuh58GUaA/MmMC+HRDDgcAZC8
o+vTWNaQEv6r1QhlLOrq8SVi+WumF5Kola/Vl4I8z1GTM5XZWGr+xaK6OOQgblO/
ROFxnyCySYLUbDqvZG2UScE65fO6Zshi1jUAXj5KQHRXVHTw0hHnwDxPtydX3pi9
9GVGm+cwt3jopif6+64Q+oHrJSg/EcMhWtLakQ2IuRZHEK4ECrbdgAYqST/bc5LG
6X/M3Qq8HfFVkGlwOEhkH0EZuybl5t2oEruT6+4ESOK0g/I19g3l2cNsaBJqpF5F
mtxZh7/qy0ZJhudS9CBUw92FJpTi6R0ucS0rrHpRoLlZCPdX65YIyQzfzkj1vvlh
atHZMb79I38Fk4ypcHOuX4mZD4jaqpZVSIv3vb5wiTSGeffHSRL4295haf417FOo
K6dCokFrE/lGyzK2XA70xzdTpsKYHvuJckssKm9TiyYs4Ux/uY5NSTELALhK5Iby
KJ600+neEXyeJa82V4E9I4kBvt+0edgXXy9Jpryi6H2tISx0zZUIFspWtfsWCcOz
EAJUKAb50P7rYf5rQOuB7zzpuUfb9jHymwL/218wCvUDSIC/v0Qme9vRSWzT78l6
9AzboawBX8UjQi/xXW/peOZjeVMadN6F7g1iPSZ2Jo2Oy3fkLZEcKzSd+0pPJOui
i2RK5hjLEH75Ecxmh5qO0fvZD86A5BfkK4cvmqPaL67CAWCQg36FgTgyzIC7t20a
ckRYwZ45ryhfha8QwBnb0RT/ywmMJS+pXHLvigkl299w6ZyWPebB+1l79ZO+IMkJ
MPrjE8/XKxRb58RNQbkUoAXSumxRYC0/criqZdYCm6aiYHYINkRdu8sEMeVW+oxZ
+FucPaWAfO55pCQ67OG9tugHUdygnr32X56lRlMXMg6MdMgGRKO/s3EzJanR12Ge
V39mKEUDzK9XbKlR3FU/kVQDS3/6gVb7UfeXVt01rGwzSosybtwtCCzx8eAe4yOB
iTFqfoRR29heyEF5rNV2uyUFsIOg0anJ9rP2mb2joT9ch1qRJMkZ5mJ8Y19/K4i6
JNPck71XBF/o3ONEUpzqCgEW31Ch7HVGl+EjRkKByVi33Yb2FKKxCJp5oBsfygPA
WXFjtY8fnj7HHdOG1ZXSPmJw+rfHrZuxORfOZIGBZqZ7biF2IJPSye+C19WwW3de
Jwq80VqxjP9FNyHXxrQ/Cej7tt+taZL9A+1kQWEsSYE07Yg6SREb+e1WdRPIr1q/
tZo89ht16ZUdj82b0nate8SC1u8WCVHFRXRkCBuzx3UWTmL4ufqzkk5rNPBenYrT
o+xDoBeOG05U3pd+g74nP1rJA9XTVIIJ6CJ8BndDtE/ceKnVamtr4Gzzm5PzELo/
PVmH5Fmx7kDfNMbDrL16xP8+2gu7XB/MPCmiaHKOCEgh8kR89H00RWsbN7IqZ5kN
HijgiRMDf1JTV4R/ssEpNzIXOum0/KDD/1CZ/YTxZC9d/Ncv7jhdn1Xl16HCzMnL
/Khk2C2GgrH7ZAmj7x1Ysb2mnbRKQRcVeVur3AIhzzTlRmWupvqYoeG7OWj0+1k4
0DpzqBT88Ih6XmBYtXOLBgZyPvYuU55ZbFg9Ys08C1X2u+0iBmLDnNu4GhDqO8I9
LFEFRBYKCgchmDrEJsDMvtg6pBNCKB17ha3BygiEiE01BrKHqR8xIDSmu/I5+AtA
3hndGYPZWaiOiYam91SnV5nWjwwICnQUAXKgMfceKG7UtqBXsn2VGl4/d1JfYpgw
TgF1Yb7Mv94JnXwaZ8A3ALKdXPHxxihuEWMvjK/DGNcc7wNoUKhN6QxSAuypjAZC
c4ehlQs0927EmpF6CCrgelB+0Fom4CHJbzX57VFLYwWycTy5Q2t19c6VIggRZO0o
2VvUBcIoi0hKVZX+BT3I74rBOeHtrbE7aDVQ//Sg9R7KMYFFab290wNsx+G0VFId
jMRlBb4ie7Y+7urDYFTalA4r++NOIPUiQa6My/oStZx61veQrmFG0Wva7hA56/BV
sJKRBS4rB20A0gvqpVffpGoCPn3g/qM4J8XB0z4x8dFEBzO4Eqo4h4w3twCXmMsb
J30riz3KZ/n7h7l3iafaIItS4/CFJZcWvRrudE6kxyMLPbo0sIxg4jehumd0yIrX
19j26Ek8wpnvjN9qVko2JycXPCKMQHMK6JSB0pxW2bSDQBfTyVaGz7ynjxWoxPlF
F7LJCl8tslEoiYcFmdBWqSxsJW9N/2G6zfG8/wKFFVqhrXC5Xsv+qkFUbwJnEvy/
hNVEQRvIDkZh6c5cH2dnzGEZiNPxymK4zMt0TcpAw/i2+ctT55r4janB9L37vlmR
TGLzhk0pFlLXcRbPEe3bIrPDGKey6EpegRuhmxn8smhRxmsMK8uAP6r9LNtSeL5U
49HQjON2fEfSHOfQs4pWNKQiGeasm2dE6+yX1Y4W9u0wxCvgnHNzgUkYbkCtBQWX
CxJJebONFxLE3sqJajohE7C9ML8XATo5wzES/mcbXZ5NSR5QXfyWL1dCRAQlzd2I
Ih24HxGifrPnkf8G8eAG2lP7j48scZx1Yqfvp7xhqv3KspKWS0bnTmULshd9ofUJ
/CkIBUobc4GJBkT5SWxWVQJkDAULszngBsJkUH+N8Kq0ex4F0q0dxwdKmgE1R1YE
A5pKaWy4/lk2xhEBc61nLoztfDE09GUYxjJD4GiXpVJA+Tq3+QqYUo9bq0ksFyMK
Emd8JtiM6vDearrIF2QyvYG41d7xjdldzYe41dHoGELCamOaQj8UJL51zyV0INjd
GDYtKUzI9Z/Qb0mYiLCaF2Ihocj3mzytgR4Vu46GTn/u91kUGokYxEHbNUywPUJI
OKeM6jjDyA6afb28O/zn4f2KSfk+gNBidSadZygTt+Zu0i0557fUdFAW+iBomVl7
ct+/MSVj/2E1FTpWPvIHppQIFSMvQiRJISc2PH0ccJPDimQPR0494Y1/63+cGvK0
wkoNZPKzbUzF9LDbpSBukXZWstu+6CFZeQDgHmpaaqjAP7UtwmKf4/q5SkEJ7wh4
cVDBrP1FQlYE8ey4Q3I+YoOKzsl65DW2nlRhemaiPNimHZmlI34XQkaogf5Pb2v+
nbXYWyh27llgtARpRHoSqHgiupIPVZuCqrk/CqxHiQ1LoFV3ALJsIVfl+GAPOtPK
xlAtmt12S+GKf7WVGpBnJ27ZzfZp34NXljf7m7Za30lglrV4TwwoD42pUCB3/HOI
4cnm6LwMJC/NO8i1INACuLO3cTnbNVqpIorHlW3V2dGG1OEOSFsFSUaFms9W2Iw/
nm3INwMvJZZsYHbY+c5ovfsBVvCltzOVedyjh52ytwUSzy9gJ/iY+QBlGy4T62zr
lpWQQxCUpZforbLlfRmOmScKlpdXfPfjf9grfGi0nU2bUeTh89NKKntnpJ4vSMRV
LKNpqDe8mGpBqpb33k9hMHlQ0K0y2jyG2fRCiKWuKfst68TDJe1EaIeseYsm15e/
1jQKr9WkmaXMkA+C647RZ1t4IXMtrcAl12YbH4SG/DMuwJ0OjqARFYgsoKUTPb+2
exhLlONmvI6lOixOnzfY2BubUvMwfW3jK68Txw5fa6nNr09pVX3/EiAwDaxQhSEN
hcYFIFKoE3LkkctyQ7xb+nwMfzqJlh5otzjf6cBfxVUT52M2snVDExjum3nZ1JQI
9UYaC3+ZWh76VYB05JVbzFXOs6LfuFEtxacbzPCGLdCfoDIwdBtbyvgCXWNAmBtv
TQvnZvt5tj4/fh3TmuWNwCYjdv2GciVfFikQKycNOecd+oSg+dxDt7HX+6ajjWeX
FMJvnaa3TmyTxc/a5rKkq7jrzdimDFYNW4n7JajEyhIJGnV2dkqk9jT5hRiuYwB0
GFbNXHTl/PYFxd3DSRmncIOaRYNbc7IHVi6UacNocrmqH8T0TS/oBNzdwdVUL6V0
Gt9t42wpBhTMqIyK8ELrWmg4W9lfj4Bi450YoYUNRCZ3JpMPkIEMYcvyEnzadNWc
C8ZbWOLacrgGTCHJ0/85Fv9mOfiS/6kCVX1I15KX9jeG0gGQqS9Nx2mv6IRXMe4/
+gIY405hpAGc/bvr5JM2uA7HnkQEKDk8aDHOvox0R0IfB8OIHL7gMZN0qdeMKCtQ
frji1kKdHfas1a9eRiTAPcA6NPF3yZ57MVO8MjCsaXbV6RvyQ/5W+9RPKs9S1ZO4
09arUPwe+zu/0argmtT9jipaM5pAKWxX1sLT2FZLuNnrqnYgKZM+Chkc0iVs4KPo
u+Yjp2ufBxdMVJEFUdd3x8gDhvk+LJ0sq/FuCRCmpyUX3ubmvYAl2z+Ct4LZmvk2
ERJPBctHXNhqyJUYuS6y0Tg6coBT9eikEG5zeuh8A7nMbPZBV+VWT9bTucmo7t9A
MpgZrjFS3F5FcFxMOTey6snUJPjW0+IEbe1DDpxyZo6fgtwoPMLURYAw5x0z7Nor
Dr4G3ARBMRX4VIVf/SCS33o3NCOrii0XkjMVNe75bC28kF0+ocXXzmFLZGhecjmm
aFh3aJiANTSO+vdg+cVtveD5ylf8tiHK9e7olkClZMafo8UGOXiV5kYbv/WwOgHP
2yKY0nPhTV4Fg0Cb8lEfYhpspNRX3hhY04zfZK2xpGEi42yyfTOuhm7+EjTkC8YA
gx+0zBL3AFMGemsTiBzoNHRoxmjTNo0YbwMMrO+bNx17AFr7wQO6CNa019Z+99Ys
+zxzzaA1BG9tdF87RNj01cEXiLJb3Qj5THS9flDTF0/nSGNp5GUet0SCXFqoKlvh
s/4BPcGDfjzwpQC0qlx6PvApYCYKB5NKJJMVVsgTuEzTZr87P8eQ6aPMPMx4GYOY
NvkC2TbZXeXuaFS7/bcqbanoAMJqQgfomfVFf36tX6GyyeoM6510lHAeBQqCtLBY
OH/81fVwpk0fIxncoatIfRsrCeFEPhXqyXI2oJbGGd9z4LGUkvIeZuY9BCDdQkGL
UbLNp5go/2u4VfJIaZT3XOXJM2b6/oPBYP/i4X4awWYJHJ5F8369NjlrijoNdsTa
xppkKDxPFcmBN75JnMBH0AQWn4XiTPPjdabhbGUpMQBUbHsG5M2UWjs5yRfQgxBj
xU0v1VeVR0hE6n0SYEHkv0WloFivJtPmzTfC5kdec4pJVyhMw3SqDxaqsj5Z8fma
B1HVgMDoGVV/MmtNZVeUC2FheJLCk7/voV04uohIeL4klseOySxO04R6/4NZvZtG
/x8yLz50R3wNbjkLGpw+qiYMtTPZvBv6lgSE/DtOf8KSG4e3YqMesGd7LS5Q1frR
48jdmhTKatZ/JFPuCZdgBwSlGJIKkjOPvaTkDnew++MkTQke8ykDu9LTwoNo2qCU
43JOL9F9CmAxkKgm7j7+DZmj8Xu0eO18Jm15ko1Gt3G1P7LEeWF/58xJmclug4xn
GIHXI33sp6+LjSuL5nomuwF1ajlRtsaxsEssg7lLuCTMJcdj4OX4e1BZesyxHdzj
8IvVWCZ0CqpCQlyNT39ftWrzCwJVWgXjg49L0eyXfSkZ55AASYZr03X9YqwOj1nB
j/utSoefzCBWTEAeVKJfRzHfxjO4G1UM3OkSgD6KVTK+xhjLkBEXDtRx9dqYX0Qs
qI8m4Q7aYoSXiZouIFOaMcPKVn1+3OspPwxVAB1a/ANTK8Jf+7r8zbDetD2a68Rw
hD6eaNejYONPFHjr2cXAYBmZmwkzv8jFbbQ1PFMURNlwCt38pJouQiXXkZzCgizV
wUdVh7fJlpgz+YIlNO5SKH/XtGrFepIfe0Hcba9DwboWbUsOgYYajsDY0OQeWBPg
pts9qsX4FY0T/lrM37oTrKAJeh+DpDhxKSKtXHbeThecN5mifEXx7oRAmd8NS0XA
PcZaSNmOSMkmytPDgpqBSc8ZVWEVUry2VlOm7WynhBmIDfctgc4IFyRlkZvUDNdP
IBdFCdOeWkdYt+1qV9Kpyt68fueYRuE9rgkluCNdaoZ8sGMEousPMNhSG9OBtyZe
+Lccqt4ewpryC7VFF/a9CDyAnmx2sFeZ6SyKv44ZUWc94v1g8FDejXA/CAItK73s
5bSr58dMg6H1NZpX3eyC1YaDARJ5HUoKl/BD4dkGQeg2c46r5Dh4zhRlpMK6TJFI
oWQ/IKVHNj6R307rtSg9eH6Bk7UF6MQmS2az8KSD2U2BSnatQ+vKr3x82/+JvxcA
v88lYXP/jaHFhZ8qU0xuGBfnPq5gALnVJUAbSPkDiLPBQ2nPDX/GJFeCKIE32VGe
fBSP/c/PFcVjxnK+yoV2N+e5DJZF5DdNZxSIVZnht/MclnQIrzfCdfAhuDqX9OCv
pFuudJwDlZI6nr7cZ/6j3HU4RHFUpOk9ungUMJ6seaIWD/Udubv9RKGqTW16buU5
LNyaK1xPPu/i0rF60EacSqSvgJsti/1bzgTHqiZbhbqWQvY12ekmeuxuSvacLIXE
fCyERlOLCFi/D5cJA8zy3IoVRWAIPyeBHnL5nT77Nd1p6PE5Siz8Ly2Eiv4QdLNd
oUh9nBySZLhUY4qbkSAAZkn4SdgM9tHxGaI4W1sE5rT+InEkWO5LRPWXy581xnB3
UmzT3ExkqzHGTX1ZbVyDyhYL7X71y8I6hHYah76X2Gi6COGA/67dQuts8C6jjj1t
5SO3b8zP8vAnCqe3HZopcC0JhEb6z2duj/8Pgo/YS/CGRAzZxcLQ/XZvTaslboUF
sEMClHFLX05yxPl+dfwWGsGnqWBVxzZ5Y2cbe/Nc8et8TwVPoB36GLquWof9giOn
Fa1eKsGg5ePGfGNEmiw6o+H71oOl0Fer0IJOHLGHoIkBJd4O5LGEipvKR0xXQDNe
6x+8qQVB+3qlo+p+IWC9ovuk+KLWbuwbv6rCTKoJD1NH8eK9N3T3vW7ujtchFgo4
EmiDzwmDBVNTzhrgaNYIemMkeMHBc/1PtVBwGYLM6X6Q2OIfoI2DIALgdBQndkBt
AD4uJkDNpDWS/2Ow+UkTF0mH+uJZzrlWNUWA0nub4jgrgwi+l8gbvxEdvANQuWOy
FYoyY12vUrs9WFKZ8OCGZfMQH3pbdECEJEA4xm5NnZ2DsCV3R8RyikJ6wofHZuM4
y6pF9uBbSkkcA6lT5HIV+xqLdS0JNVzIjwBK+i5QGIXAXXN7L1ArUoVcV5Je+LyC
zhFbUwjSgPLGqpsZoRUsWyweikG23pqGFNUmw3CvRJvSRk2VMR4mchDRywQzU6r0
R4IoeN2XktLFfnfR/4ohlsRk0Qc3rNnpFFMtjZ1ckCx7K84OqbVfFh6FqX7UeQEe
PEbz/slpTooKr5FzOIHw1WKd7YxEoFLLggHjB3jnb9+inA6z5U85va73HZE1Lc+4
ZRbFreCMHFUMmlq0qinjNYGXIaYyoMZiJCrZS/LRaHzQU1jQB1WXEawbil0PUTB0
KyAxpyyf6fQ16XqjPttquY+X1bIQq+CRoo5vqddlWpQvW9sct/K94m+EDPzac2cn
FZDxrlZmRi7f73V4f5qnXJPulXhtNVolDs+OglNREC7zmFYzJEBVJ5idZD4a+vvY
W2Ik4dzb80lFZGN5uhZQA6Q8ECN6ZNcFlKNvFn+OpKKqLNkfLrBaJWrM6ryVvlrf
VmZZWQz/TtlM6JvxpO8v+VpeDhX5+r4E48lz1ewUgUbRs9zoJ0af1C7yxcsjWOwB
WhRSBElWh7ow/O41M4Ffy55+AAo538DQKJedjpMP2K1m0yXVi4UWkIhbIulk9HO+
mXU+8cufpj8DqB+Bel0Z2fCNpMjFOcNKImUIXpbW63C6lI46Lpa+EP+B9zJ5t2iX
6gyLZJDEowz1oGSGEmMaFUl2eHTG5OeVYaajMOeAEPw+FHHNLf6na3Wj1JXHiFHl
NHoHEtuFz+TBcFmJSFY70flC0DayoKuPX3vGUgkqdSPhq2jYbBPyabRswu9zKPIr
rX+QmBIDgRJiiK1YHUETDmRUlaT9JaNEPpJId3sXB4M2HMXoShCMnfoYRhC3T+yk
ELrMVMp/P7eh+25QmRh9BN6ikRAJyat5HK1JcmrKKCV3ET9Kw+/h8XIfVMZSVrUl
oMWXerUusyHFe8hoOeMnSSs00XXO/QOLCbPeFYYVPu0ctNTSaMwf1BGkGA9GOu4b
zU/lfdwKWxcrLNr/RNGXgGX8opepUrY7GLAArAlf4n/El99BZubyzwDmtOt7fkU+
7asJp0T4ii3CVYS9Eojp1LyW4nNLvEZ8X1YS7ccHFcztaOTTFVhoAZRbGvuu8prW
lkQ2qmlc0AQ3f7e+wmqvObmUZNbM5YSWxmykN2pRtYxLaC2rv0Dd51W0L5S5K5ru
e4Y2NSoz7MogPOnX/TLD8XZmY+AH7PLO0L58KQTZaJIC6oyY3EK4lKk5n6DwpagN
tdKM1Qb4Tr9K0VjKnGT1RVLVmmeyJgmIRmPQ8t32LPzcuxe6HrgERRl5Gy+CCqgk
D8xcQLcBQ4h8VMJAWOoJu079+YEfjW+svJzpi2JGCdzZFuuMrU7RKYEmFGyZkhhH
B8HjBYXBlP+Ml/7BA5NzTU3DdwOitBmZ08F+3IUha5lTLKstZ6g+7r993sn+TeZV
N/hzXoVQMWcacg21g9ffMD0kW7hpd4yzPLj4Ari/tTQXJgx2K2+dZELAtXJ5E0g/
6O+u8gLWPT35bugLUYM4dbciIvB8uIeUxV/rmUwHECAVZul4bU/KL51cjn6E0LMF
7YRGd4sixMyhOYo4zIYBrwvWawEVJMpFNHHkmYssuiZkPIcXMsI4ihWiB/5OzPoU
aSPR/X9a348RSycg700FPkthW8nteIXiD6J+CITucBKk5QLxyrg69kQy+WP+wvRo
ykaMMSUmItWLZZlhkOaakGUY3lUj70BrEhrI39yH7pVWGR/8TRPRL6Ue46GSHjgx
YHe/TEWsD6jXxq5ps2ZJoCfwUufUKmzVR+/XnCcKpHONzIMnOQBMZCNHRaPOM8hz
oUXS06ZtGeBwIYYJEfGng8VIzDf9Oc3OXH27DL2pm9bQQtAEElBJRTudhUzkWEjP
A1S258zdOAFbvtt3nz7c94Ul1RoeeuEI8SZo8VHzkyvfUqfliGAnwlXJ+06PHpcN
MMbs2Y6V1WCgOToqxQJPyGJeqykck/zh+/7hDtFNN3WRX/VLyoQ+wvifs1KBzzUH
hEWzuCpYyzSZRdlfksI6Y90JaTTh1695q9ZYlfTk4FsKzT8WBF3n4vFiU5gnRaDX
5FgGynMst7Ss83CNA5SXx3VIoO2tWUzR8RIbhTYRyCSO09B6ZZdRPbueXC433YrB
fK5WZxg1yR6H8ybS3oL0Bnzsc7wSM0IIIK4pkRgXMuqdEFfEPR1QUm4W4t2os+Bi
WQ1T2gmmmarrhwmD+zrQDM2Jv0nSc0uxqxK39jDy4U+mBTCYSq+CpVauPoCwVk1A
ibam53GNu/fGIFB1GWhHASLc4GpF119Bf/tBLy/7BMSosFn/vQUAo7jqDlLF/Wtl
coPui+zBd5xl/PfuahjrzfZOGf6H5x3APrtLdZk4oFEno8eDiDGCmkfugVRmQLNA
Jwb+3Am+N2T9ZCeB+OeL12ZsFAhC+2QC9O8Qg6rlNYbnmAIqm/SnHM5XvG0DoPZk
WL9XeryZ3wtg+nEmJAxwDw6BqpByqWRqD2bSNwRnn1X8pc4oJHhhfb8PtcIqu5cK
iwhjj+WChoIm3iFqIaBUM9RZk7nob0lPKKIFcJDzqbCny+CzRFFNcAkJCUeYi9b3
c2UXuOMXlBxSH4NF7QqR2EtNEw4TeEW32aRu1px9dVA2rS/SXH0XUwC6i2radTcg
fTBMMafhBYSc3XsmwfRPaWQwqXXgZHwcrbh01lSB9L7a9sdhDLxrp2KTUSg2meHE
cFJlXthdfaRp7XTK5zoxl065Zzgh+K3GfNo9dTAsHb4cwX/oRCFSjJHIeBXOwGGk
+AKYQvgTWqRAZaxEt5SmGkvOritksm3mHyrux9mzZ+4jWQ22jMTf6DZWCY1NL+3Y
TIJQaAOcEIdZiAFTMULXXIlvmX1bM7gcjTajbQPfedaB6BGhhZ9EJAImJmyTNT+/
JLe6trUqNsFTOzNW0tkRdo0xkraanONEv8hB9HXuDRBuNkRP+mdopp9WXI08N9XQ
GPk2eWWkrf3FWCca8750FoHSyYTX/IV+s45VXtrigkSJ8TNNaNC538Ae5APqYT58
9f+b0EWH6yoxkHXIdhdIyBKBp/qrrt5jH/z5WeghOBpYOLulrZfWyHjVRCYYnlHZ
QqwPGj3CID5Xgc8/nR/Xoq9xubuKDPb/OzoIcSxm6Q8zgK21Jy9VeRoYpag7R5G7
8uRtnJldltbVuUob9BnmbXDpuDTaKucxAlKS+jAu+Qt+D5oAt+V6H3D1+ld3ZnFh
ENNhJjtbFDrj+/hYTSe6wTF4fPs8cEnPT6rCiJj7NhPT7am5Y/mc3+tO6hC2aY9x
e0X6urpLDEroeIjC/jP6yzHzfwYRv909+1s+781ZEUEOCfps4i9tbwyNax3BHXIE
qqEzFOsm4w2JVKtq7FNPCvDoK1Z1zCmIMWawdttxpprUI87RUvm4KiQuxt7PUZWD
j83FPm7VS1OesMUimDRSoEkkKQFEpuLpzHfPVLOfMzks8O3PvO0xqQ3umdCUUy5e
65mFsnr7WBk3AHy6AQkumGNB7Bb9ufYpfm0aa3NPhypAQVfjavcWRbI+AkHsv/1m
boJtfQBrp7TmNp68z+oQDz2uSIJUaIExryLU8BkKxesy3zN8ERQ0AObMVK/6FPXt
afOKZLrYXUMnIGSHDShCzJSDsh1g479FwrnJGmC3Si1QtaArXZdLCumO9/+N1PrE
ApEqpbthCM7QthqyUdr90DhFuj+hJsBO1Sousz/7w+hjzr04PmDqh+03dnWpfthO
K9tWw3rZpsXX9ftGC9RD4OoeJD/oAdYMsw4zDNpwCKRTn+e8Dxw2tsPSW98g5r+W
Pd0/j4WBIYdbasebwDpcQJcrNrNVuZwmmXaGd4GO+JOxIc1rMrTWzteceyJYT0MR
hCWdGrUJenhkw5ChXRdpt40aJXmfinqwTHaXhTHDsGQi13oQTaWPDBQ5UeT1UP72
nYqdSAe07RbHZdlsMwNkZZRL+W2NpGyiebDPHDsLGcGJ8lK/1q1zEY2zbLJ4gWv1
34Ka6Y2BpVb530zFxPvB1mjfs3jkSTyAplonjKSqMkdR2woHpjUHleU5ruRBxgX4
liBDsGxAqFlQWbs4kOBUttPCgUlI1dTZ/0bUhCbdQk6plVNxEJKwZd4mNPGzvjbI
Qw96S33x4FYiPGqmHjvy1GXdFFwq3MgyhlLouE7fDQ+iAlN9Vbj6Ry87xFEHpZuz
xzni6L2vU8CGejiojGX6pEX1WOJ7x74+Oya2wBrFaDiof9lUV6zJm8lI6wYIf2LO
u0H/OHLypEbMwXeCOOquMfMWOAhotjYB4tTP0G4k4rgIqPEl9rhNUzdQQRqJEEjb
1U5LoVszd+t5qG1zPPSDzBhQS+NQNzsYYd7ffdtmAqECViT1dKwEj0Ilu4bttSuO
Cey1xig7N9h3wh0F7iic8JSasBggnZ+m3ndnqp0z9JhneKBcxMPTjIgh1lXGvPl4
c4hooBs1GSoxv/K4uu26UkJwgFEsfe/hkwOVZdiC6VhvVERngo7TcReV4N9YbaYf
9KWfMPTiN2ERLrSCH+I9Fa03RA7X2S8HC9WOzkNc6G/kEpVglF4+/u0985/xEDNn
//phMhYLl1XSJNMb2eKfvzyjrl7fR0dmDhIsteDizFQPi04W9SjBwuSg/vVA0S3P
B93X+ySlRLXvOFPVVVyRYh940h6Y6ZD38Gj77GX/x03YFVNmaZLNaImugSKGdb5G
UDsJPdiO0vuk4d9cCETgKD+ABxMq5mf9eBs/xjsFpNQnlKlw9QaxFnCbXyCpmVA+
MoEr+WtGvdN/gnHkd90XdDkazYcEPtWBBGVcLrsN/VrIjeVKX+tBaOiQ1xpJaDJu
Mkqpa/J1d0iJMTsB/8qbJPL/IzLRsh5yNh+vvkaUm8sqxuZuwgWsczeKRrI+t3/X
wleSfRXvoKG1Uea+CC3GIArZALBOzWgo5mjfikAxwE98W/At39TxjggwyB7o03My
BDnogzMIuuwW3IjsmhqRfdrNhCBKGyTW7HB+jslvW9Mx04A2F+vt2TY9LTnsQ86D
ZPnrie9GY1yz+OEXMTTc4YDthIIPZAU89p3QiThz9N/e6urF+Q0LOKLmTvF+lF+A
rb/3V4/cR2NcHiUtFvwf0F0aZBiSa99NMX+FatIzawQKcD8tZCGSYv7z84bhkMgp
UNXVJbHiBcdPC+iwgnzEsdaQS8owp0hEqGUb0mX2gO4svhsf2mnR0PtGSJ0JL8Hg
8eqpOQwZAm5gh3nH4P5GlbS3C1u+lRNCJvi34P6Yi0QlSTBmh/98pQBI4yqkpelp
wabaC2dI9WnLpcjq0tBedE2zDXcOIRcivM9TuyM13lR2ipcp9Tm5Y03ipYqCSevS
uHwwSvE57hSF+pWQJveI7+xmwIKpzSFWUXsaOcXGMEAvTqh1tdVk4ufdfQ0KDUqI
owG6zdheylspXrtoA8zxGtjv3QlM3BLwXr+ElsiN7vAJgxIMlDSxFgyXBem/KjXg
r9MV8VR7hK8K+FmQrVdk1T4nJBtiw5wsbHxEtjM6y/VmUFAMWeFykQLZmnHuzCAn
wcu0dafW5XM3gRjDwxoQuJBeAWFEDx0vs6maiezYLqH9H2Fp5VTe2lulqN2OXkDI
vtUIdiN6jLvS23zQoM1MFdxSrFBT7A+EXOEmbKHCb0IuyGCLI6Vfm57fRzkTVUL7
T+k3m7oeuGZ2MDR3B5v5GG+dDQh6AEreZZ5HT+/OHDINs+B9j3zAG+fWjRc+AJey
gVZMSbLxITukPR9OtwXNbMYPEu7YGvx08K+x2l3Vi5l81imk7ipQZWilMhTLkFf/
KKN9Cw3IQezeGDhhOISEyAjcayccTA/MLsm7y14wYjdszk85oVIiO14X1FcdbSYz
fX6HP1hXAyMBu8fH+qvpdOi5OQO8QkMyoUOnNh7df3M4rA5X3kjt81A85SMK3PzZ
Gx75hEzBm7vieWn1n5fPYl4wFMcrF6qEZeHvgsFt60t2R+MPMEHba8mtuKzZHfFQ
gFoZ/wtvFqgI1fmWi9HUeqHZs6KN4gGzTZ+TiApsy1T+85r76M8KA03FR4BNbbyQ
aWPQy+vOecCgwL6i3rY+l1xtWzyhGQReX2WXvVDXMDDrEx3bhpn7AP9hTHFxzccA
Od0/etai8tCwaVXsJAWE/IDN99YY5lMk0TUnp3fjdakll1cCNLafDR2lg1eHYoqW
z3geXNEBz+prXHCDZVY3+E3UsObpInpat5dlq7ooM39WhlgG7lkh1RbT4y4Yd8Hp
tfgI3ZW6CFyixZXtRyFJ9Fo5F5HKLgQLPf/CZ/ezFyc1tRQ1PmO0CNiZNVT5TiNv
4PMEq9Pup8/EMaIVr4CbeyuRv3HnOkuNTZfVSMST1466b/kLE0r5cDdJNaG5lf88
W367d2vGU9arQxtvWL4AhtCWrtIFgT62xPH+N/5QnwMTdhNFZI9o3jUJLBPnhvKu
uCtBZTWLznZAQUos0aDUsW9dsBqvnJnO9d1srsd1bMV7usdnDHZm5VAFKg4kVFQx
4lexCvy4SsH6sW2jsQkmpIfBn1lXvPK8V81MSCd6B7pecffWXkJQ+Q/tCEvv5QYU
YHcp+ul5bPtmee0fnn3+sA3CbOMN219RTAX4cC8WzIMBUsLVaOoHKDCyVzdpaYm8
RNR2BkZvZkx50ALN3Ttstrrjlk0TuKl9pWaMd5ny3Swti8zH2abmQsGT1+6hJNbH
LqtXYILMn11KV8PKgDrIyN+nDPss68eJAiTq6eL3xTfbjKro7ukZO1pZiu7Z0X9z
eQwLEtMIkmncfvBiUy9FetRYOqjAg3NluRSOM8iIBgSTU5smmungSssYGL7/NJHf
Pd3SecEu9btZxStJT5WJwsBkhws5RWBD2z2WkmG1Ei/D6xLEYXMiui7V6dLZq+yL
XiOqsTsYUKgcurMts3r7r1VLGpGQhX0nct1PUJYGYb3Y6u/J0tQ1u3MwUJDUtfcc
c3w+FgQZaGx47SF3kxktjP1ekrJdzL3P78xz6vYMkP0fR32EljQ8rvs5qkPKoRrW
CAR5XntSniJwadtqwKLGjXlr9xO+of2lo9F47blUP1n8nzxc48ZwntaO3sU9Zc5n
WFfbXxFlCDKw1MoEiuNBKMZK+7rqoq5OxAKaVUfCGTtgT4lHFeP5d0WlUetpn2kv
z4vCOWeU6r4I2WTdlS0MUOFdbNZb6zLXnBnTSPnRAY2XU18h6pmaG3Z4Dn4+3FDG
FtRbc6rmRuJHSrWK0PeOSY3/CV28Hj/gLo4OHjpLyYBJCPFVWADKc2UJl6gSZvY6
VylHVknAeiIdpTIfWXRb+KH93Oea/fC5sG7K2744WG2BINn2kE3Gy4LU/t060w4W
R6Us/G48wguN9NVLzFT7k2/FTmamnlcnbPcVgnP72PGMg/NgukaDbrdCpGu7Mk34
G7qduZ3EJODFbpQIskIlMyxhrE5iufM+ZnP6as4pD2+F6CLixoRpfCS7nSz58Ux0
nrelKYW6dpptyB3YuuviCZB2gDV6ekN5FThFw3ckJnIfY0C4wRhVigjjPnfZcSS5
vEisGq1wPCfJewuJRpzTL72ulTafZoKxYDwPWMzvAIK8Q3yL7RpHb0Gxo41O0zp9
MM+fPGT1YeBPVGxHqplZ0YQH4kcEUUWNsSAv3oMejPLf95C/l6CRa7rSeGq8HP22
f2BoBCcsedY4qlvG2ZiqxtKwDffI7y2QIpGyc7doITqf6DFN2ifXB+ZM8mt4H0lQ
vCQtk87PvTsGuCoTfTq5Dr65eb9n+pU8TTqkTKtQuGqEHBirtwQtZ1QbhItGy7wf
Akh4qG1/h/ThjDGzYTlkMs/66ilCeQrvwtVmZd42/ruXfdLK4cyIGz/D/kqYwJic
vWlmYlHmimduQ9rkTdl2WyhJe1JXDigQRVGoi/GOX+01eDwLiBtHI30UFSZrndHa
oytuxcodFq7jq/uEJbP3s75Ht/n1oJFO7C8Rbgvw/DrlCy1SYv8Gqvnerf002W9B
xW353C9Lh5bqPHil59THmtFD8Ekw06QLMN9stCm2pIQvjO0SdpW85x/LUv5V0TrE
FJ67aNXYqj3TTEmrmJsiyDyRCIMw0T8F+qO9mZFLUphzFIfGHHFav5VB+C146iaF
oO263RrVAiIm1RCsF+Whm8G9x1vYuJ6KOgakcyc9Es/3AbJzXCKEv1G4+cSnGul4
e6cDxd0JmPfE0Q0ttb1qxPqSEYVijXVr87kBsIn+AgPMIzOB6foQ5ouxZpz10jyW
+NZsKnmt3n0YeQrzGnl/dDVdAPyuO5Z6e+xN18GUQeSbNM7yKfeZ7iCSYEKxJ7Iq
rQGbvqrw6sLeEvb6KMIEb79WbUTVz0CfceiTkEYCjdsVfltCJ2YObGkTzURsUeud
nj/bJPCc5iNp84p2RjJ8UjzD4mYF2eNaCQcVLBC/1G2+7UUQ3sxlLNHq8+4jUcsN
m5sjfzArKSqk40suass4zrFHH7hmTlcFf4T/ufarSla3Ta1fpNhH8JSIqnJv/mLO
wTUZ8BJPh9rJwKr2NZ2NwGHOY1BVmr2lT1jbmh3YwJqWnomfLc5jHo05GFjN5DXd
HTWTFSs1i7Gef/wg/4NxxrvXx18E5qO2Yp2ykDiR9CpFORSJKKRI7H4tHVpj3OsY
b6utPOIGH/s9igjKrcaOblMJ79mfyACRcuhyZAufrAem24r/H+z08Iw4knUkGof3
ShDX8LmxqgVMGlVclGx0Z5Xy7YA5NfwG9C0P5xenSeidHDjHNIympnlrqF+W8K7R
JlhxTUfvXXk7l/MJpHxHYq8NkLnnqTVWnN/XWkOoHw5mc0tq4KT4Ll4hrgVqjZAS
DYqtmB4cRhbSEnFdKLu0sno+oI8lfGho01VMJQf9i83YFRyOHKT0vDRdP5ZP9kDq
Ls58Zxj3DLsnGuVILYqcGDGUvxUVK5qvWyuWLBjMYzDFos9G+VQ1JtJvp9ALSLGq
5NxLUS80mkAZtJKhUKkax6ifunZ8QDCWL7AjXIUEO8+7l2nSM7DeEG5C3l/DTu2r
WeCY971maLOf3aufE3pSdseYFiD5CqjT7UElg24pAElTKadtOUMXJaCnCXVVZ9Xr
lfk8ipHWfVAh5ZZPEYW++qEkdeQrmUP51sZv+w3QVgabb02Xl052s9/ROwTo/zka
gJqmXy0fFEF8VtiGNE/8KmT0mcHchux9n8ary99Ms1zC9Ci0dNO2XLOUPpsARAc9
Fu/781VugXIszQvQPBP/dwPMLLxXGsU8JuYHkBoURltC0TsDxOXFeMBOafkOk+sr
1vqy3AED/Igey9UBt+rfjnQaICwH8rxz8Pt+/3yf3JUmjq99GjCZs3dL7DummPwK
kywnL5ILPj7F9IqxU2I8684vLAYzZtTBifg6Yjh78AY5CwEjJpqORllHtiSUAdaV
jHwOeI1yID4Z2uVF0TStHWRLQgEMx5acQr/H2xl7UKmS1RniZfIIa9YgglQpJz+w
itQuAVvQivkYf/uexiQjEsquDc2FvIf46WP2Tv7mo0H09pa5Ij6J66JNrK0HlQZ3
9p/UgqF4uk5p6s8sVMq5OvT3MjzmHN5BeWnunxmigMG+hJvswcQ4bycJoIt0fmW5
nl4NhT6rqsIOEgR4KYj3QIMNWxMdEytjNzJZkCnRKDzQ83odMA9gSyv4Z4QL4IAh
H+GP/WJygHAVojAqh7V4V5bnd74WsKEX3fxW9tBva/qqr82JFGoAj21+ILPvYIyT
WYYwkygV5XyfyDRcX5vdoyBHEKO1dkFMuZRaF5YVHH0vlLsmmi0WXzCTlkUrRPmP
3jPnSdXuUmkGpdtCx5BBzPTFCpGFuTZ3dang/9Lz+kEGfV/UdmaJU5qDs5/n/z4e
NmXDJX2PGdcl6Wg73Kru/zXHXENqcojq1M3PO2SDesAI9RkkE8VcM2koR/zvDOEf
q+bhUPU0hXE//5Hx3uVxHT5VGi8tjT8hYMCPmDjo92sq69eE/0+/eVky0nfywVy2
7tEnPNJSTIYWR0lpX2QmeYRi8rMFPGzeK5CyQ3CvtM9v0225IOjdEHR+nL/TbbDN
rBZypNY8GqlnG8CfOIyn6/ycTVkqElZI58K9NTKm7+Lmn2sx6JxXDXFJtVfkU377
DY0ijDFktjNMIvbmFSdqOkcq0zN1Da6OhqnFDg3P82yprnexmOGLdYsec3RBnH7a
8nhL7ylpeXPNzJ/zYDivz2eiupVysZrO+BBt0YfiBbDi5M0CxXgeRjE33CeR0NxU
cnC7aZPy3c6gOePWHMmmgp8eYRqcxa176rt6ZjtNz5WHXUiULPgmRTH+Cv1Isk1s
Fr1xeLVee7QkwYZwKTHMTkfQKKuYi69sgOceet4lX+oXIwHZs6uNoy0h0aPYsiI3
2Ax70WqRXxYiT9Vpw3nqLmpOFtx6BqsFYhJiBvH8gz9xL4wt7e8n3aTnoyCpsBUD
0XMKRkTTj3Ch1iE4jrhwwprma/4dTQllK/UTDtfVm1FMDRQIkwpj+urPYcapuDnb
njxO96OL9iP4aM1yJTqlaFEUYDs4LsTpqo2C1gWYChu8+z6NDib9OE7w5l4y3wVG
zmAk1Iiui9uUn3BIGhn5rD2oXFfhnW3BHWqaXyk+3+ywXaJO2Hq/Wp+NuDO+mYvo
/RlODMjXrlrNUTcJO+Z2DsDr8gjTPFwefor/FYL1aoO03jz0JAWUKk6ZE4RZ9yyh
8NwVT4ALEBmbm4S27hOJMhV/oN/aLAYPNnr1bfh02DqQ7AJCEcp+epJuqrqpf2kV
uqVISXnM5l7GDbhaKI18uZqczfbacDVbXOdhPba/24ph8bmuj01ebYUFA7Ewe8IV
IuD4nFBlEDQL4GrMucZFbBgaWcbpL+3xEQf+B8KErdPPm9gHNM0krkueNJG0pIrZ
fhQSf/N2OtcHkTUT3aCtLzwwVFDBVNTC0ryiGkr16r9HOZdMbHyYZKy1DsI7MTbL
1IfZqZVFwzEVtXWchwMzG864C9bp7wITpfN0hyEenXXYw3xsyrWdzwDwO1f5R7QW
TUHE4M0swoc4NG3vO5NN/9OG5ZtE03wTO+6RPM/QeQ6DWRmc2li9nBLTt1d2Wpr5
PjolsYInlgjns1BaYZXqGgfx8oj0+tNuprp/pymR8HRk02WVckiLgzjxttZ57D4d
FyKReIZNXkNXQ3m7JwmjLKLyGy+MP0cT+ooeCKaprQvebqHfik/afijv9MmNgPwh
zd3dhlY/fw6Ic0dYLcv5OTpgZ86wqyS2abSo0dz+i9H3IaR542BC7nJasFvy5A3l
C696KCsW4jvq0u/jJntcav93s+Y0yotzlja9arXR610OVHHDC1c82s9/E99IHZp7
lQkJSXK88HRnQ59UMBDM4Q+EeX7nvjcB2zZt3tjhvGOl4bllojcTAXsWSrLNOZGI
u+ksfgDBoOjalbAaPoXJ4yJ448IuIbwHU5b4TepDeaM1SXvB2xJDPppVVIvqVpGj
wFJeg55Y6BT6WMc+Qc2u3jFMlC/Ph78Tv3VnW9V0HnaopnJffiKRRTwcHiThb46N
PUpp94CHzKo66ZFJmcUg8AlgNFFJY8pY9CFXGbjEsdcXJRP5UYVXeC5M1DxbO6Wh
EJM5rqEgy78Iij90Kv8llPqK21bcSfi7/AsdvHriWQE9rlrqKLmTAcEACQcv54Du
eHdzyQnwmjtqLuFcZA8/W/RqeolS3CNs60lQTzOfIe84vcclwjLq4waNZqjqLewE
jao7EksM+GpIfZ+mxX7fTe7GATadqPiVfjaVuzepuMsKtkEXtbgGifPm0TtcAe8R
bgIBl73C+djkkmiBaGSvMbjzaap5nubJTvoS0BqUbHN2vwhsrByoWPMWnfyi5MTN
LJWB27XFX8K0RoBt/6iVMrBrErWbY16K3+E2+ByFN5pVFpCmSl5bCS6GrlubGi2K
hVMEcf2MwIAvxH3gqUmG3FRqbbfMt33kv/Ci/DjGG33ylMrGUBg51tfTIleq7fSU
5SHsEoFC8TBH/hnl5fGtaKkOnTNFo+XXxvklzpJpTUGER/8cOff+3o2mzQKzKceQ
8hMcLBhaQPQkDd6LG54KLTFsLvOVqcXYH7r5TxcoDbw5V5JHLIdD1CgsssdeDqFK
mapUTTa1S01aLn5elhH6+Evn3gJfohZG5GMT2LtwiY5Fdv199kZe6YYY5rqpygc9
XQaDjy5gaYn1RehSKVl/qEdmZBHxO2inOJWWBw/eU6zBtxYqVm6b/KhK+13Xsel+
ylLUB8kCzc3aL/bQQTusQ2/1SxNlT4hVnpN2QHJoY26IoXwI9CxISdgQ0PMtnzP2
p/rsK+O0AjlC9nlnmbLKbFb66SYG5PyyoYOTXnABXqszLXaJ0IIyDnmSPu3iQ5k6
q0GLlj7lE+Y00NE3A8R7n4Ca1U5IPTxtt7TQW/u6oucMeNaqJ8xTWNqoTwt+UCvx
hombKBIDDxbLrYS+tIYW/C42Fh+MB60VLdQXe5iIptRfUTuMD41WJKevPYy9otjo
eYUcFucHKpELxuJM26P8k7e6rH2kMbe4ssf5abma/ycljv4ySUsPtforG9kzNABv
KawjH6aydxO/l0q6FdtYg/mdtEiBIR0Q0Az7XYEB/d9Hy1V6yBS8td7n1Ic/OvO4
v8Eyz1/eTp3P85di2YgPFaO6bvuEnTrTV3fw8hNEwC2QuNMuGcJhUDfhpa8GtFcA
zv7VhHdO5W49qEspQIzu6p+pe1vp4Tm4KBp2z4qDsrzBPRGXpxA8FEBaHNUd9WNx
sPR6j67osPbLCWxNov7IdjY15Ivx8+eAik8EX2ySf/RYlFmvCeSXP5NS2CZK1rO8
jGa9TuwlL7zMwC5XnZkdPfa3QLG3RoBboZiCGLZ58SXK8i91cJ5OBMYXq+/7SBbG
bpPwYD6Jt0WuFDVgsx6AGjMQwPTz3RZqghAwA1hT9FcyumzIQLMrr/wnfEcrjOoi
NII5X2rW2hxJQ+IHus+MIWhp/BfdUIfs2YAB7fKKSyjt5f19snMtnq26IXK5jjF8
ogRssiMSmeDH/DdLs9+IRJIYoOqL9ZdWtwEnsaYTyEOLv0/wPpBNiVj7i2OkFAwv
P5XflHaCLt1JctHZI0Vgr01cTxQFVD29YP4VmL10vZQOw/1g3Y+xySMpii4o2ZvR
HaJYUQ5lG+wwdUOdmyDeW5MzNXRTy6LPZJorjvAp7T1LF/KYb/26VneXrvd9J5Hu
1Ja7I1/Y4xJ4ub7v7oz2A0nT8UcjZhSneepDNQOIamkUIA1GfJvXKLJlvKBakCow
AmFtF+He1IWRBblZdh2MI1SyC4Zx/8eZYrG7Gfdg8TobYcz2IJfb+DzJZANHMphe
1gaejsKUFffyihrO6TCLb5RFPacltn3hJIu7v5Ae57BFwQcooMP7q1QhBxt3McB3
cqX2mQ3P1BSofQ8JhiT/0j3oZX1IOBGV8BrSlgSp4HE0EtASSohiszaDBfAPxprg
RbiV2uzn3l77tXtVd3XS3UG+vPkJTAaRN3aLtLKcIJVhsmfCjFJE5KJHm/e8G/RI
Y0jN7Zps7D9A70vdxLW49Ls2FUwU4ofFHjnETAgmIIf4sHfo9KYlOZG9+W+qIwtB
f8IgoKTLHZ4G46qpTGb8PNun2UR6i8EDPLuSegbBDn8ldiO4HjFr0mFIkLiqo1TY
LaQfxltCEfKh3fKdprCc2Z4hb0SsaERFEpRWj98HkeHgG/eNarVnT3GBKGeB0MuZ
evq7JNlvJokAg7L9eb2i00XTrVyqY7resFbAV4MSoQkxaBpOFuw6NUldaIzAIucX
ST6J4x7Jqg+g8ubzGl2Nzj0hbE4Jcn984G3M8uRK96MFGMLEI7igOkeLU/dfJqqE
Kd+BxDTTfN/7noyzOw3UAahh1C8BTQoJxQp3TxVUZ6XQTuh+lfxrcnMWvOEDm4t9
mV3gSBTDoLut5Rj1uojEU0kYcYi492Ztn/7Yq2XZKzfjvN4GeYrG1RxhqYiFtYLI
jqFJAdnBtQYVuyfPrnHBjnRK0FjF/8/cpl3dNBO9Xn+cyrm/3AJsjeMlSh2xEM80
j03ikCZlKRfk0FaZNlRVGOcFtPb0GBQaS+NKpZzaOlMmmw6LdZi6uQvtL17SpUem
U6AWIZFgkhfIhWfaigOgv45cuAGoZIFrfmHaVDOwTfkdl8JXvq7vdylKtCwgIRcv
EoKY/Ym7SB1OftbSlZhGverhjW5O3lBvgD9No6MxP16KWWf6m5X/k411mHKMY3dF
Xtxt52slL29hJ+wwWJzeAE+XvK2cjIeqMOhTn+cl1SEiv5ic/TQNL4Whh9y0o1DK
ZISbBvZTx1h3bmwl1DTpLrcz2PzlFB7sOAzRy/W07BhtSxpDDzO5LxxO2Jr+e9bw
NW8uX+1VI/FhdTGrpL97Nhp0oFBxJoZPhR1Fs92t8PyuTc1bezyiTdTHSkAjeiFm
n0m28CnahxLw+he/yXCwyJS2JXKS+nCLOlfjmQYKcR127je1JNgQpujRtDOpm9Pg
ftE+aB/3t6INUjjuURRzulL7jdoLL+QHNMNDzepzcU4Dhag5Btc75M77115uApt1
qx534xxMxqzy39iK+QpG8h+xV8AajGo9ynAAMR/TPXBaSTMGnUOZqoXJU2GW3S/e
STeimOQZ+zeYOPOZSitBs2O7BkOOwNnoMAv+g+XMDgPHANd+AqnAFJTWghYAudW7
ugiudcZaK0pQTScp5oQ8L481qyBfv5hZngQlow18qntzX2L0V8c+DppjQQbrfxKx
ZlRRfzf/cILnUjJ5hQQQPUrZPLW7lvyMWUsCjghiFiIDd8TdHGn0tYy32fS5jllN
I80LtPGDo6DzYUF4WT+Zj5WLKRxwzcsl5eD2OPdWSmAbnMx7B+EXW030i7P7g1kc
FuBHSpJrRdJjUwsyrLu2OaJfQiNqmTAKsVdTjHDuK2R4ZFbS+wvyY0NZ8iNkbtAn
FkG4o7r2jzPSBMRWZsFzIBnAoFGFAkuJlyPYdGkJhQ+EmUBMfdrtEfI/lhbqqx82
DDWkCXubUwRkFtKREIKyuRSZIyh8xpr+uzVZBXxkCii7nkEqCUrRl6UYxiDU4Hcx
u9XtMRtAwBpyvzeAb/8+GBxDNhvFVEIN9KpcGdXEbCwlXk02t0faA4U5Mk7yEJbd
MfXua1mmSmG2x7QROwLzI0sI3da9Gt8apqNrG0dM3fQyvXjImOWFwlchU82q8kLY
aoJOcrNjhm4VwkSoJXvohACz9YuDbTh88kV6e3orxwS11x5h+e1dmpdmjVvO/uo3
YConq8UuSjU4HfauikH8+b9HsXPbkmHcYwI45x3+Q4fqhownAi8cogZW2z17XU2h
BqoCo/Op3qFLc8wnqU3NjaggkqnPUXtF0khD0wgtjFuKFl4alOqaO2x13NYnXt9R
OoCW60/w04UGXxQ/Ww/1S3EACo6PCkrpvnc05SEluiSZt1CP2XFaVTT01E3e94f1
QIdBdNsInSsMviPXEDOs6Ene/qJnAaIS6h+t50mUujOSi2fUqgRKVEEUJYTGb98p
IyY5jwpuvFPI0Tga80Q6KxoRYQ+QObysKwwrrjKp35sxGL8uDvq+P2htcNc1iIol
H3W2tvUCBnL3N2E79ASVZTIhDMGJC/gTl3X+B7Kli9tRNZV54NTV3WM7f9lNerzZ
WSd6GkluIty/ZqX++abUrNCuSB6e42+B5UozuDR952bfgGuJyQs1VWWPPkIz0f5t
Z+WpN0aBHdsESjQGEaA9zDZ2QVd+qv+Zt8WNZ8MYWv7WuPKhBofS0NKYfciwspWx
ae5ZrpEuA936VxAb4t1Qxn9nosL4a0UuVmlCkN3ukPCSiRlBu6t4GQijGW8Y1Gsq
dkj0saoXTBxWD6Q83XQFetahdDJ8IMhxaFomFOC3grYy5xBA6DHxKUgwC52mKlqD
xoHu72y7U25FB0s2Fy6ZJ72XNuNOy2DDNk+pMP6FbtUZoY8p/yRPuKXEmNNlAb29
KpJUEBJuONQMBD/eG5FlzqxS8QLOJJ8LayLm+GUNM+dvBPh/xLTEpgYjeU7NyVaN
XvaU5QSwljF0t7ZYDIQ7uV3wz8JSkZte5EQ2GJiDuMdWLKQqnU0l/iMehkY909cs
dOXmLfHgJWMEQLl6cZNHE1iHIawC10MMOh3G3T+mY9KIEYsWw2Qe8P5BP79ME3zI
5IJ8TpljetIA99wAw/gJFW4avvWA2rCT0OpXTRZ/skMXJDVg+0lVnYqAHEHZvxMc
uTQCWmlX+sq+yUPYfaNhImk3+cr2aXD5TmAZGDy2FPAQfsgMbE3vXC6HDMnTne7x
IFHYNaaR7Y0ioP1Lx/rxHkZw2NKtlYIeIoBwryhlEyqP8m/ZpB3qY/CFzHBQJPee
fTe0ovCtW/AtvSLNwmnLPZft/KCS/KjGsfpZ9IsJWlUn1SCRuVPKz3+r+Sh9MLye
SFMW2Ntt73lHirUlxwMKo6MwDS91vNfHibNCiGxofcOSK1hO32QYElZBkYmhhEtv
1So/eUG5f2BMH5+2ywWkW2cs14VYIsz1zTgQBwNiait1Sa8UCI8001rkFJDcfuVa
f1xs37fsWbGfANzT9TTBX3JS+tBBm0XFPRoocjWdl6Js2XcN2d8CGPvFfDgCc2AQ
DjqmarwJg3hhDpFHTec6oKlQRrWnmq1j3g4B5NDXmySNWi+jQ9cJFy11B39TC93Y
pFBkAPVRoyhviMYR7iRNqENl4iTyqCQSYYVU/G/TprwP5x8+DyNZW+YXeHPtJ/VF
KtjN4Qbi6KjSKODxSgOwWs2oSWUnuttZEMH5kd8wFJufCS/UU7gaurMSSkZAUr6W
RtjCz86mGryC9nCB/nvf4TkaLLT3wC+An73v+sIxOK2GJbLJ9iRWKHRLnFykrfjX
Z1W+KokDczqRdB5D3JYcug8OI/XOrRVy0n+hxknT8RTtiJw95wzmjNikf8VumpCz
6gQSI9DLUo1v9LJVbiBTlMMSZMr1sm8nrmsTZizqfqU5UOfimZEAGyr6s/VdiZcB
OcZB44jI2aHL0xM25lVRd/hTpJkz+APf2d3Geu6TfkrHyw714C4jIN1dgUBCNsPF
3qpDNR8UANf7aw2OmW5l+/PlBV8FdnSfNreEFLZuBHlkMqKHvzgnR7SiQTLiT1Hk
EEsF37AV5UdXlbcremyfk4YORaskSnzRnCUisgM5Hc70Fdom/lrbuTW2+rca2eHn
TZ5cSq7ybeWZeTpv0tEV69To6Rdd+p+1J5C2aJddNKUZzyARSZd4oZLCXtl1uEig
9m2hBbyfzyCLmggR7q5s2CgoPIXjgJF8kW5TQgtCoPFFtOroNX4B1OuHaGRHWrih
lEDdVdNJtvYuDosyx26eFnSZaLggWAeALg24MHJiXPVqyDJMCBlfvTIL4rl2dj6H
scjas1i9QJtUdd6rm2Hob+g2I3kmrwK8P+1xYlQCUWQsKgLp2MLWjjqrv/jLgvXE
Os409CChcaTRmwEY5rOvQM1UgfmSuwuGgKF+c9MoS/WDGwu8egFA8GigvGlsqSk3
EFuDddOxqHJCPCsjW4NIR8gcpe8I/7tMT3O1DOZ0gTIvLKdW1clbhv5CWP49gpjY
0rYk6b5A+eeCByH0Zd6a0DpfiGWAqAx/g40S4IpV0P1s5b0ZEEq886Gvc8o4HFC2
exUnOmZZhNdlUMmDgoKOeXUyb6KvC3+WPn/JpfnIBzTOZjWCpc2FMWZNE3m16TWP
Uj6ODxfOHDjio9mneuJxzXxGbVmCaKCkD2gMf4tq/ZysvRfVvv1zSsMLq1UooXXO
0PFDl3O0B3XBaZQM+FdPbWskvtVW6xVUEYJad99nkOCcU49JRCKFuGPJshHPsH/C
R9eInK1pjDinp85RrgQ2oF8PkaNTspXtq7YrWGyrs3c5c7IHDGiwSJO/GMIQpDF+
GrHsVZkQQYKagxOncvxWumo3H5NG4f41yWjzNps6Np89qhGT8067+FqDtKL18aUf
b23ewxbmelRy4pKO8XP7JdDH5RmJNTt2+VPk4krdl5/M9eUBxljxhQWG9h+iOE0Q
iDxtSDUbfsKh+EBllkob/T4Jg6+j5uIpKCpUYhS06mamOva8uCRtPDc73Y8eAkEl
orXylwDltIzLm4nh/yGUDGfx0o9+gSb2iaSUDp3P6z3ATyvALgJa3y8zYo9Nbv+7
GkASEk3GHYq5WhPHxsQ3eUHE0J+K/uBb5wZwZZVKBGSYTKR1+C3a9UM1LSZd0zRV
st9CeFQxIOsdou8Gtrink73mG1vv+O7o17aly/splhWApgUv6z3fKF3GUtCwNnPM
/cRHc4m3YsFltgj+voChQBitVCOm6ces4QYMp3hzYLG+qCiismzJuPaM+pk/GWSe
fqOKn4q6it9h6z0FBuHyi5E4Ce5hDJdJOF8SkGYvA75RjwD22FPeDq8gWLyJCy38
x9fhJSUrh8OZTBk0bzhDYpdczKdOrVAdMMtoouwS/122uX7dfaD5t0cr0RKprAQt
rvY3dhqwthOhF0h7xGqF/+POqQY94RX3ImMRgbwctvpiImV8dIFyMz/pLgmpE87r
3Hl9g1WoKqe1X0CRltexKzsIkVHWxkGqJ50YBXqaGi981NT1wolIqBmKGXQc1hEh
RjaRJyYtQEsU+lz2EtYndtMV5zWCnPNlv0L7mQFnRF4Wwu3XeqHxbeTaj6UFdOUZ
G0ONrOCN3yPtTcaUF5FxIwhcXnl9fSWPoNkxTU+tvsaVPaRoPFC0hejjSVc8mKmQ
gwkYFUsQbsXMcs1nMZFbNPP0m49ET5aEetf4UPO3mIrREOTpmnH/1gRmbAJ8HPiP
XSO/LDHSNUeMiNUSBxMbU6JtAOQ+TlQ1HRLs8vqFP9wWIpmH5B4I7486lkTM8jGM
dK0ld1DqLm9x3RX6dj0SWkc5fRoKqlgh0/J40SCbs27LBl74UjAMVeMVwiTGq/MZ
K6N6WoD547i4mq0NX5CElL6f8Zbao+wwMvvRY4vzh6WJbTGNf6LErTw0T9VmDPZM
7FnT0RtUiFlegunvESq94E381sh+fSDYCF+jUr8NYedzb+WYPq6Y+TpiSPhkyAoh
u5+FVsqMjyNaGRddO18YSBCb1+i091+nnK+McWGNteunVTjpExQDfNxYR0mg8k2p
C6xh7+ZQNFg14F5Q8TxekaDsD6WfzUgolqN6aL+tt5X4xbgiKwifeWJ/kpuf2xp7
maQu/CjCjW/A6+B3IMFd3Aqq++nlRcH0sSNeCyh/T+w3FZtIaxFdhHTAFCB44/4X
fONsh5q+7Bpcsny6c/x/rZ2nvOXdvpfgkqTtwNMPVF0aeRD5IkmiQrvwnXdLSEUO
/kCxU0cHtipIttINAgOFfj1qjnVRy7msai9pXwfPi54EQRLmyZeiwTgxkGejsOxo
Dh/6bQbQwaeKuIEkGDOgi4ytrSswQPW+hu1ZOWL06PwNxzKkDSf8gBzt+aDz3fOd
9RAJzrySQ+GMdfa3BqkoS4vFUK1EJo+3nab8sSZ7I78sRLcMOcV49SNGb7VocqEk
r0jnuWT6TFo/EAf60mGjJrYkNj6tk+sF0s/0woAPNTnXk4YSELMkgMKGlaKPBPjW
Niubq9rDlx0cNtmWu4ZpmnxrRI7alca5BhB4R1FWsPygUAsArND1ZrzlPhEUWurQ
Mp1/t7VMZ1rSBZ7k75mp69IIq5KXLh3NuVMIEPoCQryDQ7GX2lIfi06yPxLfM7ct
swu/pJ9iHN7jxjN1Uv1WROrqYSp36+qHtJkt0zVLnMYIIPx7ugdgdk+wlXoVf039
CtnodLXVGY2o1XgKIT2A9dU+PXIU2BwHnZf1OZEGBcBi6Z7XFw7pAl5VLZRcKeUo
tBcrA75sfud8t/qEDybsGHZPvOYq7KocJ0IPrmhHpX9MdxPx5q6m2aWkPSXx1wMw
VYHTZ1kHycPSzqUn4sMCvoFSfrHePzhl/p9686TQByREjh0Q7CwBxAoGTMcRWpt5
ARO3PijKyielgSmNoH2f5qGqG8QkFFjN+sjIxgYB+zlABJMY8P5v0nlp0P/3UEhT
O0QNaFjOibfWaGCg9NvBHTR4WngLepLxmwN/tkd447674ZA2NNQKP+VpiQv/bImX
z1Su4qKMnDTbR8n3j4haUOUy8xSpdYGkN236NDYGT/1uKw+x7YDh0nqXp/lW1GD9
UPxjnrRjsBojdBsG+b465bi0jvP+bhuGehRWBVU7csdsfMOt21HyARF8wB1ce2zz
h2VldPqOrATrEz1wvIQXi8XRqok+pS+nsTd40roHwMsSSF4PoBBX1ReXRXTiZAB7
hAZhnEYbMta8J9G6Liwy9lz9Mwxhu1OxhXa3a/na+jY4TPKT8USl9zQnhMJ17U1a
7s915VK5N/FQj0XazkJ73BffIoHaUe+hJ7RtgrBxjEwYBQnONAbpHA+MFAmVr5TU
do3O0Em4IGeu158TeSVwXPElelEk1SVpUmSESyfD8wKW23ABaQ7IOm4p+7Uiwab7
r/cx2Qv4npyg53EjL/mVXj4/A3zIFUUeB4ITscPg2yUXdjijpc4KifvoKkZmoUar
hniBTuR+pOfpFbvxduf1j9aXnEptrb2vVxyGTc8CSWngi/jn4t3ZAd9wrqz/knfv
SEztzmw4qzNrBtO386rmk9J0qvyl1Hv2v39OWRrHELDwmxoXOYl0McbBFyEY1i9C
rZw/I5aclM8ItkwRjnJu0LEZzC1jemhBO7fBbH2PI19EHi/pWw0WQHZhZ+X5u9D5
0ZxEPX06qwrckf9vChKdkMgLWo3WdQI19QIYcn7kH8k9je5+m5uLjDzbkkxieiFC
HZ9GfJDXQAYEBU/XZh+VRAS7ivwmcT51Jy0VxVdtBTdDRAoei0yvDNY5u78evVVf
GaHC9KoraOBI/2RuthZQk1OazSVo/4LJrDwZm8V7WSKKB9YbfZ9nIslmeL+JNbB/
NookNXHE4Xw3GCXOqtWBuHRe3iHn5NVx7PTm3a1P0OJhhZmc+zK2Hc35azH1T3tw
Va052pf8XCnBfqXiAVBRUu+1ydDW7yFHNV9IxvA514DTAxuPFQJh3+Zr0Yt3ctao
AQIkItZruJlX3fPIfD0VuVybJGF380L0Lo392Y8GyrUfr/v/4LOXRVvRrLLOyUGc
WC3mp27Mq2zcv/8HJfcRZJanjc+0hH4HP7gbET/PnTolORTA/s6265f/PUPAWabA
Ww650rJzWvS+1UjTOcysjQzlkHNDtpE4zz91Ey60g+Mcnuq1t4IkAAxLbA5s3TNU
rvWVSfVIgwPyTyk0lV/15AP3tL7WnSXRK79XVAf/HHLHOejunKvG4TJnHLx3pUAt
cbQlUW0OHBe6HjxkweHn2ROyL2K9IuNoFb6VYMVH3XQsgKg7dSBctQuPeTkfBti5
6WD1JTdggWYo5hYKBq547dn6hHy+eW/rJEHYmLbLcvQZBkoMFX3mnVc37ln9FAW4
qVv5JQoyZ+47zNWnP8AwlNx13tqWGcKbuTyLijjFjQzsvCPQvxiqj/h3jRRZJq88
9QyjOBmcThppUStOtHEhVp5pO1QGaMXfrKJfcbunb0nvNNImAzEBK8NnTEGfTMn6
7VpxksuZfJAnh2W3ej8q8eoM3pV3wkPb8uB13w6A+sofdttg8zZAAwguV+hcmEgk
wwXS9P8MtMNSI+8lc3+kLrrN3vrln57CniOYLtV50p0DXtKIWwURn4Q+FndYEQk/
4QEnvO27DGFEBgeerciiHMwkf9MTn5w+HIQv9zl9zLyhNBqeYaZU8WpYHdvg7oYM
C/SyyQRq/idgjm0pXl4B6ChLkJTx524Tv5k0uytp5m+Yd6X+WUVj89ufJgdq50FD
Bta7xFRFXlqlecqGK4N9uqg5cmUUkj3+UJC8lfXFjMeDFS3B49YnoR2a6+D9w7uS
EkOmThubGUDw3S2XsJmOwplIWUQ4Kncf9PBPnZu40pNXRm/h7t0iX6gnh3F0Fh5m
Ci4+f9CrOte5007T0BjwY07kMQM7hMoh3Aa4ztlicUMGiLEiMK9LpewG7LPcZ5g+
TvLvfQUa6lOLrFztrWaR9c5+xevhWRTDuWBGyi6aFmAutdRMXXj0tzZBBHsqVjwG
1TgncgwFw9Vm8CUmUSaem7tYgGBCp3HY3fPMFSu4yaXNusHQ7asw4T4DQW7u6n00
U79ldz3c9A3niIvKL1x+IRjWiLE2MoEiPbZRHejUKQq/NIbucjPeVAjQP099sjN0
ZP8HSoDQ4KfLzYxvp0vpLS9/OY/ud46sLNQdWy/40eYkZtweZ4X+1/asgmIEXihX
xuIJa6tnpcRXLGudkoJpE28bDph2fijdiHYPfjKDI62MJZNcXdfd9pmQQdlnQZJG
93W0we7cpwbhXHEIXBevCTOuQdvOmnxUpam58ayXugFJzpre4BfPEyqafACLGVvF
xXq+Tjcm/Zemr0YwBCdtA5vehPes8irucgYSXuM5rOaZNtQvqZKgINUYCUW7h6HD
zAKpv5RYZyY9uK7baPAhR4ht5HtbKi5aExgpX7qQQ/TcR/BDMEwhRFl0bFiAKC1W
zjtygr0EnlUf05vZCYV1zu/NeE9G278ukSE6GkhMPI3jQAx1+XLsEC7qZm1y6JVj
VQ2OS8AzcgHK2NSUE3Et27iFGxxPU5IuGBG9TqoOzH+Gt3KdY9rWxbr6i5eM3mYI
32dVsg1sRSMBTMSkoI/8SFHJkuXfRtJZrj0hiGFYsDP7Yk+jnuMxh6GQ5VEEBUzN
MmPeGqCX0ecmmgsNBuUKStpcSAWmPJxHk3BcMBjzuV8tEE9f6bITMJXY5ZuhXFMR
cnPlvz1tK5GHE9IgL0HikqcCrzBrqDPOzr2mrfXAiSFVBrDzcYLa5rANBV6fT+L/
mjoPB2wtyTa/jZsWiHY2f/jhlX+YMm7afs7Wng5hHfAJNmkAijrDy8Cuj5STp6Dh
LpmhzG3FFyP3EEeF9prt9Qs9rJNqNBUphwF6eapsM1FBCZ3iDuaT0wrDgibAiiv0
e4j3uFwpVwmSvXUoAsz2FuXQnaSVgM/xaubv1xpvuquzL/li2cpMMdevgOILY1Oa
sMT5VLOtZDI2pC2G9TZ3gnteW08YzC7wMqENQgEIQJr7W7KpkbJShs3auZ/KbPaO
EiLn9HceiBtlya3RXt3xt7mFGqqHd92Dfywru2xGmLfg7JcR4wOhZ0eOxArh/e4Z
8WPCBNqTk7YlIW+QZPiiRYBXgJ1xOeg+n5H1OiO4Bc/8eFqcIxqO+gHs/uN1ZrfZ
OmCgXawHZ2OJxvjTTzpGpZoAHO+owYnSd8o8xHx9v4Mpu4efCfNMKVVgLL2giKKb
HcBu96mQd6HJIfEx74xDVu3eryTsfukZz8bk+0Aqj43lseLZsRehdMDTcpbVywMP
OfeJbWhYDfRnOhe3cx51AsC/7z993zM6WZvHsTr63fkehZl6wgpGhXyvKUaRrXk7
PTYaJ8fEIM/FQCuEZbvM27Axl2sEBVHAh3ziKk7fUbvm2rm9Usym7u6l2exdpN+b
hwn1MgoCiH07LLX2xYQBMWf6bJuyFQAS1tR2rxXap5jQRE2quGmIwFWWHasRUzyq
aG9CxXo3eKYkJbhwYYA6+OLN4FYW9+eIxqAb+Gvcr7AHWkOnFtoKXRMpyBr8FrAb
as3IzCHq/3ZIFfRTgsfKdDKMX6SmHAtyg6wzTLdC7XeMeEcZF1r8z9wFbgnVH4/m
M2/Xex4tdmXbHGYKb6JFVyZjuCFn/UTuhHjyhKaCHW7d7jdhOBiguCcNP6fzMLMf
zPXwcpPH5zEnMJaFZrnUFQAtosz6G2VSEuRAd4TO96Po9IfHwwLpHA7085x4lH4a
f5/dKwdOFjZycxJa7wAnnIQpsOOaKA+oVVUIkJeBsq4Zd8a142Tpm+ACFyRKssvD
IhTPQhARf/JnEseZWTa8+Q8BIb0qE07hI3VIVSJlUxCCTM4TIceQw8T6Baamjcx6
aBkbygL7agBfwvNXiapsIIRRQ9yjldyApJxUe6rsf/SGRJmQ0YyQWZ6THx0cczaM
YryLVea9hswpC2wNO395aLsR7ilajfDqLBKO92p96bl/bJg5iXxrKpb5441XI0J6
XE5Y7V1CF6c56hLzc1Q48gkVMotLQWWog8R+xxTNliQG10CSuA7hHnzlEF0U+ASx
/zy0NlXiuRhYjQKbo3l4+2+S3/lARFucMqCgakKDLeJCSQX9hA6c2PF17XPFBfAp
LqxZfl59o+dRa5aLhA+AYogeDXI3agQxP6VidaB1O0a8dXPmD24DjnQiJoT7z4D8
kf6jIsok8x7pKGkLtixMCXdV59+6Mfc+Og7oFO6JE1sFxvXUMMzJOekPOia2GnRg
rXR6Mk6AUXvAu4kDlDdOIgzFpweYlRxN5GyiDzhQ1qmjXv2tvx3mFmKdk0hJf0rj
QtSEiKCm8epIUzafgPT7CaPkH/CXzd240PZ8WsvK/REXNrW2iqxs5XeealLoi2Cn
VFzJ5feP3RmgApy+Z+k9sSmoCW015I1rnJe2YT3olzNxBI+Bey1lvznjnrDTkl8D
vYQPaSmCQg/XRbBX2PPu8BHbeZ9kPEGDBNiLkRxKp6x4/VNNwFk6RJvEHBkJx2ab
Dw0rVpgiRQiSis8z2TDW9OZ1ib/1HvOOfGSy1X2ZiwRYbriXw0GnNrJEzVirgS+T
5GUs/83iZtFIGVO0Ocp8IPbfqW2a/PY/kvLWRoNPs826wHhZx+HZd2R0SDOffQ/Z
OxOi6JHeEP1zGEzBdxkO7UEhZN4uAbqx+24TlB71dVQOd8oZ4sfMsd0i6hcIed47
jrngZ3jVUhwe+01MLAbWNXDc4YTbf0rtZr1rRVhq+kvnNVsd0oO82yLxUJ5lu49F
44Z2ntzdMTzP2ds3NyUtd6+SUZbtyS6k989PJRmaFyjvdANzK1lkRx+5ukv+a2q9
CUjg2ugL7mkjf1UaYA2kEsMe1zgQCXzHJ6CoXgakxgZzbh0fYgO7wUD/qanJPOPE
QFl5M9+NszmbG+NNIuWXMfj1UnlUz0cmuH9U594T+TSlUYY9nTfw63IwySBtmxnT
LfsValA4Q+Cq9BdHnmMPy90LvqHdad5vX5hxBlLZTUP0D+LvVQqzIxpqRi/UbT92
u8YAzyvyRdzy6J87UUCpuK/da3MxfJ5jbmRteXuGzymOA6tE3ibiKfuF/v9dMqU9
twldIpHI7S52sBQQWGhHImAsRVuA8evjwek/NuAjGpuXF0vASCHJKgr/HzHO6xIV
Rr+UAikua+TA+MwZhp60YXU7madqdgCgrpbnh5P49i8R5jMMWcGarN8OtckEv6BJ
A8mwKTVC7CP9WqNtBMaTKAitIf1wf3e7JxlriiVNE+ZiRvqf9zGkMGTdDvso5tHd
PckH6wHSIAuip0qT55PWsYbp0h7+xUBsKvrbTop5R17Tj+YxMJcbzjc0B4CGzCJW
qy9bqsbLJ5WVqGri6ZoMY6Iusrs7ZN6CFLpkNNDr5wlQ0KuVS80HK4GZR377uRHt
k+ehACg84VylKdlBynO4hvTIbI3wy1z9TiLuXYEjPae3jWtUBdeiA5GH+KebcHGR
XEIYzP331ZFWv+jz3fVk/iPA47PpLb9HrazzSLn24XedCGzvSrq/xEa9oSkOOFG+
2l6pHUWKcRsWuvznkMAnBIlNGv7sKunJFnartOlhe16nQEVnG9cQEdXWxwYyoHi2
CCwzDx48K92YSHWdUaoEmwE06wZiQGKj1IR4jR0hi2hnlJRc5FTRxCbTdA4PTyoE
nFGbIGQVRsYIFsqZdJJccdy3QCRKcgxF7Oo3tZhEex6K6LegcT44F5WKXN9zzWTx
ggMWcmGdp54a2gPFtWIlr+T8yoEZJnbyQdX8MTEqlFZcjD1x5xQC8T2pttJbn7u1
TXtk7G3+7TWl47XZstHuecrnRLb4DUdEBmM0mn4VtYhAhmRmAQSjJEGEBOklxtL/
I1L+GmJCz6813pdl6eR4I1Begtm4KNdnPwDrA4QEIz/V2MbBYlPev7W3dFpyUzia
L23SyoAyG4RzT7tJsFTuAG1xlgEO2uMoD7u49EH9XC1YYTtefMBMH9cMr0ni5cpz
fR64pXwhORTR0A3PAuqoGDs2K6YHGLuY5SiCYpVu09AFfNbXAP7aIiX9WPXrxKOg
5yxG9GUdM/kgb80NT0YkVu/oA6CZQeL8yPHt+lM3Lqh1ua277CrZtQxg7vuIXHY4
Zmac0J9lTSFR0GxYmOajK9pdaKIz03cssMkqOKuCQmfx/KY3YJ4PE/+70q2qgb2i
K5PmkFjmxq1iRplgjmQNPUH3DyjzegJMmVQ38WWKueOvYxAuw8x9qQPXBLrIdvaX
agMizxqEI3Ukj//DegRZapeyJtSMARdgFuQSORPE72+MmtSZQHA6JtfJfyDYawIv
tIgGvwEbp9ebQ5o+505X+4IkdhNzJluboOMZYXTUN2ZR/hSUSuDF6WY+mtwD+cFn
8nglBAQYH2+lAGitbtHKfRT8kYtCqMq0F6rb9g/SLOk7hAzCJ4rDhJFWcHIvWqmB
mhJ4n2HvFsjsIHt3k8cusbyIxD4H9vP0qpRUCywcEzmDjRtGji91kMZHRvTSDhh9
xNYSje2oFMX9djZ0s5EmmB1QJ2yJaGEH7I8KYRFCqmSYVU4vwcRlZBDyFX2LxnqY
PTpGzqCbxmweOqHnhTS+QuAWpTrx+ST7Z3Q5YMPehwsqwQ8dcBvBfQ3v2JSFHDD3
Oezqg5RdZ1NM5Xh+RcDkms3KiHRzDgyZu38Zi8E2yCMgEgEBZN7qFyZ7J2nOO1Xy
/zE3sXA7uboWluFFewyM7s5Uwr1XbOVtHzpI9zqV1ZC/0ZMCCb9YRjbAk+ILyNtE
bH7J6T5cwGZ6AB4WIYG8ofaZo5+3wwmaCYk5SxF+cgMnh2C60ci47N8q0MJnvrLj
i/vLP+mhY+nxGuJSnRrsu4f90CeSf/pQ9uxHqxNdVd3SP1pluqtdvGmx8m4cItGn
9Zdk7kUoQZnYsTUmSvnsBAzkSJSku2WQWSR1St1t4Skjtx48GmEFS35mZmrP2lSV
r0zyn9ycy+q735azTZA1iQ5znArOxeEuD9y/gD/EqnNTgLfG8RaALaUoGM2q79oz
RS0xTQTcG2iXOn5vApFBIX3wzK70IvcFJE9a6XQy0OO8fhcagcfu5cp/nb0BMVg4
VxlbB1fexU1OdlkmY+QWBMUTynznwq+7ak8qAUL6QS2BZEOPH8mnCe9sVm9Ft8FG
Fq5wFUMG4/yT3eMoaUtvpMFvfEWi0Veygx+6Pl9ZjmGxg+rMY/ivKnYwxY83lgof
QsDBylOj+NL3E/pfdhiT9nGeBNaYVZFUipJ8RUmuGQ1Bemy03+zym+7ZXFi1uS0y
NKPtxcAlVOqnLb5g4BC7voHIJcwNj50ZMLWyiuF6d9groVl6bgebTKmE1jCBN0wt
A/KFBPc30jICi6a+pA7xR/FASBrxsFG7F3q6hcM+LFF79+mUNEn4F2h8KuIQJCI8
AfHxNTKePiS9tKpKraKnjY/4nMGEV/xSwVRIQw/dA/avsJ3LwxPLgpPeAN1dKE7C
J2VPw+vG8/cnn7h04Fi2tZgte9hlEHNUlrYsTCEwVs+p9gSYOcgDI1utnusGM7YQ
NInudBlh8ymqQOrosaFQkbU5sNcActQWh9v6DBbGjWN3nlXNTRbCij+i66SO6Ii2
LWvBrALGCMJCUi9Q0Ok540xEQE5LE7tjzDnlQX+ukMB6ao1IKcwv2ip/wHn3Bojx
7TECVbSm7M/fNubvNApk9iszIhfKfiRaDGlWHj06MmPRVOzxWyMiqVwBu1dqQ8qe
x4WO+MMESOb4BThlq/D1WSi7gqrtJnBomBdwSxxWpDQXg26lX/+ohfl6VNXBbIMy
PPMAxnaPpfSKwgRkQr3tvqGo4ClhK2+8OVmDwkLfbI66TrPLb8Nh2FUYugq9JoKg
nJJc85Hp55khplvXztM/zJIWk7geNSdA056ik1OBUbJzespx00hS/Z2gDzEuOtIG
u59CQIUeCFtQHwq4wqyq0pyVbPIxUuv/vpVJ+nx1KTpQOd5ymktuIk1ArekcU9EV
S2PhsPICSpaDsaexXYD0bHBNcwTi94nrTi5h1cQNR3iVqColHmUBLLDKtXgp3S8p
DRXDlF65bNNUHQOAAuSXFQLP5zL9aGc3FCiRDVbToXfTY3XxzsKek7Y8ZGgl7b3G
mavpL0fKfQ54hUfbKxHfsxcgEiLAJGW5WTrJlJo3UDY2wReiP7Zcw3nBNJLYJmmZ
eiKUdEdQrW27FF+Ikh1+fH0dp5O7zq3LsCd/QBGUDcu1Fp5cjZ+Fv4jgfuUCDFhx
F+a6ITWTSiOfDA7v7zOIxgum3npfyEemGHgB3LV4SSatctHacY0qaqcPzKxD7ZVm
McR4CQXmftWqEUtDGmPTt1Zix/bsFQRXtaamiUzZ0rxawWwkISQfgWceQBrkOqiO
ziy3b2Y2DJoyZ1pkD8W6mIJtxaF12TSkmJIjb9pvU/85GJCzLQh6P7OyMdBZ6X9n
kPBAsVX86/AjSNXbxx/OjsGyzB7/ihcBLwKLT1LNS+lLCSeeDw1FkQZiCpPnB1Fa
GfVCUApOwSxNfagWDSwR8gOLy1y5k+3//mYhD8h0QhO0eB0kX9FTbCPnwqJ7XcOA
OOFaZcJ+wjMhW5xTCv3MMoCeprmMmN/3AIJ+Spy/Qt+sLu1BpNzlLUlVlVh7ph9d
F5Zt5egGX340iO8kl1/kMe6Hulhdd6q+5urHapGy0XpdrvXoVHnRvMAdnjVXtJsm
FL78t4SQitwyu9FLlVvnZ3ebf7pFUEQaI4CEMyQMRHvd6h067aDZ6oJ3VZKXxWD+
sSVtA22HmuPNaN5Dyg0FEvqx8O7I9bp61AgvOSRTUwN5qiCzpM0vBEKazmQ1Yjmt
kDZEUC4eKBscCgSVaaQDg07u75hyvU5X3rFPHxjw2+8O8u+tFi3AgrE9F6kFpi9O
5D5MORsZsfxKjWDCl7ENccjSrPDWWGh+zfAPRuU250hg0LsvoP1u4ZYs6hTlATiA
zsp0WTkQpX0GLpNpqpheB4+bkkX+AltZ8EkHR2lvoKIvCWtM2wh4f/KeYDz/npNy
+VpnE/upRTDYjt7Tiqj8YoP6nEMCZSBh3deAze+nWJv2M9ILaPmtLmEEtkZvtpRh
ZAK/r71faxo57huAWmjzfhWRJIL9kkkS7oJGbhPWu/LsaWdvJJCL8iTXaTuWxXJ2
osfeBsuWdbe9u8yWHs5FB9xLrLkPK41g4MJ9G+fS2hwCpsmNJySJoFYH2rIfwwcH
CIWgNwLGWoncHPq90My96DB4lg4DG6NHqTH5mJPUwFgB7p3RVKpIX2owD2RyxGdI
ee60YLBJGhi4vIwYu+/8WWAQ6Q0YSPtf+atii4lROyz18YKnEyUXdhf6H4qgh8BC
OMk8scIkFWQ1C6Ck6OjHUubD/0XiGjhhNNQjmo5fMWsVIjSBQqbyFdy/06qVIEmP
jHT2LVyQHKucOSSkfX5ZqRAR2U8fotlZ1O9nZ/cX6SuwCyvuhhhyJtniu2Ivjgkj
vJlMZ9LKzHF7/K3OCC2frjpLKgk7vyrgRh2WFV4NAum5iKd8X7eSRo5wynIYIZje
N7NAV340HXTueUnBEonwYi9MZo8DZT9ReXx7c0bFi+L9UFR+Ql8Wy241Lizv3md0
dWWAhWJr9qwJBfaKqvMIpNgRvJwevcvdP9IWZKiG5S2NZX/sABhMgPzppQ5HoB+8
7kH5LRmKLmnrgIB0J1izxyUxtKL823oGuT8CS/EVwu0n6j3yIn+sP0wEMvDDt67b
wLN2fDuILmy6VkngJ1ZdunRQ616XqaEBoy6tJ60wN8CW4q9Oaz+60Ih7iDdpwbSd
V7Je6QNVzHv61Td6NlkGwj/7JcHyb3tm79vhGZh4lqc3RyXFxofJDJz5zf56CVri
hBZV4x5TIk5cczmCMrS9nhuzg2MXM0fJs3h5YEBMy1YQ1EHBSZk6apGcpjWQ7NHV
A2B16bkgTCgmodBrdkckPlqL+XgVlD+gUjI+SjKQ1evjboTqRHr7qyE0uktLE066
1Rs2JkeDj3oX34yTa+cutN7QfZibP7RGWNWrzCPkD1eL88sllhPQSUP5AxLkTTaI
vACD3IS8Xr9YcKxre/OeGN2OOzyRu0U4hRd4oxz955unM1BbomdWx4O5vtQ6sDLv
csVbUhYntRObIb6dWmOeuPkkaTevkUiVyAFQhCyHkbIk91rVkVUtkN+r2r1DFjaJ
sJzxhyza6WqOvfX7DPNg0oR3RgcC33W/A9MMk5BsZaMmckgY0J3RA5zXtVrFxfHY
TLxafT7d7X05dIfTyPxEtgClWRh8lnuD5fs8YAfjpeLd+CwStcX2mFHNph6dJlpf
QOqGIOZEDZA2ptbRJFHPWPz7uuf7Ns0rR47JAVO5n+oZai0O3h6Lz7DW8Z7h6FLW
MWneHFX+UTuNpV1uF9v1EIsIWbQVyPHzalozaZfXgrqP66S5yvX3WGHPNJ0nIAdz
pfc5IC3ZAE63kFsapzCYyIA/jZD+WM2EK4+w/qaehYQMpwfzZjua2cKXqoPQxQFG
GIY2/0H9Qb6lSqKDlcTx6kJCWYGYG3LRNZCBHgwgkf0NdzXWCexA9eR4gE0nteNh
1CFPjMjw718f8uDf3c6jee4t4uByoEmVzhCxVpk9Al9+uI81cXCrIqZMoKwhR7Gj
U/HOfa2CnvxeK6h1kofH3YBYaijnpF40TaZjoRxqN4/3+rm1fbIezfbHA5SxYmg6
XQcG6SVhdqAU79ccSUwP24UlSLUnOrbq7RRAU7YutPYWYv0TPevPcnukZrkYeHXt
dZQlDaa0ygYdhMtmst/asiT0TEPZeMZ/B6k0qwTZeh6k82PXf8/4QnWw6ShIDMLL
x0CGLsoijreaLvtg33JOALitxNRp5H5VwoHiOfLDWc8AqpqvBTiKq45Q6yc2d8pi
jGPPN3OjSRSQyiLYe/22+SQ7hCxR6khSknaq1/QDWp4j19/SweJc1daBwph5B+eD
mJ8UfWS0yoEGbf66MYnrONZViGLZS6grSxqQ6MEGV3SQaOPQ0Vlln3mmK52Wy1+k
j5O0N2pEGaU1r/mPKoJLZC0eTfBVWy/zo3TXQra8cePAdRbUhOqv8eUQEqbBSrDO
a4lMGce2kH0KspKQxtXZFUhvKihVWY+xaTdmYPTgZzi5pEji0yQ11AqZBBeTuQ9x
5vi3r9YUll2IVeKzJAPjgoXtgNG0p4BMvihXlTdvip0C8DKJkPzx3lDDh5yxjEOe
N/JfZQcioeSYWxFjSCu2gWwpnCvKJto4+Yj/4EtC0/zTVP8gZHlHpfIiN3C7Ok8m
6KUx4gx1PR+lPQgxUg1F3PGg9iK/89NgeQ+RgjVRrCY8ud7UAsz9crYt3wFNIakc
Nw8HyUO7Lgh1VIW1YxH0fP1pDTXrDkMXOgMLG2610PblV2gb1GuRNQtm7mMcRTyI
1gWK1keGus4G1WZTxI9Xb0SSUT3qom7MI6NI79kG0NU+xW7A3dDfWmYjPZnRHket
7uCeAz70dfwsGSpIAd6Dp26bjSfBV/BtYrKxLHxm1R5t/TWXXdaSDKAZTOzKhoZP
PM7JjD2Ji1Rx1wADFU50HK/dHm9I69+mc6p8iUV1Nrwxgcyze5hbT7q3L8J4I89f
FTK9UGJrtVY5Boysq89gismFFqNq7u8UlhvjtQWHvDUaFhGLNafTKwPLTFfFkFmM
P1Ng6Ax4XSCoy6bNdxuyDIXY5UKIN8YngIBFaGIEcMQzXkvguxhXpbuoaQuLPR0j
6PLUPRr4FLePXQ5f8A7nFhQ0zZwp1coLEDbvdJg8b7pof2xcLnqtx3Zr+L3d3NSC
x4R3FPcrc6++J8HM/aVKrY6jinOutOSfOTrdwESFVyiHhTOhs9u1JqDJPmcQvrX1
dOwIfdrdine6UOc8dx+nQ3JxiH5vuOHBXOTPkSvZigXaFeq/J7Zlza3dwZxS6MUi
QE4vlA2Fb28M5vJGuq2BPxAcK+w27ZFDZEt3SMoCflNM+YMJ2pMbKUSnpZlsf37A
ai2eptQIVhE4sHAAbGzlaAurUQXcUdWExWIvehiJLTM8Wdkd7j07KXen6c/4mxUA
4YLm6lfJHg+bCJuXeOzLR/0+eZ/YhkoJu9eHiCroqlGRuOgF2z9cdgKCewlV2Ld3
UVq0eq+pMuJ2qidhbWBW8xDjZM4VcGMn/8VScWXOo/3bYVxkHdDexY6fn5FebxXJ
DD/aoUySKiwyAkZAIgF/y3UCg3dyThUXOAQpAA9rL5PXz0HGDtn5HMKoyEK/ce0U
knUFMek8SclV7x8aHEfSQ7mUH2+aQaZsrqPQJ2WqcZz3T48FLEUNpvwDyY61AyjI
UT3FNYAvF/pZ/lGxMTWtZwWuZNMwQHFPP3Qfi1gldEoMgfs6afoMOE84Qeql5Lao
KyTHlU0aYY4n0tcL+V9cYosQlwgtuUT2BudkZkzs/Ha/kqSNbW80+tnhIH40Ynoy
mK1Om5yqM56rhMpm7mnxzK0ZnKlQeQNaP5psOW4+31NSx6DgyxD05KmamXcprHdX
ikS8CZV420kuhc2zO7Zx+dJUAduf1p5nJ1wYFp2SWXDycdDS71sdznVDmDAtO1zj
iXyntN/KCtyhlrDam717/OD2iaeyt9OKkEgl/O8u4IGQ2lIBNZvj1BJ9HFtBfg9x
IIBZcsWX/ajukqMbhnZQqol00pIi5g9WXsjwjSX9kNtDZyIihIsmyA++8gg8R/wx
uc0eef150kCCCLfDayaODXeCuEtWLJWDJkLm+8BRIYvEWLYdoEfqDqGhAkRcbg7o
1TobIMn71nUNAJ+WriP2Wm9ruGDimY5CwbL/XTXUzMXmTFPULqLxiSB/pNP5HuHq
Mq3nmgGGdcat9vp+edZ7fwbzIgDh3Mq6sktSGOushlv/DE0M/iYMBoM1O6dM+tAv
uuCcaxHD/s2cjK3yH6oOBWyS+QOdO1C1IBct9sYUpRxVC496Y63AQQEzAViUigXH
+5mRhaPyrdvuPVKVdFEmJ75y4g02o8HY9K7iVgHXXBePA6XgkZlY9BDZmb83Ad/j
SdQbnUzsvHu8u2Nvge+oLdDlXtIQnkwGMlkF/5DT6CVHyb4La3EsAUoV1kzJYchn
UaucVU8BSUxBc7uDqsdFSBmH1v8bSLLsF0QyGC8L4siw7Jfl4v/7yaEKBGjmPxNG
MTGIHJqLZmR8Z5Klze3XfEViqMgSh24tWEychpoFh88uCexMVVc4Vv6/8c0A4AnF
qjyXYwf36xHVDV479FT5buBWEOUrLNw9b1UfFeMQP8RhRBFMpzVP/qJW/2Pr9Tf8
s15Q53spDKNoaou4ZqmUlL/DD09za6d9eaYuF89XkSydVIg4z4N5CDngMzzCiOg4
Hyb1CKV7xAEblvP9F51wxdGjg9AOYg1wBWFDWFmqWUYwcFd4szrMgzGBZyWY73kk
eGB7WMamQzIJiUzkrZjog54wIVJVk/oUsiFUDmL5NQziLe0zZ6ZrTO84QM/K9zbL
HtwrW0LhQaNIHbTYRKTSFJ76pLf+Hq186eUrOnfhWi4KQs+86aSmLSHpq3HWq9Gs
piPRP7lv6DliPuQGVGBMwi+x5+9YXVpLWl4BZO3UWUxA0VmBJRyDeGrgMeZCrnNF
tZ6oanE6rS5x9Nri5LLaaucDODvuzjqMPBhpQDTfAul8EH4j1RnaCLzx83RYPYiW
eluUlUKeIdoF4CfC3ov3uIOVtcCerD/0N+7O2MO2SxnmqRdZYvYEu3ra9Nghc8pi
vxyuLOnUs/H4bCiQhiJyJZeh4e4QB5UZZ2p1jomCq++pjxb+Khp3ZsAaRfTakNd8
omqTHB39GH2vk8Six3RS6OHOI+ofUM439CjXkqoz+fZX7igwhZuAQ4w5qWNaIdEg
qZP7Ge37tPnnUcNg+/ZUZhy31r7NcMDvOH3xhQYP+EMlMhT0o3PPQUQCjmxd4aVu
tvKER9lREH2O6+1SeI/HOZT1DjHKc2Bjdu5qhasAc/41Sru+uuAjcKNl8Zu3VWPU
hNIp9eOGomtEXshn/tfsLTtNVQo8ipDzO3fATwcbCCVWGvZ8d3zdrz97BBSLiEWS
p9xHE/YUAne5glXCq4yX8sip4xqRJMqzd+2yMZQ5yjCV/quouclLbmrJCcLk0Y8g
2Nhm1g3O/I2SJMw8LUSHE5RlQvYg79/WHaHuhDnY1hDt9IWKc+uwNG02zGBef84A
inv3fevl3s8ut76rAOnAO2nWh93ZeY9iOtR6Upg1ldLLfuUG1yaGjxdAl6lIvvo6
hGT48J9564v4T/F/X4cLlqWGoeqLvpefjlY7jMJTFVxF25D8qJnHw/z91HTf375d
0Llf0hc4OTBSKL4mfh+IY95cqiIRpoMzKwilLLRu4oHC0MzqdghT6cLbSAJ1keTs
dbndQo2vPPnJi2r6OIDbx4ZE8N4kWKIMKm5q6yAlU6CwSfYMEN4Ux10mDDb7ShsD
Hy19iOjZL4EALC3LJuUBTDWlfDBe7bH0EZ5RRi5XghujcGqTQexgw9+KgMzDR8mw
ikNQMWG0BUnx2/42RzKQD/FMKHVmGA4rr8m8IV+G3efGuc/qUd8ww2PE8yusqw9g
0wOjPGvS05A8e4xJBzqw1iAnoKOTxUw7o57XRhZJ3uKXI/oXTNBjaa9AKhnzj0uZ
Moezm+hotEzi/0pnLusqmyOKheIT1K1V6OrFxqRybfhWWY5QduheIwcXPdmY19Ft
OsDqN22tocuHnhn5blb4tDFR2W7vdziER1GbTrRQVDS3VBL71XdnVb5ZSOEzsI9B
axnT2pZEEhBN8TZoKfkQQwjBgVRhwc+TgXijPPCiqh9YU2KHrgUeV99c1PY3BPyq
10/Zjsd6BGe2Bh/Th6zFcCFjoaIN1jgo0XMFmb1jxN/LTILCdk9NwvvEyzHaeLpf
oCma1I3z9/FhgKl/BzZ3FrjOmwYI9Gaccf5whnXYKVdchf0Q3ZfY1x1034oL1P6z
u5r0FUkAZLLxR5d1O1du28QVcz2Iizi74wz5zjm6lJwcwihEQun32aZdoZ4jzdMs
LKe90PAgXmxlJoTZuVoZd2m44MXQgj7sQ/oDR8BlrBdXClsOJx5nxJRYCeZW16+V
IO7y7CtDve0FsP1edXaJaG5sy4jluSI8tPiAdeqo5ekP8dZ6rB/E6c9LF1FcOTnm
lWW1QXJxGCQTFl0RzXYKcTatpQ0URAGANnErwtAZfN+7vMQKjcu+IBZTT48V8qF+
BAfYFrPpJvo8gWwrbx9OeV82wW5VlBBno/zqtAWnCKlJ+absMwBCueSAXNqQussR
GZ1X/0na/CMmv9Nk82X1RXs5Y8DajAlUKGsOyO9S+vdiofgSASlOEFCtUCcAgZ18
SKMKCRiBPrgMBiMxxDwcedMaZzgu4jbnAE8ogw98xTo6jcL3lUTso2HpYPPavg7c
3UFcXBTP0atIeNYJAFYE6GtTuFrBF08xZpcTXIhUTYD+GXt7sUS6VxqbDgAHqcDk
YmQHVIHlreZewalzUf7m4XPsXjX/1TVk/QCnPrrZbU0iYYBp3cG8Y/u7kWVCUBXo
a9m6vx1JPlnRwx4G+QHjHspQgvlQDZz6ZgAesJlX1Y8EBMKq4WUsfAHPZhNtoVqe
ZFlRBBPPPe7NzwHyjYhvdQ7x4iYyfFSyOtZv+Z1h9pkzAcXV7LS599IX/46eT0PX
ZUNE0nW4GrpyzimAzVONqNpgfSETCF4tzON6gc2Ezidw8zaIQWNOo8WKl3AzNh3M
NgCoBq5z+Lz7eawXnEJ69l3YxvjL4zbOcSh1HCtsAZdmI+r+gqAwIZ4tlWqqfJWs
gLPumJMrVj+819fC2tRWBWgehd0GA3kHQ+umqd9u5UldFNyTucRst85k26xTa8HM
538TicNFX8B+hyRh0KLZxbvFYoXCNNMVZ4bMWO3RQM3K4PsdJyvppeX+d7NwGIMX
p8Uhe8ttqF/DtcWiEZ5l0/921WUlQJ1k7QjrmHOJzVL1zSyqQuV3xI+7wG5Jabvi
8puX/GqqtHLwb1/q2eEewsIaFjzxrfSpIUeRu2mJym/JsIPH1BYbvJ17Oi2k47Yi
kSfoGYAbO2KPBIfssFst4y7Ne94WO6+iSCQmhp3LKSuHGLr3moJLNbPjVBZA9HkJ
MhoqftSzZUkE0/XUVHyh9Xi6Ao+dCioGb8oxNmCmg+PV5TOwXoErzvjcsm88J6EI
7Sf0kr4n2VLtcS+cxZZfc0Y5qTF/xpqUItVEqz0AIkF9Js3O93Ea3DiwTTv427Qi
5c9MqL1fMoaRygIb4F6Y4NvT+PGac8YsHIrYDK7bxuQWo3RL0Fw7wP+jc7lQs/4A
sIy8wdBKddt8hgTKWuQ8xJwYuukCK41jr7mDpOQ/QFc/JfmuvC+2U9Sp2ugYpNMQ
UlcsuW2q66zQBG+BzGhcvelxyaem56zX2+abokukU7O5n2NXm1xG/ldB6bXnq9Ke
j+cc9s63/bheUN3E5ShpBFbvHO2das4nlXQ8/dTtfRd/1oNKWHDKVuYLNd4a3kgd
rhD8QdqZ9yb/kDzTkD4+1YrmwnivPr/91KtGbxxaBCBuOj46wyHgWJ5CBfTzBXCf
OZ7fIuMECLHPDMdOKHJVoLNpWqNxIcAS/l3Y52hqFqic5dwEJsXjYQvirPGvC96O
A8Gv6l6I7oaCQPk+1yTAnaBW29mp0Ho1hFeMuYg6XoXmNMteThibdPkGppjvldOV
Jz9bwfcgbmawGPvVtHdEGwWOTZqaYsCQnx6Klx+RPQ3t6c0lRg0+82FNj3o80MVu
BRA6W2IFQgftXTmEPAH8CU/sd2v7I1KixX15XkWn2wRZaIcoc62I0wfO7LxQyUuP
zAKEwWWV42DoRMbgi4EJkq9tApGGCjcvYwX5UYwDOkhpatTkE24YTrtu4KeGXDpl
cNkB6Z5mxovzEb7skBEx4eBMTyx8sQfCdvOaGRdJ2QR4RMQTknjiNQ61HetkZIHe
ePuRzfQXDf/ImZKLyWu89lhzDRVjl4so5WOOwGqwYJGGP++oJ+Y3KCJp9/EXAzLA
cd2rWQ6oNpZDhpc4KTc/Yktkh7qh/HGsMYdOTbl3wo8bALyyMn9cckFjJUgWd/Xn
GaanC4oSaj1dj0GjkRgky5s+F9sxTHZNx89der/SXL9Y4weGtfoWDZOLPdwMjKvQ
HEuZyNPM0FBD75Oli79nSJciCJfeHraVWAvoWJkMPBSOOJFPLP/PVQS3QfnD+L3y
TKh074oVhbgaeVNbWf+e8FmsCEmHeZVQ9xe4BT5Z6w2Uaxf0FG96qfTbobtdXIlQ
NVqTOJbOt8Mdag7FfIAGyKi/K3fWXA+ylCpmjpgRM1aTkpS5QtUMvImyTxRE4gkV
+Sb0KF4REKm8lPliWKzCPfSoCLCfBx7/TAe4eTpb2p3jRNUW+luLFeAJgIjGK7jx
QiQC/ylhVHSIvxIK0uM4su2slv1kHpMwAJFLbvXyNbYW6R2D9757cCgU0hG4vIZG
w7VEKRjIf5x0l1xber7bYFM82r7F5RcORdMND5avxbDjG4m873nLgj7NyF2Z6saK
cTxtZl03QZX5zc3vMXKEhRQEI5S24pVNnhy//e25BMk3wGi3C5YpXt4ZfSQNoNNS
mCCL2gq5Kr0KvCjruM9RhTjyBuMsKnW87EX5ciVgheqvPe+cdC9csZGHgSQ6eCZx
IXWdJEUOlTfuomIYwtT89PhtdarG/osEERCiFmpGlTjkKmdQsgH1vMMQzk4H1aVl
DlzMiH9QnvyrI3RTtw/yt5Qejt2qzAf7bdo8LOXydYUQhf8nuBC8cwqLB6kijnwW
82paTl/QbrLqU6fafNoQMYAiG3yPIl4LzOtDWtIDeGL0F3ZLefcg0VRldp/GiswL
lwqcywwpU5uBCl5CxnZk4GTlfT0EpwSkDnaEjBP3R6KM/0P6yFtRPNXxWNaUG9qY
TdTU+MT7dqql4cmILgQn79KlPHdyEouYFps5gSyo9puWDQsvc0GkjckjkH87V++z
3tLvNYFyseMbsoXKA/WnU5IEt+2n4ULaz5tbIekd1jans//GCm7GtnCcU4P+loyV
att9fWUfxmST0YZRzQUhPkYbbAUsN7/i7E+NUmd1OFxYvLiHVIBXLDP/qt0xVcjY
OOD39R+EDrzYYo59352Z6Eo4dLnojNqP3UChDJWTBdZO5C3myYgDWFX0o/ihxkxL
ckOFdwS8DBtfRo7DQfsWXhhM5iZRgIwhqSkdoHrXlcyJWcyClrfVNI8Ql0+pUM0R
AZGwNdO5RuSV+RIrF1BqHRTb5p0zG920FvvIV00ELsGyJQ1DrkXqV7zNO/uWalf7
2wuuQQZ4GJs9OMlA8hZdYvVAbOg62MYeGqu0FiHS8/x1mK8iM62SvExUPD03XU2B
f+RuBWAG8O7Ip88AyxGIuiwIX/OC+GuUgEZirCa/I/bHaM+Kw4CjlN2SchMkL29f
+hr3Sy4fn1mPuAPj5z6FAfmbdgPH1/6UQflYESvY1v8qF1oUEbOyVk/Et1LrqBH7
YtYKqHSgGOCLAS+LGeQE1Qz88q1W4o0j4v7Hl/4L/R1y4hvuij8lYYUL8H4jkmqj
exvkxAPw+fPzLUK+ivDg9wPljmRUSfMkeGEfHWrUgLiL67fOZiBhbIDDN0k758+g
zv9FJHp0J9xKw+jQ+3y5yNma+9ahk/1qi4iWdCWDrxWesVyDavg/7ZCWDI7NI4+k
XwwOcJ8I9nKm2MDojIsidEUcI2hfnoaoMIvdv8qRJce3HnwWSuMGMuo1N8e3h8sE
vhqWLD85TokVjiFJV1R9+ilZizVAMZ90+guRy2PRlAa7ZR3C+7znRYsucxceSb+N
0yuSyYCrkq7fwIaHWaZUQ1RCwwchKYjA6MD0s7Zef0D8ApaVvspe1BYRtiCP1oKb
+Id/iFaRlnbE6wtWyX7iLQ2j9aO69WsnRnDVwXPjRIjbU9gWKoiY/C0vufHTWABY
QumtvmcB6q115sqQZ69Q/ldDKd9pixTaxcKpvduPgXB17swlE5CIONPdG2bfLN0Z
yiSw2BjK9zg9NVX6XLdRTVtpB02QzqrAczQBjuBYxQQSNFC4nyYlsDK7jVvunCh4
rpttlp47odP3e1+wuH2iNz9U67ikUv/WCb3lCK/+qoZ27/7Q/j+P+4LYPB47FjT1
PjVsu3xHqg3SqUb+PHfEdtaeGCWRD3T3qkRPuUib8HmvTA34N6GfD1Q56ensYDbJ
MkkqKJWDR9N5EmyKW+QcyOAT2A753GJ4dga95yhKj6GuWMPfL/viAgyC55+29+xD
AWfD5xH23bmEZJIPGq7DnvVmdZP93eXQytvTGQ9x4fhhRCrU9FjJQk60DX+c0OLY
Gb2NxRMi6Qb1muhDw313/3SzqmeBglMeqMTM5jMSyWYeibsdnNrpGQnPTH6Taqia
z3QuoJDgnqAVJM+6CXpdajjlq+vKoU4gfgP4AtB/Kq16CYhfO1cy5h3av0/YJlpe
GPR1opIoh4B89ZgFN9sFv1tcEtdWeXjThT1NT/Nj4zU92S7sS7dy9zHEJjJruGpY
UrfkFDur5Psklls/pc8b4SfWCVTT9IpnkcoUftiG8PW2eM0HzxtqTpY194nBqEv4
BFqgzeE0qBmk4wPQd3Nd8zYCyScn91gGDktcpA6y655OspvotOBEQbjuvjodq+qb
egclyMJjzqbQblWsj9Pt6Z2WvBbjjaLN/5dR+lhLkSChltRfp8vuvWs1AblamTiB
hWP++3Yk+cAYc+g23cKdyZ59RgBApWlWgREPPq+YX2h6TVtnCVAWZtFUVOawL5u1
SQe45L6X/m51hoXQRGcYizjK7EfpXcLG7f43IO2SMevH1S7Tgrg3m2cUvB5Au6iu
iUt+9dBkq1pza49bf1nWeXyvHVLIYK7itTHc8DG+FR2AqZdNaH8mR87mwx1d60py
tGStNvEZzVXD/usQDpvhAQOsT2jrkT6/lA2yLu0Ff3AplhSF2TJde6KAU5+JTJkc
dsUksWy/Q8r8vmDTJID1ThA5wFt+aMbn+r6/8vAM2Hc7QdTvzXrOSuS0d7Jrts3K
XiE0bqoE6KyUTPOmjpH3uxhTa6Iitb9najEj4ecE0ppI9VRCzj6BdX5Nkun4x026
MGn99nexqk2oEM7LqhWYl+t+MmM4rIuvuBFlk5JRYrfmqrBClqDyccTFRWUPRP+S
Ln2bAg1FFfREd3BL74LkZxMqZx6zyxhswCKIWhck4W+hNtw5TcLhXnYcomoeNAvG
yt9CfH8EXwExGBrkh7MFXiAqrSdIScaAkLPzwNOGq9lmVFHaSlZmxtTo32l4iVTc
6lYDWS3QJYrw6E5bVnclXPtZukyELT40nGmEMA5UIeAPuo2dBJiFnTUyDkjMOwry
LekeWou+i23Mb2ZePMv3OM5h9gxyvcDwHmO6gnnrH1ZicLyW2avW+vRar2rrV3uZ
6VRUh2lzOw9tpJq1SdmlKc1JWOZTfQ04i+XVYP7FnbCAWtWzfy+LB/hwUpduHyia
OzwkVt2GQ31/RbOwDKO3F0lG++k69CzUM+Rx3V15HSAYQTRUyFxGNsylNWy848hT
P3HL9dHW/UkiEip/YN6/uABaVFCcI+uOJNrMjOr9rxfmu+Z0gOMHUNIwmRDxVCx7
bfYdtgbvCKRWy8dM2WcNQUe5s1PdzFJ7L8jn/iC1fB+21H9SgEEbCcWvqbvzv6Jb
+mzwNbbuIixB2OnEZSv5Nm3eJidEU3dC3PeDZSFmOnEuz/WxenGogweOPr4M/4N4
Pz/6uCFW8jzF8UOHeXxYeja9Z4nkyBCDLLobVw8i8um5CUWAitxIOFTg0/UpKIwb
FPWIyjV0u2uO2YH+GAngJiT2j4ql3nm9jA9USIMNix+GJEdo2Rl4OJdqCrk6bvtz
KJ40/c1OKk/rGXOUUMp7Blybcbrh75t91VcBsn1byV/5t6T9uGZ0w5ZjNtCXDaFv
SdLgJj3PQ/bcyn5yF1rHbsCTfqfYrwebfnC1CkrUKYEEb43EZfzqmgqfT3czYHNE
yXDk7H3nwvagbOSdnkhJrPYgC+VpBVFbJmV6z+6v0iJoihzU1PECIp/KtELtLk9g
d7Yz4FUmjcG+VNI/XYDtUFZmrId2ZJRXpfqknIkeMa3ipT9RYyH/pQRdKskUX05+
twbjKaT4BdmCXKuNiWoRBcqgKXkJb2Z9ZOEIYRJudB4peYWRmEG4OwUrE9HlMZvz
QsGCIkcIn+cSiNl/OKBYm4XlCRcvNIDjOQckAJmzCCPfp5nBrgqS1cxX5DbPDgAX
7GkP8zpzl33ZcQfefrgUE44vIgZTFOxFTA/GRmEUn4fn/cxWhek0FQl280jbu/nP
82vkNftCn/jhmBdQjwoDK4IRi7yyQpir1cC7ibQheK4jdfGaqrS6DsOY6hrwdgm2
SXmeifJVGDNgd5dqhxXzl1y5w908TlglwKTGq1Z71vAx00Zr9abh1Zxugz0iQr0G
CsS1deZbsVNwS4K0/KmzjT1YbBnbf3sDMJIu2s2Duw6qxP6dQ6BUcfcdcCJKqnP4
StqbDGxN111CRyailcyyS9RYOghQWe/UUKVgSIJdeMnwFrIO3lDqgtlz8GWtWco/
4zdVIvH/2XVFEcjYwY6vsB8xtCBqYH/hGLV4s0n317Nd9sYCWXe+md5PJoWlPnDB
t8BQbMtxLKR6JZBJ4GgZBR7u4oCRQUcSe1Mstxg1ERyoehsKljneXBSGTc6mFjAH
1OQsxrhI4IWgbpV24ALbgOxYw6OTwzTnxrAZEr44QWYM02IKb7Lvr6y5lTegL9+9
CYQIB1xyWfr3fIphs+3niOeVEtP+UuK0ZEYT9lZ+qw0HPVzIwqyoGUqBHrO6RogP
qHzLnXUrjw2+QfAl846ZomnKI4Sd3WaqHgb0pnLxTUHg7S6Oy+th6iDX4QKDLMmo
2E0cYWErPES40sBQ3on1ESDi7rmqrcTwoK3TbWx+5yLlFAaYoNYT6h6H7UMzsKPx
xq53CjE+Ad6sMdewuH6rsrdfwazBwWb5zn4dlqu13fMadGiV52Hl5z+F/Z+Am/3O
oSbXBW/Q12MKBLL8a3TZsemB30QpR5p8IvxnQgJ+5WDf4+Q4sB5uR0xkR05OLhtv
TewwKzhX+GtJ0j0hjBciSl1mPqiAIWmOfjs67V29IOI7LPiNmhnND5KV1ESkpIlD
cs7pQQJ+FIRGfthHryfsBVmX0aq5tA8NSV43YMDyDNU057glQ7W/IF7ilen9lh9X
oLjpa1DF79ST7y1LN5FmqSVTWmUaVF7gfFi2qKEbuzqPGjAA7yqWM1c7sVNViTJe
HRN+m3jyoBL9mXYIHABecbGNoNjDGoJfUUF9tbsPF+6hxDYobKn/SqxX+HFabWeg
m0HlOObbK+/DS6I54DBkJDuqu9MzhUWF4cz5bb9CM8HkXj4jYdyCmJYvb9HyyiKE
AlPWS3UtTHF2hVfOGq7MzznRyj+jqLg9+xpx4XjCcJf3Dh0ZBc7s0lxne2wQpY76
oCkv8MYPfoL0fbCBim7co9uihDLhdSwvZs4KXz4pfVHJsEkGxcgftEgui9NlPKLS
4c10pySBogEAJV6DypwUMbjMejPmsQNGB5MQHyvkQwTxbeaxLqKT7qSbCKR9pVFN
C775TitF+/PQbcdWIGldmAMj8ofupz1qaXla0atq4VSOj+e1sVnLmP76i5N4dzBj
NqqWbOb3bcdDPx5DsTRST8igEeQKAW2AuhfT1jHOJEumgpzJFUPuteF90iXvNbVS
eSVm7KtvFTweLv5WMzm5Iiz1bSN84/FGEtvM5S8ktseQm41M5V1Zo6C2dgK3Lxie
4HFHnnx9csoDlm4iS0/Md0un8YvCFx7HtStEi6UVmn1aV77+c41qYFfjrSl3Zlwd
njYaZ9XdTcVlvN2dVS8V9m2yFtkrvfJyBiEavuulPJrOMavdISYhQYLA3IvaEaHr
xXC4Uy9ug4Eif9yHI4F45fvs7LvFmRuy4cEmPtQpzcxh7DR64U/btRxozVSCUGPf
bdc7XcK0+orNrOrJqNsaqU+JABIPM9SzUu117ZZjxhPUhC/j8a1TRs6Ub/VRV0sR
hZiPgzgxdPgpdm0J8zhShJtFhpG5upheW3+YWeZDPwTq7amCojMJ+IZvPQvSf88d
IT5y+7y0Fbg1ZARVpTkPdgW7mI+W+DFR0O5wry187QxIOM+u3gg/scODeNlWGc/O
S3J3vd6lkeu+BI16rSE8wOSyn2yVWtr2VdPITvc7VLhx+CgeAjz1aXz9yea3OxiP
g0080j8qxaL1sjE2Kjp5QUvFDmbATGS0DgcnsXSH6wvMUs1zu/yf3JnLSomJNlZH
TusGNWxYVTwA6gP5uOjJGNnGlJ7uir2JtgdH3eN8F92+KSXAtWYwOPfZ0BH7e/9b
9os8QJpoCK3UiTXSzERbxlApXctTgVpaa1REim+/vU8jp9gtq7pJPoA2MP/GIFrW
9LlPCLjAl1b6BRpY9flqP1vMceoiloJY0EvG646itghcb6VTMqipl5XjVhb3MWB7
ulXvB+7W3jmKC4sWlqYI4dxnVa3tO9O0Rz3jhaCS22mwXMjFrsdSQ/kIztLzdbDE
YEdmoLgdlNG9/wVFQ4fhkrp+eTXLgcoa1GsYaIt4g5XKueOoEQarLsfYBuEMiWOr
RSwQJcthWPT8a9g7ojgp8GI+qbB+uKxLzrLA5oM4Q5PfbsfvLmKsERav6FnokSDd
68453KJmDDUq7d1omBi/1kRr38uuNl5xc84OKyQKDl1czvMCBQpEzzCK/Y4DO8on
tt/HIEoUmloIOI6wcVKfI6k+6AQYTUCAziExv7TOHtfwBRlzESSrYPaOML/J2QeD
A+qQ46rK5ZoSvJj1KTiFtYomoF8d9eHE+8PGMG7JmK9WYSL8s6DdtQPznrWxr+ET
M7naHUkxZF+XCqMBWcroJaJSasYQ1pDgcA81M90XUF6GhdauR/MeCdDQoTGCxdvf
gspCwgF4y/cvbTv5EQIX+ji7bC34tFQc4N+LFdKXUKJ05SNFrRgsYjeqnddJtzqc
zsuzfAXCyGe8Vy7XKo37CdrD0ituHVrR+WTkAjwkzd4XqPTeNm3zOblngBhq7VBA
qZx39/E9OC1buju/9eXOQasM3lHVW4WHuNRoDXgWu74fN23aRPe/B//RMAnWEk4E
3zuQNbDZCV+XH4BbihdmfOKGbslaoEgE0o8S7EKOdTsnbFbOpSBWpl3wKc2YZ+P3
6yZ3jYtQhFzNOk5fHj2qRD/XazEu7E3mzqC/fx2MOU5sN+H9vSB/OY/oVfpI8U8r
28vl5bHjVT2BJ2fGutVp00aLAktX9ImakfRH5jvJk/7bYoA9U4Rhr9m5LHNpR+iR
gP0UoQazg20+yVBtWYyvYmDRYWNpUafK4/IjoUx0yiyO+tFbLbk/4G4vqJsaauH3
w2sF3lvgIWWTJdaKxTHjilfB7Bk1QpdULZwRqip2UMBjyVvKeRpN8CC0nBoA8f5s
dLbA1cxqs0CbHPNthXVO4uvJD6G0LucplUopPsjbeZwQlJHCYI5+eMX2TMLj8r5n
1bMFQ4Kl/Sa4xmANWRNIfNTKPQ8On9Gq3DqFdzHCN0dpkWFGTNfqI4eHK0GuVZOu
tKK4wya7+SXeZNsdgOlrzbtNoXD0phU4KFf4iAFOdD6id5JK6+45EWf79FTsgyHQ
uJZeh84bctAo9l0dWUaS63bUJjl3z45QU+QWp30Hc+d8zmIByhr5MOqJZDfD0hEI
+IciSL0blQaa4nboMDvUgv/R12A8V/pu5XGyB6nm30il5LNRl+YNKI9L4eYylDKe
xN2HAZnEn0hSkqmhYXTqEhRSjiDgmL59kjaO3w8rWilQ98genM7S5VWyoSK7CutF
rCV+eZSGOdxtCXtpyyfVEh1gteCpImXtUbUlNSWibbGlFPdzv6bbQjHEvs77j2Uw
S+hsJvgKgMhD1QTuwp5mrWzKJJCizwQIxWzFSyw9bbHt5lwcbMG1hLBFOj925GM4
eIyf7eWcWvQSwezzCYh9byezmQyUWoPUbj5iYQkg9Lw1T69C/dNqTLnzH9zuLaX9
VeylONiV9tWQL1xxMEXUeNs4JcbLkBNdUPwGPBcRTOsTAWVnW33kAi8VzyU4n358
466KVQWpxfYATiCe6M2meHbTqjXZksPymw6nrwQehGVpFx0ZMhLZFqtGB2xkhrFq
fqspnSMEBDzI08BfG1xZ+x5G4/4CTaL7z6a37hOkM8sgz3n7Ha269u4xZXER1g19
LK6RIeaAaEmnDD+C3tDcDOnkzP/NpS01F0NU6WW1Ojz6k4rLvoaoBeQVeQHMGxS1
rDzZ/hC7ZxPAV5mQxbLc/fJE1VDIP+cznrKI8EaYI7milh4tc+s1O+MqCpsQ6kA5
HsPxX5LJHlyCWq0BaFGt+SdJ0hsYRsPDU/BRzrcn0x8OZzC7WGBHPk4IgHU3pcde
60efylOkOjrq+b0HMmie2ygx3s5uTl4o9pajLEC1+5ulyPQvQhOElOah8IX1TjWr
FLYbo+UT5je82AztkiYlU3m1PoV/mmZrqoZI9w/uVXUx0j7GJ/uoC3IH6c5OXy++
fBZy5pEL+bIgBu42+bVjA26cT6aVxPMtu/kWQXgnJ3JLSF9YmK5wiAO8vxb1AD7m
H/9AN0BjYV2d+KicxIMtAOcrKc2OakCQUT11+ivx+Vdm4UtwJ22nXgMjlwiwZcb2
SENnn5L31ExyKcs4yx1IUhS7ur3bETDaH4K2H+Nw7qJVwsZ2L7ajSHJtNzR2aAJj
TE44Q43MroQJr+XbKCq/U6LlQI5pte8OtpVQYLOLvGr/GyAGaoI+elZIfOebpATv
XTba5zUlyl90YQM92KgLfrhDYfJzbSLsvgUN/cQYRGmNqkvwBigcSoYhGlikX6VX
pfDXIZbeOTROqNF2GZYkRbmLVlSSoDccnRuxqejeziXOokgWfZdVW5miArS4MRrv
2k54Ckn2SECjIkmGTyb22chX7gJ4amjkStiHgdsnsQM=
`pragma protect end_protected
