// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
LQmCeJOF9P9WXsF4SiLX9bMgaytfvXdiwU5HQWa66hvlwFbuV/LbnKK3O1RGO0vS6Sj5VjhbdIm2
1rRow8u7zOQjZdUU/jHZGCA0jX8bUK2X49MjDP/SFAjO76JcSX3Ckz0egXQlJrvFfymzXy5uyAJs
QEyHhHbui+fJYW5FaE8dMPj1UulRzJq7jcpniSJbp8dt34xurA6/4zUEWEmpWQTM4EeEFz3flyJH
D76QQEpsC64n4KYvFId17PydU8sYATYgHou2SoLEGoVIHXyes1CedJSOP1Ckh/ckSfJz1WGFqXHc
Hfg9p6QdusEFcFmg8xuA2iyv+QnYNGU7u4uW3A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8640)
MzRXEbIFCPZb4W6cOs5CugOB6Bv10TQ1S3hCm7EONBvG96uaY0dxg/hHSShQrdoSQhaIdVBi9uKQ
A2POHVWr8ptkdA2f88av5glaIRC5IXB1cM3XiPhxkEgcFc+Taub5xpVwIgFidihYn8sm+RhRPzKc
PRysFZtXrBNFwr3xHkVDOYLPf8VVnEYkSuEbLK5vZksTekbhoFKTEYyk9xGso76XyfNcxwGe5grZ
FV9iCShS0mtP0pfnRtcT0AC+UEm34mOvGyCwoSV1lUqYqLxlWYrSM3fNKvj6RRiaC7bRDufxaZr0
l/xvdTZJQ+rYbYZioTVLH7fBoxGdAbbYmFEyjZnq0AIoPkCtzZ38jSosWFcebBDasq7cQ5eL66V6
4t0wpVc2DwROrvSUf1wageOzgkyIeh8qOVDiAAX1zqdzqblvXSMrk3Zc7ordH9L7sg+bknvxSSVM
NkCGwiTfoMUNeGtZcNNuOsh+ntEfiM2+5TmNw6AP/IHlB+OCHCoPY5tXhe8FAF82Z3woI3qvcblG
OBWqHxIUKYnibmv+7tsHfbJ7sm7eu8OjxgOaxxygt5N3R+P1UbQ6MhGQfda+qlzVP3iwzT2w9hnb
jvgxJTS2aORVbGFtIfl+txU5jH0fe7XzuaFqZfKBlXEtdnA3kUMJBFlrB0F7IspU+DRZhAg+O5h7
phUF1fc8qno+RiGNochnpkfBt21xV0y04f27PMhOOgEFp2t+Dr2M3jpqHleySyx6avykf0Lnfel2
JVTs+FgSsLeMZMcK1PmbQA47PYU8cBnc3Tcg1URN9nkFMdvJ4t+Tc9ITLY5D9/9Yjs007A1ru5tJ
qj6a2KA/U8uEUqQORmtf2/JnyVOn1nUntvtMaMPJBdnGiU83f4RP+2xSGM82gOZVfQ7CzFucr+cE
mYNiGLtoFm5Aaryd/fbRvfEEwwievAtAk1RPlSgKK1TribNQO0yMAxtHBF+vgFOpCAo47dyVUNwY
Koh/oIuizlR4nNar+iu4zsoFbXHj8tTS8yhUPoc7v8xlhxRHt0hlEYtjIYF6GrMtyINn8nMdVYGE
0L8QtZlCQZmqkRvXwOfkH9lkmJ6db+Wnwm90swymVTydf7zl9hhdpI2X9CXK9eePvghJSLBOI+CP
w9ddksSyW6tB26zygdvFB9THxbP0szTh52/gGCcXbzyBVPeSCailLO3SFPTqy7bZigJODJMweFYg
e+MBK1ZYMkVZF0VZrpEhOlid/i68OGgj1CHl/sUxPNouzbhSboGTYqzE9ROzI9ty5RHDaG2K+LrE
DRSKb3zYNPR1zfo6nWCs5DuUItYBlmRj3Vb2qsqqVx8TpxbbxIGaOIcqRSb1EfhBRsmdCGJkuDJP
BKSQQff7kmcBKPgF9DJr7ULEoSllmHxlckgweI0Ki6ZiPNDpyWPS/hIBf/+QgPYTmjHGS+GbMm+v
47dY9/fJkGJRTJlQ5SsGleoTMSfjMaJK4AeYMgl/j4F5a87TdsiHTnliEnIOl+Q5utzJ1y2Y9iil
BtW2Qgju7yQEGkY4cQezZ3kNRAf4TcgKcwq7Jh3YjIFOZD7n9mlBRrneR8FK73DFjxev5xN+T7P+
QBmmx9p6Ebt+L4l3FyXkzTYMqmVHaRKXN4n2BQwgJBRS4qcibApVILY8CYHt2+gCIjOwIrrC4zWt
0PjaDvR1D/Obwo9Ugx6e29NRL883ygsJRsztGNdhAD5levRqt2z7QAv1/Rr4M5S7qcgoQqn2gxI3
vEo1UEDeKWPrTZg31rR4olaKaLX/gwzL3DmVAa0gzHPqPDiyzqbkuWMICmPFpKLufX725PuqjDc8
JgkzdiIT/PYiWorDc+/qbr7LagTzeFKeDGsB0Bs07U4VjoqKYl1G9D/98Mz0loTRcn9h9azfuih/
YqodQN0qfEiVFlP6+4n/lgD9IYT+6zQNAq9/TQpXaJ92SYWigLxW1Cm69jr9CqFj+nPQ08QxmmWx
48E3Wt39Zj5AhKuJ67DbmwB2Rsd9biawRCaye0OeGAQbTA+ingiok8F91VxWDtQYzkcstzYEAOYA
ZN3ZpUGgL4xf8/WYawVh2uK1HplkN16r4GYfwePLIdN3a8Fw3l7G3mpoLFl/lSRPRS7fhQI4wtu1
neNvZpcrPY6LKBuIsLK+dTyVPbebmlQ4JmP8YvO1g+7NVKeH9++6sxKO+RsZUOjcTcJy7/7iX8r5
CNw27WMPtD8lYkmgZJ7lzIWG1XHt6se9i+KpJWofW9EnLuQlMBkAgfMuIhmV7bLbc0n3jD2dGqWs
w3TxuAwtecOsu7Oai1xbj+8bIyNlbP7HU7qcKB13Ng1JFzNzoewbHNy9nSS/jBU5s9ykATDTjlZa
Y4h/yRTmOrFNa/qlMxr/TuepKeYsnJz9Ou5Q6eZnAdWBpaBqfOXduz2JDknVQ8xQEIFoeKLr20JI
5JJSJ972VZpHcBB/Zh2BBSVZDbAOhoc3JAXGcuMECu0IYZlP1pRtVUIaGAdWflRVvFEzgyCK/kuz
uCnD4O1hrO8jgopSevdT1p8zIJ0tTGCpc1YXbYcTV0Nr5pVe9zldlMR8DtLrsb3XgQQUL39uR+D3
mdRJ2as5QV1Ji00s6+ql84ddEWoqnoDVOUbA+Hgo8t9NlAcMmCED0gsv+jHeOtOZMplrXxYs21fM
BKfeMfLfhtxeZDBm5+HC51vmIDElYuJ7b10nli13LqXi1SFKPyQxy20nN5d0fnVYJ08XXxlBxCoQ
8Qiio4tSW7PnFDeFyukBlt5yoNxhVOjCuLkD/Eit91I08rwGTuWYgEy5nVg0O78zDwp+Ktb0IMic
Bwwurqfr1CY3gCoAoAkf02SkYQ/+jIyS2U8ZPt7HopuxYx5lrkLYukaQDS2ngKzwnSNAWNGNRRD4
rsSByEN9dxDHChRxkV9LL6J9Iky4Z8iEqY3aG5MER2e3PcRfj9Ga1EMHthCgdr4xtInfoO0SBs8j
6e1ffAVE3qMCUL8jYIEGOaqCXE2FSuataYmKmZspRm6a14kVexC4dT88a+/x/wbDhqXqrzw8QkMF
zWrfzfOr46enAosoByvWnd8dtic6N4YU03sKR/j2ePxIuL5PGoqDfLTQSzmB4KvONH+fnCUfp/DG
HyhcG2kvNX8RhC+DuCwVNUznmZFcmSgeQK30IXz2VzpcjsuHKIJMTlBernSI3t6rjgAZrA4rPG4G
YBUnWqoXZOlpRrlf41Y6Rh+S45glzvFWuA7a0Ndsxm1LkugjhqlslFGuwtgseuITziVosS7G2SDj
ETUPeoKHnaOVcA8ndj6RrZarC7EmWTE3GKnyrk92aOmpGlCfv8LvUUZlft7Z7lsDW3tNJZWIH07+
sZ4ea9WjU2MPDLl5R2UcCMgn/bzliCAMEwhxXa3DomRKgtPV6FJr04v0RBJkjCQHJlYgI68Bc0Lp
att0Ya9zCeRHZ7JQi1pvnRCZcAO31VUTGBpgEsPeveN0udijOybv4S35uzE/RoEW6lcb3XKMQruH
bIqmeETUJSeNssT5Lg6pHan4TAQwFtphQTJWFW3U/pYDpJacQHsv5LNy9pnHWL8fSZ1rJwpWmkP3
OH+zVmqh+1DSiUxv5Zk075mgl+SkjPmHSRx65wPo3rOCOFlgJtp0Y41LX+02yaA5VwnGEWBVN4KM
bLUAlRAuPEsugWvWFGwzgeERAy4H9dkvNRAFSqfC4r7BelLhqMsat6Zvday4SfnEhqVzNUbKzMqo
wTkbwAe6VRbklwG12YlMkbrEbeAIy8YsZunvb7JQRX8onD86yIGei8FQalOoAPjbVMq38+W2PQoc
KWjDQx12bmb0OK8/QvSYsRDiX2VqB+AsPR2IKN4AUlnEkyK/6iz5QmGDKfpMjVaIbgDeQr+y2icK
+GkxyeBzUcHjz3Qz9je/QRuX+vktkI4MJajdJHqJhoVZDjv7cAl6+GZQ48sngwKBR16ikEvjUW0g
Ap2WCDF2FpJU8E0w9oW+CiJIBlMSz2mO1h2iLeG/HGAqhIyMRYbZScxZUm3wCXIlFgbSOCuWNFFN
L+VgJxqMPZIPTEyHoPPf9E48U3hQQGbcalZgJD36XU7bQRzoXmbajHiCneWj/lv89nkd9L9/I9Fe
5poTxPnBx7aBWbqSgB06y824WwD4eA2GgvUauOs0Tyc2lWIQ2EV+YzuLvDXoALg0iOM6WWyHGTfg
6GTccC3BS9I3myuo37/OR6kdpN48ASjSKtb39Ikp7HXpSAYp86Yc7uKjaDvcmPXJDRhykxAV9FdH
39TzQIKMTvZHTROL5XiMgm+h6AKa4EymNnBj8wKYaYkHPnWAeTBY8Y2pHBJoCU8+jNN/IuJXzPlw
RoWJSw6VYDXoM04rVvZ2gjqgM7THG7/Cq0YO1+S9P5RX10r7KflYRn9raW6OG+SRRuiYWhAuo2Zy
DbS82fF8rnBlAVTaoOSZGQ6OW8S8XPFRtI21iHmAu+0ZEWr5wqd0Lq12UKI+SjETnQQ+sCwdnb6D
hnUlAcId14Sm+8KVWXaMdbTAwH4K0bczvZOL02aXIX8EuJ4P9Gyf5I4YaZ6ImMQ2ILAoNNv1m6cU
p1rCh9veYAJI9xPslrwIT5VvoYwHbwLUcUQXWsicsVzxnGkaqaU511TqnkHVwILLjPpPw1MrSKhk
bbTck6SW+g+Sql3Ce+KlNPE5UT8cCuf+4PfBFOkrbaUPpxvR/G9txV/A+JWABS8S7Jj8U0F4N5bn
xBHSau+8j+ZPu0E0MTleL7uzRvT+SaocqlDOOnB9khl4PGVZB0d4Rz0TaSGFLHMhcRgXA1wNkLQ5
gvWmFeMe9LbVFjIlt8tEdKfm7RwMkCzF7/go+fxL8V2OS2aEzSKlUNOtq0TjcODxhQLuco0r9Gjp
kNDJ+YuEIXcfIT6eu6WDwvsmsDVTK7MBg6fr8okfCjA9USSIgy82kSt+yGZfOt7iq+8pgyDVDd4x
rxXmLN5kTgUxWkiLbjR8Fyw/yU68A3JcdVlJGRQHY/yj3JrX2PxYLrDddyG9dmbLy+XJTwznOWB7
FGMnfs0mLF42yfmuA2s3K5exZScasnHETKFDFudQn3JAK7UG/89lT1O70KVLph6NL0ZG74nQOZGL
pmXHrYT3GG0M19lRtur+UxwkqSJL9Rj17rn7swt1PrDATu4awjmnM3XLC/TdADq+as52iYKPX+js
ZNJ85eVDhFb506LPylxgl7Ad9ah/foR+GiX8l7j/7CMqvwhdno8iHuLKGUzxo1CyV4+KQmrprRto
WrYSOQmzbbAoc7+9Lew6kSsMmoRJ2l81Wriwj14b081EQlQKuXeEx0i7ELqluSGITHVS6fuT0TWW
u//Ptx9NtiWWi31GOEgo5IqeU4fYtw20pdu87PutVzxuCbIvtfNNzfA7Mf+gN7rG3lY7XZdN70mo
Oz6bLck1fksGPytREMJ5V6BpZr8EmwvxrP+FbtGIDNuCs0/yFbcKut78zYrJptEhyih4KbuD87gv
79PgEjM4LPZ+M7dh9MNqYKtv10et/05zmcHNBCCLCkySWVzPRs9aaXQDd+JLjc1HIkkG9i4UnnMl
p0kSzWX+X/dfjz9vo8+Q10/KgRvN6N+nuq+CW/LTSXnNx7hlcj0A1L2q6WKiSA4hq9NBB1xTFoSy
oR2jiwCP7FxULY9YCfmyHDfg0oDbGRUeGoE5DMOz4447Y2Bc2ZdKfjy/69mVvsqz5/sws4L8NmTV
MQhMuRp/VffpGOcKsy12mxUZvQnvopcnhKWJCC7qLny7yPmtwtuYjZYJkv0Yf0/BFvzpXYbkZyPo
jFtlB7BAxhBj0dDCK0GGXooI4rrvrCqIpfh1dg+JqUo1K4tIRzf0nw8DyFALVBXe/ieqA5/r9Y2f
Y6ur0xWHym9QSkUywZVnbm1uwDDOrh3ahMQCuoUDGq7Lk+wj1NOd7axAp2uKcii6phDPjIIMS+0Q
CwTWrCYoqcnUC5jtj8F9fWOyHZ128zzmAhiBDEslPoq0KQvyS5VS1YXS7/erZBKRm7PzkLOmNRzH
fiP2nI1KXdtv+xirqWJeuxStSSE1HPmmV1xFVks/NnXkxLV5UolPd3kUSyPRQnjRuG3vCzpSJMku
N0L2nzYwk9VqYLOPMfVvPA6zDRTBiHFF+syonOXrmm3dRvgeqnSatCFS8HRxkfeSM+oN84YPqCdT
RP6n/jkAB6YQZtby4gDzgBtpU75Qky22xy5Wk7jLOb2nMulamg1JSHMAC/eImVDa3U64FNhPiiwR
Q4GxP1w5KfTsSvtzfA2GeOUkPyjXP7udeWRwyxEZgUcdkD7QmbIxTwF9IxcSMFvQMXSy8AQdEWs0
4YsVhvL9a/8TaBIcJy6eeIAtQm841tuoonrEyDw0XAxceFYTYIcMA0IXaVQYlEZeHy9gbhnP6P2/
oQoV5laZuwLH5Q5+zNtvqhVqz8OhDlvjrcceLXOOI3QZvZ5fUm7tZXVLkFxwM8kZuVybmkhX900Y
8vg1tTJxJKlNy24V1fB9IuSa1rnTqYLMAw3f2XbYn4PhHB8Parr07GYVP4DgyXmhaN/C793BLRm/
yT/q63YX2th8h8+5VwP1rvZ+VwEVRVyIqFiQll8BAPu+6636CgPG1w+5Dlb2CJif2O77eMyvWC6E
edE5Nd08zwCTHBqk9Lr25wgmIbJm3E6ivUeHijsgROaOHGSMeukwKqPgCQ8+ylbmbqKr+5XG1vOf
cFdrUuidlowv/QcUA3NHNRN5Vl3rLVKGdJZacFoOZYCqdejxYEvSQ4xcqmX6Iry/OXplOgxc0zjV
I65f8dUZENw26zli8cWfUspcDAvgjVJ3dign/hP8f6aoZMoG1JAPbgj7+tWU9ImSbcvRIDQhg8Mv
JmnY0b5pdzs1i3BjAPSYoMM34n5KTaCPRuJYJtVDYe1QSB+E0zti8NynxsDIMUsraJwb3Vuqdoys
o8WxWk5mYRl3wqcmleWFALtyhP97PIDA1UpLTrzpSVez6aqUvv8JollXZ5Mol8kaRX09v/9MUJMH
hDvMyGG+r0dgALITDXnyA+1z34FGr49o0e31Gikggzz1kIQuhPJ60I0qQpw5xCu36+ujiA5DegJd
yT9rRUVTwoaGFXHUX792LgeqBUujjM43iW+ivHthAuXPDRSFvlDRWwTsHQclGyMPKYPn9X5MImP7
taEyMY7bd05OmN7SHg7NvUgb/rsA9xysP2frUOKaNh2fHz7cvDA/lbmX8Kuo+gj2RmvKTvrUebvG
i8q6/LhV9bABAYM6z00mmBYv3EunyWUQ+Q5Q55u/+Q5zgTNXydyndMnIMhTWnw/mZWDWhDnzZOY0
eS/yBuPUIGNeVyptOv5JxH8O1a31ReekQ74G5txIayyosREWksfc3rpZHE92BS9bXv/H7oAzLDtj
IA6t4nNyamXBaNVnJ3voB91PWWQIlXSOTpEBO2JgQ1IVQX62WOjHGC2u+AyakljRcI0xQZOB9zr8
oPaOAOK0s3r4XFRdh++obH8+G9Uadn6SvZjO7GH76rbes0e+2i+WVHPennIdAsDgYaBVrL5RaWnd
nxZirID8N/CDUAcu12tTF/qBCOj56W+GJwTPx7wdQFIWa9iSeY6twbRNsjY5NBx5bb+xoMXG23XT
ergnE8wbhI9jKXuHXqHqdE8433WXojtPGjmmDw6vBewpPflCFU33+Dzac4+LhyNBy6POICWK3FPd
A8FBYjOs9dzXlTYkcnLAe6LrW2VkDQpuAFq3NFyzsRzUahkxFQTP5p2f5vwEV3lVZeydgVFtCZuq
28qW2mUuCYPYaivcYexBm+off+iiMA2fC9fLdazKESxXxofENPznHUJDxqXQa1+dA6DPnr7OMygr
Aauoyqji3eeiEMM8Hb531HrGhYxmgd8Ke9HAw+yFjdRRbumF1rqGjlDMNzP2GufI0xnf2QgxgDGY
jNEluu7dSjQ/DARCjXFBSisXDgiR6eZclu6LejV8Pn2jetbVGZ8LwWDvyMwXKpyBxPCv8mR2e7A7
9uPeb+hY8eWVkNeIpXjWNYCnBnAJD48YWN0BakEFzGx7Wridv3WXNl3EPnnQRrf3LY+CvHxOXoVC
dFIlAe0tSlkhlUUx5g9snHaTfCyWZC6YH2JhqEUL0BgJ9J+rf4iPVyXGUBuL5ZzICa/RcxGUJrUh
4L02LMLln2dtC9y+5iyczuB64EyjEX61SFT+MR+ULmpJ2z7DUgQYGfby/Jqrg2tHjCUn3kOKY3+m
2LkeqzSID5amO0GhTmwSzLa9h6K7OPoR/TPKv7bbBEWIJf7zGJh4JerLI80tdOAFuq4ESwan6VBR
uZVVOlFvF/a9Zm3nekKYaLmSl/FVTnHV5SMfWLsXYXPJYqBAEf2S7+Mjiguvd1lr954tXgjgSaa+
5KpAb33l+wpiRRmsa428wXh+2zjV5m32yUA209ow11mClIVN5ooon2KYqBjaGMRFUFtxfuu1y5su
XM2K5y+zyo+tXnE0VDj1nSx/a0alM2EaUtW7HEq21psU/jKyf8UsQqulsVEttRPOj/VDgWz2jw3b
fRDy/o9bSCqyAsKF3I9nmgN423fzR4Rv/bQwDQwApIeoiR8X+y8VRPc3s3j3y4i8MlKoYj0sq9bF
IYGJagVr4E04AskXbPQ6L+NykxKX08IGqrkg7JWWZbU/0+adzyL+00WxgOdoRUkCq+uL7FOy/Bue
FesfaXjSzyq+8mjHO9I0kgA1gHprYP1GVPgkFKpoU+NL1goBYwO5RCpf7XMmFTjMxll7FsWIrO5y
NaWS7976ZjR2D37bgFo2LAQVglC60kKjSwbtdF8EZPj3ZZF9mwPyfsXXq+BruO7uPONhYYY56fR5
Lbmwxw1bR/skfG7XxS5zJaz6gB9OHwodlOE3Fze5wbkR0XKvj/NwOcgA+y4qYmzRTOlOSru+IfG2
lUMLCd3O7/fMXlV5xipWMoe5c4D6gh60Y47JSnNu8H6VNeEd6i4/NZAIgZcHfjyY7uhK29K0t7pq
PDx2ZcQlTBp+jyYUa1iEYUq5L7ZTQH2J2kJ0bm5UC5c8v7QBM/WFVSPCOCiaDeLROoqtF9eYkSnm
f2ybvAEHU9Bw1yiMm03DkHpAcuG77xzMkuyeMDcRkToVZhSN7Z6wVm0MUXq51UR+52jCsL0HNugd
wbYlWCB35SKzeuxLjWth0sq4QpCCUWozjhHn4kSnwLuQibdptYDI7hmwVWcH91K5MNNLANiqDf3R
yr8AGP/mAY/0RatuSMxplSopikMYQEAni2j+wIGUFcd4tNwn86L/HgMo+rTVRWxTiSyRpk+iGWzO
N07Q6Cp8jLWZxwd8JaI/6tOnk821WmwnwOl/ozvRU3x6fILeHkA2mWHcIOuvXPb2rrpg+/13dp1O
aQNuu1MWoTyGT4ynIkUPoFztDh3TGeCG9Oe4N1fjhY0BJDNM1jtfmwyDRtu6M0YGbpGA50PzPUao
obO3j5eq5AxhFKE4CjT5NapE4BxiQGs0GRNEJ+09JIVkgoFMth3Fmy56ztNqYpuKtBUGVWKnwZzP
+ht+po6R0N7cs4cC6BEn73Dcw8pMy77Ds9PUcQ5S3a/H6fsIJ0aD/f7LzZ0QaVBxc1VmvzYsbPiB
N/6vNRvBfOqIWaBQNKmHWH/TSynXlunERtU8rrCyM8Lc/kG3AZLqzZfkwTzBjq0tOt6zqUVLJFrJ
KcLP3PCE9LfHiiQdVrLxJ1kDlj+jCXl3Rh9ihDNQolW8To1jeA+KgtnWlt3bY0Hd5/sLyvDza+j4
FAEzRBpsYxnTc2K2HssjGR4vN7YidwRaOpfV1Uk+dsxm8nYWKiy1/KCHRo2q1Eh5puXKW6MuF+Yi
lXpk8+0aMI/x7k753/k+rt/9y/4tdYjXQZn+2m0VWnI5MNFqfQMxDJRJDN5rYOkaYM956dtYnV1o
4Pek8tbaXZMfMNceA70ZiQrNGckn+colnyAEWD0s5NsVFS9rBTUuuG9y4vWyWHJ6esPAC40eOR/3
JDMqWFqWjO3xKVD0JOa1I6teh5VQUqwxQU9g5pXLW1+EMdb2nQ8vBLisWKOGpPGOcQ72Ed0yQu/0
oan7zb3H8Ppp1YSVIZsJKhTY8a7+ywx9l4p6j8TRHDb/tYS148rGOPSBiqJ6P1o0tL8jIoT2Iq+W
L1Q6irhWOgfHo7jsQfFSLbcjqM26Mho2+zPI34c6jVGuUpbdv10n9wfpfdmJa0hXaVqb3m8TNHru
HtnhGB2daDAx4A9VOwD6NwBMBPOP5U0trwKCuWbfBiHM0cgeo8fUiY5/nWI+Vj21/Nr03XDNxoPO
zHCJPHQggfXEY5a2RWkq6eLxMAEYzpgG35U9J8i8L5iei9QUHSQshH/gspn2/1C2ivIrFe97yHZ1
4yEFyjBx29Q/y3e9Vi5/FZdIs+T47auHVGrD730TZ4rgtCkrpFta5cXfKht3ISZZmS9CveX9uvgF
BUYUlXmpHwXgDETlVnpB7OsDiKUFY9TqBGqSyPeqV96BzATJK+UbjT/EAeKg8l/S63uhWz8joK1r
ryEXmnb4FTY2RZJXWG+6S+nA8eIgPqi2ViX9aGJ58owy9gmjVpsftjNP3MvnsZg/pMVwfLNZyb4t
n46CFUvylypK3pD33w4EsC7qPUsw/VRahEh6nn8MCiWnvxy1kyt01Ly5wqq6x/Pcx1TZFufe0USz
qFw92l2rRDIWOyET4/gpwBrLjcMc+SODudlGFPG/1ej0DVfO3WLeW2iN/Zaoa77K8vPiVkPf1FaV
KfYgNrLdzDaJnlFxOOLFppZc4gvz6mogK/dOHIeGZ4J6S8ul0u4BMk4t4ezwT4QPhuBjh9sNQChh
lFjgClSPjvpUvocn/8wA4WWxu5o3EiAZRcog4QUYiSSJSid9+/cv8bIQPfxrd1Qq/YrumS9QdHME
Bt2dR1O9ATXbnUndhNTm4d8Yy7sjuMaohX01g18fyM2vuhqBBRUMe1eNPGFV4LsCTT/4A63mBzPJ
nG73na53Iw+yNx5zGDKbeS3ifY8bRy3rvPTrRat2LcAcDeSpLU8FiE0rXRnepR0dDbJhXX7G3m0N
zXo/Eue4sGq/Y3Ag2F/NIH4V4U8x6M3nVqseUnZhoYJ0YnZn2tFsXc7uVmGRRYAykJvHlZF6CNRe
lifW0gXadLBybGgGq4mdVYe79c/T4E6pwW7bNf4YZohSYtOVA/qJXEJv0p2Zql95PLLFIALQabma
fMrzUC+uxnPc9LVJs+DS+PkbDdV6rDpNeRmXjswEzDQViH6Lk8regoMc7lQZ4SHVi/lFy2SkdJFb
FHv/4TVde8YH27G91FoWfVcoG5br/Pp1Ykjim+Kl8U/Xq+R9kXLdb+KSmRs3C6rni6+syjzhDli4
wEOXskmYr03bs1uf0k+1cTbwaA3vRRFAO92QyCVeUyPzwCik+U6CADQh4EsVo6uUCIGi84IG1Gz/
Sgul6GYeg/EZQRbZXIXFfC6BMitdQDGsI8LAMEY1GlD98xi7gY8xdiQioQiAU2KzsDHpq+dLjv6i
DX/GWloUJJ3ix7XFccnKejNNXnH9zYykdDTd0Vsg34xm
`pragma protect end_protected
