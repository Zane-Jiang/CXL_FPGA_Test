// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
qqjiK3RJbUUDBgcgBDt6t48DEkBabzNorbNFsZ9E5jBcQL3agoOvNRBq5mWOCFR6
ebXvKC1RaelYPcKcuX8iAHUTkWvtplVrOb9uRGwSxLL9uTe90pkkcpe3xuK6zw3K
ZYp8uOSohEXvuPLZ7LR3DLOTy7gJ0tU9xBiVij4J0B0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 26032 )
`pragma protect data_block
T3q8k3zgrJoMzKcL1CvwNNojjKAPWfTApCbS0kLsUee268hsShutQ04ztFp9VK6l
xuME1t1vBwcSIbJImZDebuqE7BgU7QNrC02TiaapxQAzcnLPVxkxPtovYSazWKkL
Jp/BQh11vdGfY4I1OHlwhlNjnPNi8qZuz5HGlED6jrK/WIcXwOunUSk1mkKN6MtJ
VMRM2Ia++TZAChrXCbzH83vEmiyuglAxdyWjTaqe/qI/3CT4xCj4mvgI//MNzl02
FVO9iaEuNDkJdiC9UH2U7UoGQCL+inO42bCWKQq2vUI0PZ/V5qAxdFXfBMnsQk7F
D88AxVpixsXlu12LlVUWxDZ2oPPxuxZIQhqphF4xkPWcv9FCqB6f5U76YXHdkh8L
9ksliL5UuMVfn+5j+A28XTz3uX/67gNrXzlQ5Mdbs0fZ1nkHljyqZriFtA0p4c0N
te1qvVYAB7IT7aaVQeAV99ScuTmLrMmUtwmr8THTddwf5lCap2wDJ+DK1MaKkxHD
nHstRVNRNa2AOIBNsXbf1DsPzfJu2QzXR0JqfIHSkzULmYWmJZkibW6PV7qeEwwk
XBdXkSuoJOmQouuaouSfV5gDY1aEwphmGUVfb3VooKGsmQzEobd0B5hUBF31fiY/
vJBzRZdyDa2w8z9puy/xbWCGZNreuBKfWvk6Gl1VpUN9fRio5I3HEhckqGTZQdjj
aZX+36Wfs5BEPESxjrBzmKgC1b3FCpH1RekEXtCOr7uxca/TCJ7Ks9vzIPcp/Pjh
SgVug8+qT0BHecbHcTKpWkjfOMK+kfasuUMCaJkUAE4wJcY+L2OfSKUIMzo+tUWx
3j3QfJW0p/bu6AegkNK321TrFM3Rjwshiuxvn1sEpbXuebU01p6K/cPFaDZPWPJc
NkK+34xziJ7jqcbtjyLdfi/AWpuYVMBm6cWlGa8Q0Z5rn4CgPRwvQr61swIVuc5x
OgFVP2aUjdr6YyZbFxgZdn2ZQ3KaJYTdO039auevbFEuUbcHfwV8cWVBEmlTVIfw
2JPTJr4oIuDF8oqlmIr0PNphiBnLMX81wi5Vr8psBxOYHHdy49wGulSl2cH8I+0m
DlSMve8S/ypyV7lSsU2QNsO046dtXBNcDxZGquF1PLHM8LY8O+lz3F7r9ITRA9ke
QrzgN1weom7NKOmsO3nWYNHN7BB1kq6SKfbr+YDzQJFCMZm3i/z5/ZBTdsuMIVQ0
aoCCf/Ur1bc2i7g/GakCYJTdH7hHwSqdRCyOnNzCMBWcoVaTRVNw0TY6azfGuhbF
7p5g16pqwNeNzv3Csobd5aA6CvFo7W1Prt/oky8w+cxKjTfoL0coxd1MnMbw9Qi6
QeqjfjtM7mGIj+lfyQVNm11AR6cNUj2+dA6p5PVN5hLfv806YmFUgXFiyFHsvlDn
cUofeaPDnybpZrIiU4HyvA/2pLTQLo6hP6itdArTVaxiGM8UC/BWlI7ROvPEJfNV
7D42onrWJdhUHzALa7qNhH27yO0nu/nM6V/ysr9fLEEAkFYH6NSArAKkx7SEJR7G
9G9QwxCLzF2iMWs/CjREenKLQ/oeSYDoDYb+iJGCq2aG/MRK56i5fxFm+RdMpvne
xobbfCP1A7VW0rGvHZdbuusSoYoNXa+w3hGlsHmQ7IEFWm2LIeFTQcNl6f5ULwyl
NOvLoQyGoSfx944tYOMrkqGAXUVK77NHzUT/lTkAjZvBLjFt1x6pFhNMy5HHnt7m
5ghbGtyZY6dyIQUj3DZdICBTEMQYezgpW2LLMfI+dM6um21UxN8wAoodIzAYrQmy
F1/0IJnD96Jer4n154yQIF124+HtkWv5GGJKi4Zc0eqsukS7YHXeLSj48kEdWQ4i
hKUCfbcH6t1NbBYnou9gY0GP6Kf76k8mwMeT+aBNXN/CsWjVIkvGosyLlkYuTW6F
JolmmDOrVPbP1THY27Onpp9N2cMx5olzJLB+X+3JRiO4cSHo5JSICUVV09NRelIQ
tEgoJNq4tI2dTbqe+gOJuLt5ecoMSZHA4moCVC0iP/D/UiFPhXv8YjjWoFzK6vZk
R4zG/RJQyq6pCms0B9tiZNOOpNxsaGVckgRl6qm+7k4Bmt5HbyZvauCHLwn5skcC
lalwifx124R0SDUjnJ45aQLZG0WaSBa3e2f0a+2hV9juV6WHR6Dkt3imzLYiaSvy
b6XNnnBHm35tKACOlWQ/+L1/xRDQXsWa4/KQfU9N8gnjiaTf/p/eUgMe5OY84sc6
lMB4vj23KXncFXbKs9IEGMkAljbN/tu2JsYx4NUI9dpcMPo0+Cvpv10lt4dMV0py
ccY8Q8bccUnWyo/gh7TwsL9gCnMpOrEZg6YzuZHu02fHV0IeNkI04Oww2S+S0Q5D
zBsKrixsN3Q4oPWuz4TgCexERIDEX9Bcl7ltZQbZnomBHAFqaMSzMoFiRdDcFJrs
xmc8waj0C8hBb2qUyxzJuBSmUZUYpP8KQwElfaOWJIeg81FDECVj6RJx/iUs9XU3
ZEAvux07QpRJXPtCdu4zaFy/RhTfXT7OuEJuP9nVduZQPTYssUIcKA0u+hk5pz+O
FtDXxNpE7x3mnuxyRaHPUoKgpQHW83PN6MVkMvUn1qN32IDesuDvKJilhmvq1cxf
/6wDEjTaRQPdysiJUJemLwKO79jz9Z46IoBnjZt7kTSO/OQXsoENaA7X2vgcuxYa
NzZYPb37STTR3DYuCsqUUI+dhFPNvHdY6Jm3Xmc/+FvAaCYiTxYMJxdOP0bCHtaV
PQwCEUhTeMJgFXFGOoA/rCgYV56rR7eiaxgUbyUF7bGke4JWNWV2Brvpk37+0vUl
Hf1p1Wzhxk4qj/MvRVerNdx7Oj4B+5GzrTqZoRncoJXwlEguYxXAfvMFCrop4ufI
OzxiKOuJNhRT7MlLSDGJEAM6EQg5dLDYGzEQ87374ueCwKGW9kyFmEo7X77KMfzN
oAX0kgi/5PQv76Nt77iH7iYmYFl3m9qIrEqrndQIaT4VSpZxfekNsanuC2cvy6vZ
Ln/Yjf+IYOYZLvHNr8NRCRW9ZuKUWucW6Q6rO1QkFOmPFMltnhKmdwU5X9+Ftm1y
7AxOrB+Awn3jEQbw8wqFSjZ84AXeJrSLVsO7eyoUd8z3flCqeXj4DYip4osGP3uW
GF7457kNN6AMidqKqsMeNJkL3Y48gUn5+6cbyUArlHlhwjeQO9msMBgjLSQlI6j3
UqAiFMkC87Nxyymw5sy1jaWlwzegT6PImELB5QxZC/JSWpzZDeobdOJJIX2f7ae8
I0qs6Q9TZ7J+6udrp089kM0YdU84o/yZpbjZVLUZ5WZNLE4VagHqWEnfBDJAmvQi
/3tBGg8bsjDK0H68cqXnPSLUqG9kuX/qa8SCIsL+TeqQs5cJPp2i9WnZdVQ9zr9N
8RKY9LO0xCLn6yD0husl5Sqcl7V0cofMaHef0YDKkdHxbFsMp0Kj2ICPrMbEuoL2
FqtbfVVw7mEH9mIDKV8OUDN6dGcmwqLKrif16jN2Yp98SGIWe74fUv9ovo5lT4gu
LWeffIeTXyDtt5BcjRNjZ2qrGmggIQGUzpbD6aKwnk/j7twm0bXSAd3cx6fpk5UM
1fja9Z9DOSqYdNyweBQ1BO7b4lnvudnXbbX78uxs0ktzmd0kGl1PKJo5DMPouRgS
r4DrziHTB6/TwuvR7hrKwAPrMY20/FUeuF16vAl/AwNQtHGddwyUHZTrWEHM8y2q
pX5nN5Joq9ZYDSpM7tf6hCt9f0aHnzr/ELrIqq7WukHLjYjiJuc3+7/5tqz2JCmq
GSJMydhXFjxVads4L38PlUl8nP4W+2xK4uZHCyl6ZK9kse+C4PPVWfaGFB3RdvFt
DJeTPKC7FP1I1UW7NjU8WEwSiYS4WvENDdicSc4odnjExXcrcbLFPwTIlv7chfgi
Op6l/21IN97Ee2dmD3rAejwMcZj4wBqPwEw7BbfL3metjERfmoKoXGoJRXFdb8gE
VE3+/6/hzTo19Ad7HJyr6BxqLJw882yKxEmfy7b/UItZwq31YvgWBxebHJ+OhGNh
2eTcOIp7uVU6QSu+rdx9s7DkTwnumLnFyc5D8R4MfffROvcHAZchj3143u5F/y4d
YVGK1sKVZZHosAvSqOBhSbL3ie8JpkNSXvIMe1pTB60Fd10dYBVFlCBFESiZk+Rk
PWhAi+/BbWGhtZyYfm0O6JOi0HdL69hylvC5BuCKQzv1rPfKeGUckPO/hkRr9w2y
o9R+LVBP7hyqEdSw0VpXc88ImiZI035O1ki5YSwlWzqtSjPxEvjE6OIZZTZAD5Dn
isfBebYAlMRtjUfj8BiovbrS5pQHyGXyNDkvpph79QolNx/S2tMnGxJaqgR+8fRS
khVXh/9EphhXfZa4Z85WATc3d54y53tNkK4HakOTIAPjsSHxUHnQF3VIlUXku7Yv
EzpdV9zxUAiik1E+sFQlDAgxv1+OCu103Lw1uvz7/deWlHD+r+1avcUg0OEwJtm1
8DBe6olOrJ6Ea52GLKcLfAs28n/nEwYrNPgyB1Guv6WV2Dksn8/LjxwDbRdLkxKf
sQ//FSwz0ynmrGKt0XokViFEUbAj1BWuP6B70Xrua+jjj37GBeatIp5dOskD/lRF
cnvUcmfLsaYxcO406Sh9P6dpnciYKM9Yx97UDDtDOxlAgfO7ncaKdhwnywH5jvXh
kpnTKPQgRVTG7eFRv8qXaJ8Gvwy9GKUucuZptqIcWyiKfJRpy6iGylpx33Yx5eLI
FFaloRTZS60zNi5wDIz70CX/jmfmIuFjGPJ+V/7LCZTa0vI8LSCPCJ+XY+kfSy5+
ETaheQslaeOeJNoK5CCt19xfnMjsI3YceIPXXImtxATRgVRGDYyju3jtGWn/EVge
gFpj4MuwPiKNczSlmZDZZMr94h15zjdzYxlxVU9NddHAPsXbHUuNM3lT1f2q2ehl
HrQ4GshuByXAjW5jTFStAJMWbNf0Qipd8haA0iAPN/MDLKY7IjIVugwYDhd7XGzO
6kvVKoHywk8/w5aux4lR8JicCTP/EkZwQrzCrrHleDiR6k5X5NU9I7Yjl3tioM8n
et86auQi/XBKm+bQWUP1n/YUhRHrgvfCEeviEZEPt741M2WQxtKfdKjXbnpteR82
83ZbFolfGa4ht0EOdh9LeAqFnJLA+Rb0oyJUjXe+hMP3wE7d2C5wnw3dsenXJpjo
RV76TZi9CLC7u6Vr78N7Xfy2UaMyaDP4jTLplEqWVO2Rgi+AXep5y56dfR+yKajD
qL5iTk0vCzeHUhwrc/ll1INl554KQxio4nWyatrJnEtkOXAeMouYdUdtYzt9Xc/W
F4w7AcWVcUYVSynrd0/JY1+DNz0bk0kM4XVLrR4iz2ZL/5ZpqNJ6f2JEKHdICrUZ
zUELuD7qtB2aXZMOW0L7dRVEF4Sk33mCh/VyMDAbkah7cw3i3xgC7UIeKXnC4fNv
GCQ93/YHP0MPe3ZaA+VvNRIqvMGHpn3swJT/Yr6yNcn5cfE5J1LO2ePYYJWGMK9G
tSdPuBn4a/gqZH+JlfOLAJr/wbTU/Ep41rS9GwR+00woy/OQhOYKFlcXye6OEAaU
7HToKx1kPgf4USmw+Wjyciq+pxGTy7tPLM908m37nh1t04quXsgrk9NvPx1FGrUT
JsQcHzgBgouYDXXYGrSIaF/oEuo/5eXawbm5K9gHcqSoTo82FO0xMwzLAYBEGGoq
/l/6+71Vom2Pmrhk1bp1c/O1GNVR98ramOQZt/6RsxyDtUoJiLoQuxfVnNnI6gfk
JpZEJHYId5MhVbqgWtDi47FdNR+xrhVV73gtPR2Kj/9M9Ria0/1pUUlcjLq01acR
2cBDlDO0fpWoDjTw3DCEnCWoROKZQEVNup2ujowumk20IGt83bwRES0X+7dMcGuy
9CnnvEjM2GBcJW0boalOFMpgjL5+Be47u448WyNfIjfVv/9b4Ac+98soqbjF2uOJ
4HYQbQYbeoq5L1OyhQUf09Xufft68UOLRZ6MXuvUd1GLQ0n9L2q/ndYmUXsfVVx8
a2hv8tW27DcOd/sBc2MV15EB99MKv9kIRmPanQ4iZd8yFQLBKtpXRluAPB0gDnsp
AKwEh1lhm9NT+r2N240bs39DysGVSz0PwC9UZc+TF9lm6m7bq6kyySl2iR7r6UJp
2P8KG5jHs53kgw/2DUioRbVifX4zIF6yCIvWiWjs3UlCyJhmTG0AMPEBS9c7ac0I
je2VBgYEg8R8sz3CyHJ0N15r59EfhchOBhif33XthOiGx25gqpCPwhTTctLSJdSW
31+oX/pR2g/Ms3K4hXllsnAax/JwNm02ksxWAlD8CvGMW6e+DGHH0Xd98ZuEzuLd
UaDTa6G9Xsf9Z1huLQUBdSCF3fJhw95PWuOOAIyPBYP4+a80b+je9Yp49Z2rkalR
3vwhI2Ta3maXoh8HBHXa/ovAS3ZInNfZxKcTq4WbBv7o2VEQhAjk9aWpsgxPOhO2
G+uGo0vrZd0PXPIPBxNH7uJP/Xs8qM2rL7WGkea3GIev0egMrN3SYovoiFMnsIQn
rBZgTaafqIgO8Xt0JgoKW6LqmksaKKHgepLHblxzS/Z0RW2lOly1YKAURahrPeMw
eTZagyVoj6zrCBIQgsfD4vo6X2s9GQHfavuCgANutpO04qtK1xparVC+Ix7wYmTp
LWobHrYCLPxkeuk+5X/qSv/d2o6ZxgC77NgJmNxZaxTvIUhtvlKnHjdcCRrZMPGy
WJwOBMo2QqNuFVxqZ8yQ8wAML1yGWAE19U1UDd2rgxaZIy653s7h3zQONCiLqCFz
LlCk1dO8yz6iEvteJrIY1te0+QSwQ1RzhY8snSYsijfNy9PkWQTt8UzrmlUmNJ6i
1wxz0QAnW6+1q6wNwXejN4MyflYIUc2vJCBnVx0K1UYvseBK3cJVd0pSua2O/TAl
FcgBpRPZlb9BmiML0FGaEOzzt53QReX6oX/58CzriqlfTUM84Xaz02i66oXL0QSy
Qb8LpoxHt2qDxUMqsgS3LvcZytU6uuqc8hHzioY4lQmK2v4ADWTl1lFfhAMHRH9o
W3LdTQ056lfM+LhanShNcGaT5dIkHVrCfJ3yI5sIbsZR+ntgXvfcvYlJCpKasuyw
q67+cInhPgquc6mhAXWmhvbBHohBEOluGe+FmE6A6vfboev5SSRcSk/OFfV2+eO4
ONX6OhdBShXAHP0qrvftFbzONaqcYi6dXw0AuR0fp59uO2C+QRkidBkq1ob0pw+i
pIV/khsai8LSk8Hf5MaAgYG5YrEgCXP4e9+L2e+luvxvLTQIvcBli9Sz6psEF5gf
0NPwLpEXnfnMrbDoDRScBgiKmvZLdzU+9bxxSA1iAnlSXUUoUvEvouEYgJpb+697
wEoq0J8b/G6Gb03sRS64agbKS1Mk57S3Qw57LkrJKJOb2123Crq70H5xN5h0pIZx
p6lDPEwInFPGOGt3r6CJg+8uApk5w0NiUxkz1mU+oBNrdKYFzFvAG8Tzxtli2med
r3G+ibvqp53/+gJ0fwIIh/bIF1x/58VVzC+k5KbKSHfsoV2TlJiN382rGmIl/mkB
DIVPbbyCOEe1udOtxaekUufLnFNYVhbhzs3vGuFDOYxYLH+Eu9/J+6QEl5WrCwM1
QzY3deC9J9p7E8eYfac5c8KE+zFWKTiVfnJEkVkCbuzdk4ZlXtNg6HzWq4zen16Y
uBBcIpARM64/3RKgSVY6rz9Xc2JpfhzNskodzmnmeTKCf23K5Xi1+GzhbAPZ2Ru+
xFFrOv5iJbL0eyCqTTRNLbUd6ScKcUVHoNbtzk0ND9hs4lmudYC5rpJ7ffB8O9Su
jmk86jIRSyeGznkkVg7CzNBAJ8U+LdF7DWXzmNAK+TmWIvUu4lntsc6ByeHEb86L
WISB1gU+H4SLRDmV8e9tcdR0DB4U5+gzgt5sOo44hu9SjFlclRqlpM34guu7mIyZ
LSgEGQdV0PlIVsaLWABIot84afBgnsXT22rE1qCMMmyhdFvAlAwsHrLXJnUYO+dK
a+3uk39XPfBQ3UY9LHXgkq47+/Mf/IKc03BV9a61hCFaO8YC0LubYitV5cGNglzx
gbKEuWNJhY1+v1OL7CYT8SnoMP1R/f1YzLEXhHhQ09JV/ybnddWeJpSiOqnEOeYJ
PSxgROBltpVSzM9kfZrakUMY+JPtaPuk2oN6QETdptoZ+gL+aXWkyytwzZl75+Eh
Rut4x4NH2SGl5NdZKEDbmKL3xTu09tWkx6jQAjhMtoUUC5SbL+xSIqopL+e+0xiq
apJmOMQnevrBy+cWZONisLZmvn80o3Zg3mP2QvtSFEg7VYONpTRoFuC2ouVF9Y4v
TXadc2U2izdxASh5fZpfi6xECYygFs6mvUs5vLvcBA1YGQe/LO/VxnmBOKhYwBh+
qpyuc/WAW1w0yrZ39DaL0Ct5YW//8JQw4iArhJoIqFBXJToy0nPggJEKnSbAenNB
+6zW5+pFSS5Azj6hVEsbDvxNGbWqw4jPMdu0W2G4V81nzRuITRcA94fi8bHANKTt
VPXxrQy6oBBYEg33QE+DgmB9qv1hwXYq4OI5KeRoPr9MhHNt0VcCstbt6SPQ6vj0
HrhIcaMQBrDxB5qbxGVQag/EdnRwdllX6IUyb2mMymzk1Tuc32K0Xw97hHBauNNw
uUanWDddypNIs0wU5BuCmq8S45PKEkFgYO40zKV5Z/dw2iECum4YQr9NW5BFHvEI
5AQHvcypGu/qYNlrsi1k199D1wtUnKEZj1HT83jWb+0+HYK3CZ+pIiHD/ABN54zH
cVYTiqVb1007hACp3swKnvrVHHWEuna94p71ueOIj6xnAyhN314w/3RvienVuOUQ
yBt0wDbGC9JBH9N1bisQAwC+e+OqVB1ipuSlpYDZ3PAa8k4+CfXIEV2wDWZmBxtG
ylN8+Au/Fry++FDLY8iqj4TYUERFGHTI3tK7JU1VJNABeUUDOwxqA+IqvCEHRQ1j
MThAJkjzo/vg93Hs6ktnxu//qIb7PSL60v3vip176gAVOPtxewOjUcmxVekD72PJ
12IWn2G1/zv4BB8VcfmwVIzTBn21i0K3vLjYxi3SRs+LDJJXNCWahmVgJc6go5BI
VlGKBv9x4u2bvf/dWCx8bwWJ9+BpVGMVUUJX8E99CROuf4pwdhIvYZ/F+iHx2J64
9LdhROCLumQcHHjxTYaiG66gcrwf7YkoEnlJc2zreRhbngPC0DB+OXMdjJA5li/x
yjgrzutVYW/H0ATha8SmtfAuOud2UO2tOgvgJljBFV/915y6YZ3JDTuYuI9o0pfE
8eiL4YNHrLSlhEHm9gTuBySVxT0JKn2R1dl/kaGio5NXr6fgIW54oUM+kr6i3WX2
MChkxfo7dAdKnvd+825Kkfon86FN2cmtKXarWMDlEXUmQBOMfvTUE2lIsvbQZKou
ZPS2N4lCdiIq36tCJI4G5g0GYVyUUYr4VHZv/XPydYMwcML2XDVUiuafGRCt/HJi
u+Oxg6MSvrfpcueJ7w8cWl2iPYL4FKqRC6eNcm+iOWuoxT9BX/bNV8ryKoLl1TC5
hP9ffJrr7CYlPmkn5pJNeJgF8gn/9FvPrgqOWNGjxv5HjXoDXM5fJaLobMANNN2u
QsfVChmZUwT0QQek2xyfJ4U39ryQK5QO0yloICK8b1ts9uZHzD+6qcCDIM0f57n+
HYNqjf4gRzLZyorCl1BxvTGnL3xHLphS8KrdqIOlp/8dvC516F9e41L4xptpFP6c
x1ZUyHtXxM6HjCoXWwGc9eXxqIaaTKC0xJiLgnmea7c9b6Q4cpxLRDLiAsq/b4Sg
s8dgCfirYsVPHizrOanncH9dAQtJnfJ1LVlZDKRBjiVC9GTLCKNfpAT6Y2KFFbMJ
9UgtGLmt6oLizAwR5MkZxeTUwOyBdn05tVUgKhVFUNnWvaw0q1QQEmFvLWd+NxOu
CwKTHf7a/xADIdKfNXxvcO3JICTbE8GYSthUNoRTI62OTWZRVZk01s0qazAtQ/aN
dMNQ5IBFPfxU/02LKwxvadinK7+EpVyN165f/zH0wXV+eTPjNfIhM4+CtV4Xe3UB
fn8q4D5zTO/YrPwauMVOWlSw9/QU0X5Jp8LWPgZg4TzM1ZhmlUpV72R1rg3Xh9rZ
FFWS1x7P2i4AljN3p9Mr8pe5u4V9SL2uO+nVI9ijVbKACAwW1wny2w0kiGC4R7ix
M2IHWqyDDkgZ4KjiRxrif7LijQahroswZoaM7D9gOyNolWMKCZMxBEYbmYnmegBR
oDe15cJOVuGrSgQ4NQTXx2H42Ow1VYOHwBoHBuIOfNJ5USN/ONcylHh64RX3fVe9
iZZj/9JW1uvftZoDVEri2nmA4qzOGf1gHvIlSWigp8ppBNxkZguHpiFrSiTFUUww
iSzuxJhYil0r2cgkM4/xGwz/lUmfM5XgC1EfdadxrheehrcRlBDDSqfxxvQzA65z
1+7+bCmHaPNNTDFjxKG5AnJjnJgPE2SFNtkoyklFC56/anxG6wgyQVq1Q1rJJzoP
8ZEfBKiLWZhuxQXBTHdn1ePO4HpHSoOhytQ48BZuc1cyJRsi4d7wFWl6zvnhXSx6
l1WZD8LZcsipLIAGDtUgLlcP7K4+X/I2FKMZCYYW6HrtWYA1SNOkqC84LImdK+uR
+UAyW9tIZrWq+eMlx0jMvW1yHgHLhyUqRDhXfHQFDPb5qWrSJUh3NpP7CdwJvGaI
ZWs5bv0rrijd9uV5kwRQ25OiedCl2VlLfz2D9gR8wpvd+snkNZ2Yry0tKa17r4+k
xHDM1qaxMhyiIuIa/Q6yV1qbqJrGu4IYXHt+eIuT4Mia2qR0FzVRxuRFZI1mTgT/
j0+VsBHQC302hosWyVuFJDpPVak3W6j8NgJtGd1WjQfJN2hU5tiZzftk/5iwcLqJ
gjC+DuHzt/l79xEQKTumDaUac7GyN94EwQb7PbjrVJRU+7OiGDR1EKDJQrt0uEc9
5RTf5KsG+WQLNVctkHbkAqUfH64Hegk2Pl1NAs7HOf+xo8iYrPwkCYyGvTiifpBi
qtL2iJsybrcnKUcMGLfJk9jRF/ICKiJeZR0XG0S+/cG19knzzm5QWITFkX7UlP9g
WeCgHdlSeb/RnxtvQ9+ygx9553bCbLAQRUj5ZaT5+5u+pc4ZOcPVbN+WUIWbSBsn
lcuc7Bv50PSQ1NK2ZKjpYhhyCgdYQOa1Y6LQ/N05jK77Ge9W3jQgM1fqUqhXfMqp
Av2MuR5MUg6dsJKIdklPOS1M0sX7SQB9/GuuCO901fkEVYn5sfBPAFA6Q354n3Ig
sp/WSvv7iDGJiYHrOWB/Q3Ilonzs2/q7yALwQxPsrtCuP7IwVLkv2AJmjTPpPBQW
i4UmwD4RWNubEYqCWc2OdcgPCmbZQYmKsCA6Np5ofBnMlYf6CbVPk8mTvR3R9Pk7
tr9oabQStDB3mc/KqOxps9MpDLjTXmMnedmROSgULEZG88zAU38v/y6R/ct0yE+B
Uhwd758K/C+74MifQzN/3X8S5Xj9MoJ+IoLC/yc2deyvT8whP0AgnBHCKq9TuKVa
SImtYVTCOOaYWMpFkGuBmuVcEZL9+Nuz4H9bQwbOIh0WnxaNmiK+LS+dmtZc/EjZ
QUw9lwPbarta9s0OXKFz+jann6F4J9AkDq9r6EsuzreHkiHJPNGXYB/jk2XqCNpR
HJW+fRm3gSQh1zuDezUK7YWmqMtc4D9QCo4LbhLXLfHCBFBiOjs6nhOZws5+0j4p
fZWh5Q4emXnxObuDyUkU/LoBf0sOV0uiKsCLYzDTpda7e+WNgSkxZJg2tb5Z3MfC
63qoX4BkimJ8hSNeB6hJKsgYtV5TdSKpV7uuLuaNqEitmVbgmkXtPG9eehx7Q8jG
xJlm8HJ9ZkEf5VA/aJvIyBvOeNG3XfocYxFIQ3jQjsu/S9ssG0bFcK5p1rCKb0da
Sy8NfhJ1BU1JHlws0+tX64n3ev1FUjulJadKJIWAHL4f6KTW63Ctoplzl2NdI/e7
qG+rlBREAbd2FBtOrY39loI/OmJqKw4GHmSlnxE9Sw5byX0FcssXmAWFshEm7fjV
vYyKWg1YWiKTDL8a9sGgGTl2Q1PZwdczZu/+D2SRK+VpKalT8U9SGgBcu9/3KD/Z
Ua2Ct1BMo/Ru6Kil7fRJFHCY8RT7km/zKj/K0eoAyTqEuu8Vmv5qUBGe9kDa9EnV
v2OmaJfiDIc7/LyxWPzPMPbt7aXYpD51h/8WLxNJj5gqbVwEC2HFc6JvHHU0hsHl
wDC86kYpIf0yDNaGaYAP6Nk8vqQHbgvje4yfKRt9imTIucfF1mYQGnxYL8i2u8+X
eGa8ouEusCC9Fi0qxCTHoczqTR10N2D6wnZIAbWMoF9fPJyU35jmeBgXdge0hUf1
jeL1o0rjdRLYgcrrgodBt61/9U3hSTmnCcgcNNzpTabsKYARE/KVQnf2f2qi0ng1
E3yzo6Z4yz/fCcUw1VnPEi+Zg839J/t0G9RXWGwOi1x0dCGAnZLrcRlujBPig/nJ
9PyWBUIgNCBtcGW17yvcttAQzbE4UaSpgfokadXgpyUOfZDtToWnsgEGEkb0Rz/X
vLyxx3FBBDEBH40Il4b++W6iwv/qbjVX1WYoTR5XONK2jw1YMBVqncKD1Nqaax3N
/HR9g5BTb4WQIt+25XPKd62AIFA4aivXbPCRNS8pUPacmULQAwSkmtHDWnKWa04M
+9rOXRvUYVxdn3yqiR32WJ/Wr3CIQhog2aVtswPLjtWrNdwSDEso8ym+u6nBL0NH
kPFWO5dbrAhsdoUGkVu2YZ3r48AfKQRFxkP669hn+Kvv5V5/Z5h43d2M6wG0ePO2
zL4oPwiRZAEs9V2DOgivzyNjg2beG3LcJKrjeXbDEVh5L91J3Atbz2e0CynbNiX3
DStpLN/0Nfk2cCRv2hfJRmymkwr9hY9iJMRhXZUY/W+07h55XmurBxNrffBxNjvq
0sMiokCpx5bd5o7kk7zBMkngfVRVTdjh9+XEH9x4ZXnvqHB9Zju1HOzEC8u9A0a/
zZ7J6jQZWVLb4bdyBJZ/05gXwVtRO7LVR3qBVKHyXNR5uPJX5iSBHOoB82mH8Ycc
J2BshdmaBR17D5IwzYyuN/sJr4DpZ/hSaWD8Ms7WnkOJKKmki9gYOK+rWWxkx5rO
ZsyTgUW2Pn0BVFak7kBdNQQll/1Pdmmj+VBX1df/GfcBhJv+7wuWdXNdATL+p9Xc
69F3I0c9OasE+ux6XOL06eocnhlNi+WNhXFj5/M3UlAr6nkkQDi0rTsEpMBDm3p/
n0Obu9eV9BX8cfyZSxPnl2BV+UyA38xDEpQbCcwuBj4DyHtyu5EGqSS8PEbrkuYV
etuaucVzM+BtsSa0UXgio3ETRE9siObMNF5GorPj9yJPzQVsVz6IKmXnALXNUhBh
0a3eTxLweYQ+Ic0wP6lIMVXa1o0K1LbvmVdZ0aHotiWgVSGqY3O3QkxOdCoCVU9A
u7AN+mdVxAtqoYyRcjwy3RfQeINt0Ye01ZCXKNZNzjRZGAlggAdIWf8nRtiiUEZu
A/jBkSkA71e4dmyJxrFKnkZBcjfVrZTLkIKsSBnhJVbpIyVuU885arDxT4UIsmsW
GiznAR/Cb0cs6+IKi7i+BFFlgQahNZ1SmUw64ZEnrNt2mIC53gkeyYT1BLitEjqn
yGNeSmH+LqFtFfrgG6F7BaqJn1tKCDWLVPCi7d8ldhTiYSU8ov28mJEtbGHdCN35
wYxF6KNG9+YLOV85wk4SUYHjmhafvto7OGh79zzIm9/ArDCNH5rwByRO1jKuqJx+
t29cYrsoxFhzol+NIklizruBzH7nFT92A7CxujhiMri8UMj5yRsmcSwNWTEDS2i/
LpjgU/eZ+tbMfpHHgknHvhySPoLNqUVwokLR/+iFEOtiGQr9IEEVJtEl1CR0no/5
YgNzv6/3ksI6U0ej++2plMUoLaZlqGupCgzcq9yqPm9jfrmq3Cq+k1rhTwA/5gvr
LteqH/RUXqqs5wXxRYYjb0J4ciQCalRDfqSDN8ji++z1kBVdtfOnS7ka1Dd1aPlp
HJPyKk6PlO0hAPVYkC+w/F92/30BCaTJteBNtDIpO01xD5EO+jLUJNVTkhbKyWn4
Ezs6wVLkZtwnMz28KUSj+3WvP7PEVWR4VycUSTfG97eaITdkVMBPN2PUpL2RCl4M
Q2nhwmQ7t/k5QjD7QkOwtsgoKK+mo95uW2xDWJBb1aMJK7Wy1wrjE9HXKxbGLilz
bOt6KGG7aKbnZdegUXu0DmwYGjJgeXuciom3t0CUSJ+u9/9GMixyRqZno+y3CwyK
jKGl2ZYffakfEfRhKqP1lRaWO3ysUL/fV6KWjUC2MMYZoyRTWkUylTu7UtKvbX7q
7p7Jgy+NPl+87bglJYDRc+ZOAknCsK3NuKe6aLL4isT3zU4h4NBfpURrlhNK/j5E
ILaiyV3ho78QJ6F6YkectuTZV4wSidZYrA6QutiVMxQIyjmMXyr/O6c49vUMlEM5
15s5Y/QUokVtZwMgpUHlq/7xfDWr8X+2XQWoJF84iVmFN350PoXr6YN3UmR7AoWg
zoAibdXEK5OSv1S79Dwj1uXJ3IHgD8Iq19O0Pm4onzAuqkFtk2mrk76y3ZV37wMV
lEMiZJYN6JhrxCcCAsw1AbivSNTW8g/ari89ZbECYy+7FPunQJLg1Ietcad+gIgH
jXu9zv7JyOjpM/hc0+7zqnthV031xTSIViQWivsffeiawu2kSwWkSkY0VgxLUIsI
VVHWgCcZ0iWBOoXkCGEtoSBtIotzOoDBNcy/jcE2PaDF+Mb6rUG87F46V9JzG+/u
jM+Kp42Awx2CSJ9jxjvtQ6UNHPIsU/Iwrj1ualQvD2gtxZMzUBWVT8WBSOv+Dpbi
mxa+LjpLJ97qChCKY+jhQlASwS7HpupgR9QC1swyOOH97hPZ6oBv6aOfOWxSBW+O
fjJQdxdo7KffuC7Sc6n8/KOGKdhJUcGP5Zqq5A+6EaePTjybg5lvLC3FMepDDETp
J1BqTDNuplAHNcUCBY852/XvtPztxpCvAHY9WNw99FJ0A8B0IO5ewmMpfS4WBtfT
Tey7yOiTw9IJGQ9j5gnyR4PinuDFMPQW2sYkunNXs4wFyrf/ttgOdXItbHAkwZF9
FRFAFA/tI+dhp25plUAtLX2Y97JnaX+55/AyXPP8pcCAgeFADQ1J/8rbm3870rgm
axG4YetzCAdExqd2cc3TGchr7CHmLtKDYn1w7WscxjKxLvxumONkf/Yk2oeiP80M
2zGzMZX8WoAxYWVdJ/r7gdKrmPE/Am/PLTnrP15zFT4W2wTQQPLC3grLi8pu5JM9
DIf6wqvE/MD+sqQi2B+p1zPLD3x2WidumPJPovbFvOkmnHmZC3+qsIWei8O8c7C3
ua+ZWk8L4CvmaAxUo3wNP+5WX3RC4pjeIMbQpIdU5CT5YhezpI4vTB8Tc+SvNZ2D
IISOtp3Cdk+pF2RbX62yFhPedNdTan4jFvJD8lM7c/uakJCcMhxj1+f7dP7tQquy
7drRui3NAOFKJ5nSL87BbsvpCyrmu+VbLQaz7vd8JUc1VPGdq4TnHAgVds+whKlt
0dRTbRNjLQlNqjADJrVH0ZAqvsAlUJUlJrm3widAWlk47cqdJzA8BKpqmx5pjTjo
zMxPmk5eEKCxd6nz+ZAE5H10rB7p7YhQaXUmHRHgfyyox79QIs/jLVFoCRyXFC0w
cNGrGctjcf9zniXmia75Lqo/3M6gp1CyXs5yVnk8KKyCgbcIyNxqWVXMQYzWaG1O
mvS0bC19vOMV5X1sO539IRIqla/iEZN3anj7rENsSVqaCNdRYq6ZmVFXTw2Wl2gN
jXgDkbNqmVjudvJZUgZP4LCjhvrcHBwDAHtJcth+iClV1IsjqRY4PjAxPavaRTTq
1AZFQeswwsU0IiUvBXk3TOd4qeB1lAy53PGTtYf59adnqkFe3T7z1ECVd4qzT3nl
YORBemhPJwDNwkXoiqUS6iZxZdTumKQKqmLUUHD5WvbXUkT+k8hyWROmXpni415n
PP5Egojtw6/pYUhaXX+CQPZlWFuo2SWIMFhMuAVYpPVIJz6az4ki9spkVqG7MgLl
urjYGh5kpo7BaU/04fGQ4e9QIgZEGlobThBd/rBCGYqY+UBUfSehnQdjfO9CcvKo
fIXj7Qcws6GZTXgA6rNM0lgOgUjjgg8yHIGqePY01b4sX9U1+WETUf4Woczx4odM
+ooOkzH2XkWTTJG69mfznTRjF+t+pQAgUl2H+UHISzUSt4ce1oA2andQz8pmWBC+
7TRoXjopAeqLmiD+ysZi5krMn/bt3gBiHZ9AYWbTaGtOHtakWM0h3sKmFGH7WHiJ
msZ1TJxKvleafNxLI29ALP6/6RbtMbOYCjKJBhGuF1THSfmlfHxTDowQXpAgBQ3s
mJ9bidp4VtR2x3QXrtY9KfZULdFDCul59b4TXW/0NZJlE9oPjwm3BrD6QBMe3+PJ
5NzicagR+ID6DEq1D8oVDKfChXr0oC8lc9FCH7NRYZNbGbRN6LNOkCunKD4h3Gqy
7MQNXkDzOUnXbEgR7kT6U+AxrIoOLDTic1Uy5yYz4Q/Li8/bj0ytsa4XzfFxymqC
qVaCNLCsMoRKWslf++1ncyMEooKl7aJk6F6nNqFsMOxtOQMIXH6TFEXNCRhtvHri
9J7UFTBk2pcJo+pa7qjyjbHQ8OXTLhmO97cGXS+5WXOeTYdYHK6fbWg1M14/rlyJ
kQd/oLtMwaqa1ZVd8NNeiWpkhULQbYJ5byvTHN/SVnxY+QGOpsnuhrSfF10HAbX5
C1U6UaVxtPzXjJluP0HN0+f/B22AKf5kIFY7JwboQVt/sC5KotFEeYbWVf0amwbo
Oj8c/jMkxcaLL/EzQ1fRJIW1gVz55KdHKv0XWKgIPzaJ6OoHZphv/nlXCxvulQO2
Ol1Ik21Eofn/2CibnSa4XO+wE+ZimY6711K5R/DBhBz4RlSyE+Jbc5jLBB12pUR+
BoJH9/Te9Zw5wjV3xStGkZykeCjy2N/woQz9LrZJTokwsYdnATe6olywaDfE77pj
7et4Q9ZdxWp7quP2zMJD0sgl8b5Ex6/TzKJXp8Ysive8FIMkUXkezWDxNJEgWwpE
XQEBSiLRfmzAi013ICj9DRm53IpzxkwEkpwIHB+Hnr2+PatfCHQtKCrxPXJEakr+
2X6axdXtrsJDssTvOieR1WyxTJYIEK77/iMwbM9i0zYIbBbhDdVq0h/AIJMxpGE1
gxCMbjrlrczAvXcH9tawbSmNqIJmVJD3kQwwMbhkSh3LKFuBPm6Mv3514VHt1FTo
LEbwhG5ci/UH8uI04vNbJ2Mlpkj6hzY3AFq9xFmzYlgCPM1Z9z4e5r9E47RBF7xb
xvCS52TQaeQr6sNfwRvx3miSVYaBH2lAQ4V92j5DPjtC1edzo4ERQkcvZ2mViclE
HylE4s/yPFNPI5lRJBrMOFMjc/T08Owd3R2XH6MPbaYBbIwWCOKTG6JMcT3veW1z
rOcL74Ri8xi0BT9FjVGeBXvE9IPOAQzxcNnWhoAdsM8dWzHoChiBZbr16iTGIPP4
QNLz5xuCc1tM87Ipi/StJ9iBoucDb5uw394b66kEatiptTl02ZGgEIKSrxGIOWiZ
bISGxWzx9UPXCAgNJXXHXqeFlIW81VUvsrKFfR4tgyZiAIpYtad2rSCFn+8I2lmv
Ibni7SHvxg3vhiAnzpwEgNu9aqSj6nzqgQMRuwLcrqi7qvIjIv9bSLGMEkFQAG95
B601RuGpm9VQXKH7Fs3SKqox4Xfb1ckWxDaQSxGw7M45cmuUvRgaZGqKXzGfZc27
UNuyGgXOnBUUqXN7IKF408FJvQPPghxKxaGaerRBmEIB4Cum8vW1MZCvzwrJ7Plg
NYI5AFEYVlcF33nu39inJlvoGvHTc8KZyjw4Zvzavaq4rjPU7/nPSs3iakFGZcpX
4nUzWWdyst3RAAMLOs6BN2J3rqOADyTUnY/ugDOF/gFyCfYdwNbS0OqzgYYDQ3bF
MSl8MTwtAV5qy2P6fj8yK0acoqRJ5K+/vRCRnv728dilUOuzxgMfLI9DfMOK1hZg
6tMp6TkICorrLUK1rq8wsvtjT8/yi7kv7YzBCFZ4ilosgv+CLLGaCNpOQ5Wm9CqD
C7IyTDFq2hgIS5jT+aBh4Wvar8lXts7iI8kPpPrA1n50vuUYdGZMuc63VVd52JFL
vGCRLaluENRWH5a4BKiVUuQ7BZEBq64K6ThYhK2cE8+c607D1Rct1ErRAqESYxoc
vBoONzF59F40ozc7/bHUd+nqN17GtPJcN2zxsYC+E1DwZAqJDJhIRKZrm9SAEC1B
kCvDwBrb2kXJeSbRXpkyOG0Tt0/wUtWp8E3GCXrrJrGpeQe3dPu715uIDOV/Kxkd
Ovpm7X1k1TIwIdxo4jCKAmOzJDhlPTC1+yGUTfik0wUa2KEaEtzLtJZB4iokZZdw
Pwzcwv9qBEVbNOSqKvMwEQBw9QaCWfLfS0gJrEWmLlyvlJXq6+6K43K1VFvr+Az0
Wg4Jz2pjctrt4pDNTox6ZhhSjasis2NpAKVNydiUYb/8FEwbe1iaPnVwU0Jr16yK
YRQCrk0Uuu4nuNM0S3MHyH9+2lyjPc7ZyO6GGnNFgLCqw7Lh4FArVSohYc/DCLU6
R6/nN3t6m9p9Jr2lAFKGtDwMhpRJJjKSYK37wmRAgPBLuyLqyPClStYHe78WF36t
jqzdX8VcTws6mQ5fnGr1QXWYthhRM0hlPvObuU83Pr2QxOlwNYgBnjILBPRe9dHo
xo+kZNtxdy5F/VQ2FSC5wTJ4yn7YugPEUqCYHOc/fh/7tJa/XFjRgpgKT7mN2puD
ABB23VJFNfp7QbPAg9+vZOaRDyNiSd7eKz3FsCrH4Kw32Tlq3PZSXbmPrbo4PB9M
az2gpj6ubc2H/Ny4yqliO2kVe3CO4xASyY0GQOQdt9OLmVa0/L1wZptx6IJC1KCc
Ibtjw8aVOriPSgoB0VHG5C5jK4yzijT0AXOgTn2FFHwPeWH+VIbMhrR7yBuMg79l
DhkjAiGGq/tPI9kiY04YQESFCBq25NE6jW3z4AGtgdSVS8RbGBZA+vpqHjbNzJuE
vq6I7KXH6gz/kA2+1GOp2QpCvzjxcDQAugWECRO6gMbIp8LBj8U2MYvwkjHAXHpB
0KimlniJZDfM85OkZmXnjbo9ORAh1kmZloxR+FoIUoNIm/b0txZFbvldJU2dRBFF
tLE6y7wlKkFJtIiun5i8Yaao/xwrVHAplJm+vSOC5MRGDPfGuxLMYmwjzyUmnttC
Iw5QkwTbkg8IWkT4FzEbdaKRxN7+W7pA5alCKU1UJhv3QsEZTO+lJLJwzk0v41m4
FuSHJ+3ID0FjH51wZgbWL+nFcplQf2sKwIuUcGJKcTzyct0hcBGtBU5Axdd91qC6
2pcbh8ty5+7L/kaTBbuqmvi5Izew48v5YW6KzEwS+OWXACBCwdsgVrz3vN0/T22n
RFF+ZQo4VCS3xDBHag1zn8UmXKSRICYHSe8/4LVgUcWMdY27k7cFMIqKWTj2+Rig
ptKrzPXOz+VljRdlvsyGq6wIlEn/8qt6AXBCDMrC+f/zI+MDIWjJKReA3CoODUgO
ty7kR5+CsKnViiqx3oirolBdT6bpxyCEFuDrXLQ9MrcC7KgPZsD825qNBYck0NKM
lIA8dn1Y0LpBBwc7iwB7XLjzgjjzQddr1nZSx8ghvXRmcVyfoIql+GbxLnLZg8kF
tLqphQxQEA8YWYw2Yrri5BNIS8lsIlROLAZa9It55+VviJRznHveioFJUIwDlBRc
R7J/FKcjLQJ04gnC+00BoYfw1nvVHjg8aNEy0qxY03QAaxlguwOWYmcSXxyyeCkD
jku4qyfCnTeIStncwpvYumvPzbs/1x6vqM/KWsmIfEW8LqqYyQFQMzroX4Y7IGXu
5REJ7g3vzCKdBxF3EcxyjTygRLTd3z16U5BXb5L2ofQ/kCKcU9wkE7vlQ446E/PR
HfeTkh/7zj2TXUN+UEKZKm0763Xp3T0mzgS3YLrwpYMCBLv33AbEKb+gPyDSgRHl
Go/aT/NKG3XvQOYT4Zrmkbg77TxsIKtZBRXskOxZtSTNAbqYctRQl+1JYYgPtmqo
PlWduFIhxYObakATrn9ueLWoBEyyjjw7OIKanmUfQp5R4cwRvZzYoNlxWI88z/H9
Z/it9dlQkTP5EuvftI5CGPmc1IgFEPwafVJ9bNXqJfCBJWEu9CwGY5qCuNDSJg+v
l8asujqI+kW9jGBfsKvFvxd4LAF9llyZyD10o3PDQCYapQvmxjn0fa3uu+314mlx
udc8Ka49staK1Cn5miOSJlg1QMVtevSeRe++BIzZJWZWG9qspt4zucIydcKkRHDx
OyFZjKLeS7V7WhAXHXwB/im8fb1x2mLM8jjrwbf7NePI18Beiz5ANltOW63UNjVJ
Im61mXWDuASGTCAseQ8FRRFqluYyLF7jMtzkEZPfjIomN3Q/HSgxodFS684fTGdk
NpRFBPk+e3cvsd4/VkTs+VxtssA0c1PrSgYKq5+ZczHNBjRe6bPRCLRHYlEMZaux
Jdr+ZwnCQvHoIA7HVqWjvqboX60a1CMFySNGKQL6B9QjgctH5Ivycriy0nfJOjTO
3dvyT0r4+VkLy1+4QiEhPQk9RwAEiZuPTD8utURXZEA1xq9yWsglouuZIbzYV1Zp
3opow99llLRR+XFnjN4sPODO3nRPZ/0/VwGqOB2YWKqB2k7KpsZx7g5ZCHXzVFVe
Mje8pis6Nm1/8LlK7gAGTifN8s0Um5gulmoiAz2WrnWJnGeVEMP35lRZzZ2qfwN2
WISQ3JjeMK7xczxhNEmv7D2e+gRh538l7ei+h9WLLwS8wFrWQcXRgIVjsKUERUVA
/1Xdg49XwRh1qjWbX5uH0CiKSs/aikrrpWpndZEmMXN3SYmBu6suLcy3CapRw1hm
uz91zCorwk7L/2B65SoV4nYql/JELBZoq6tNL1FZPDSuCe4j4tm9AClZu1FLraXX
9QD9QjacDa5uCMVG5Yq3Aq3F720fk6LUOW5EkR7kLPcisu6meUt4PEbxeNKmUBNx
svxhm2zVizsbo0fYaOJEhNlvg7WTrEQ+yrOx29jf+IsbfLd6x+EStRL6vkvVrAwh
W0Cro1D/GMx+uykUnTVcHII9+FwMBtBGHOrsCKy/eVKP34IKQcshW5IhkMeoahKM
LQ3xiohbTstVfHf59o4m25OEUAkGxIMeOVtf4WGPfngctZKe5T+fhICqIvoXfhDL
3hhKA4DbdgdMId4CAK4XONqdjdjzHWL5O/tNyiCYN+nz1+fkblWO3Encg9fH1eBJ
88lraS8FUB6YEowKv4O5LIdRK/GiP/7e1PXZKQYiuJ4TPBbT/bxz0YuHErtrSn6m
pgUAPzhxkqqZtTtZMnhowcf9EyI8ChbYNpjW5BIiDqmS2LWs8nz2yMDM2TKa4U6l
6XgErych2REswn2ThWFUWqsAVmMEAbtqntrrtW3crOgqX2Ix+56uMTeMticKPGBR
1vKDMSvbW4ysx7+3Us8+XAp69WInop4oxrMAzqYFpfb2vFj3/yS4/sfpElVdygx4
i/fR0J+YL4Cn/NJddEIC0tIbUmskC52XaZ/XLyGT82TjH52xCVLmpW+Ao9DtbMWH
bPc+HE6K6MV4ymALCCnHiQdK2w1wAT+9xdOyk9+jB0p20+GrULpeo+PYsfCTmrtc
F5RQsAW85em+ZqRstNoYBhR6Bo6SBqw9OCNY6HsNBzRN3vTVaOQE6yeqx+RvpIh7
Dyh8RBr0tn8MyBpi9VnYBe41L9O0Cd+iojq+YMOUa4F8WUa3QMM84zigwe9LTfFd
dNQ5aESR/KkS+qh3ie7ohtIvVdR35lH+w6qvHXxh1ot6qDeN7Za1D5HCT+qe8ZF9
Qatw5SWNTAtjjB1mG9kbK9389+RC59aWWnWCn6frQhIS+IgA60Du+BGOuMGNAA5I
7XobbVMNB0xtb3cXCbzqmw/+HLIi38OQbLBn2a+tHqGLoGQX5jgsFb1BszmLyMON
q6fA7GWwHdGOsiLQI1zi3GBARg6a69DjwQgv8bOehUnIfGz0aSKCeiyq+dDNXghD
9vvoGEH1yUg4RBCo0XRdSp6hGq42391eZgSbNhsMd6JaM1IxI4/nH4GiQO8onVpC
1eqA9hP5E5UUsD3BdEjT32SSrpbNk9094fbFUqP9I1JrpNNG4VQMtPZG9kuM2FLG
TrTzuptI6i0hwhuEmuNpmoRyZ+ERlqntkdX6/+9qNM598ZtM9A+fvonh1C0BOKpK
agKrK2CEqgv5ECafA/IvKJbAiNAcWrUEUq3pV635bzDmvqYOYkv/B0lS55UEyHtm
GBsjazBHPgaWM3xHTxMdFP0j/fmHX8YkcCNDzSd5czroROLtFNA4Cmd8wx+KtIhn
9IIxYUHRfaF3X96c1/prrIJZxxYvjniv0vDob7VVpzKugH4wkBXkrzb8t8MDfW6O
soQ/2FE2on3KMmveMsFgSqWazI6HbzoOh1ZtoazoHqwqbY3H9RH+xlbk8M+3lji1
TGGLC3/11FB3hUPEJqAdHGauH1U2e7C9PujqtyKe/8JTzh/UE9jIXbsHzJiY+Nvt
/+VzyB9BpWSkyf1uxCIJxGAnSEEN2cXn9vEyQ6LjEmSvHALxJQ6Oq320Q8LK6DWt
4red+8YP0+L5sZfPhqMC1s2P9I+RdvlYPRF4XVypNtoqiMUHdTm94rhcw8KHN9U+
P/GHfby3IAfs9Xrw6oJk8JmBCD7ho84IdOmtxAyYVDmuDM34x22pqS4Feotipuay
aOyiyNRXV/td/zul55zBV9qmRnqDNnNbe17fJBZ0Hs3FOJb+G07jBDAzZ68jELDS
wAQ2T+bz8Dwui59l52uu3GUDPDBlATV+CqnwP27KERfu+MPV8zDSObqf0fCjNt8J
IkMZBhlbCEC9KFyPcnprZkNTv74cLeVp0n88rrQjOP2QYUx96NmJMwuks2eliteB
kvd32OllONbvMPzVVM6DaHty8Thl0jnZnjSLkoyNScNu5+efRYeXDd4W85DvzqEQ
lVg3flhj98iFwlgrndnUdf5OQOoqlEtPyDN0V11rPNF41hQWXI9PYv4/mxOxHTa7
sbA3UM7ZQvTaMY+nusYkrBijGFa3pTDTXGBW5aTZ/An+yPJC5fSBj7sY52YPzsCA
ETKYUae8svvq6t1g4ZNbflid32WYck2kTR6o2K/UMnPDYCDXMk7COoDzPxexcOER
PqJoXqcM97f7VgRFqbl3YgrFjTGOg1RPjQgqLF5MOEI35UVQaEiP/LGigvts9Q1m
Q21EDnug/i8HjI+mIoNB7mW/TbQAi1hbxX9sAboDsHnntA/8kl2/0X9POOsb6uPN
Rm0gk3xHRLP1vMJ3Ed6KBRzv41eQ2kSUigXU8cTUm0qp+z6/P5utgv8EkIKiVD0l
jOc+bT6c+YDj984fMLu8EED6NHfmdao0y1J5mhjzyv3PMA393DQK6Ne8vEvWnEL2
e4qzJo2ljfFF/CIniPgZcVKWWux4WmkU3EJFJLRZdeQIoYYOHevT8/1zcGjNNSwT
LFVs3t/btw9nbNVA2B9b6v9Xy2cpS2+0W2EEzqEHMt/zFP2L1+HtJCSYbRbSvuEH
WYW42xqmBkX1kBhhi7fLSEtKKoFRanCSdfnxQRE5o4CuCua/DCAMwt8arpld67Yc
nzNKJ8xLHCp5QAOlc46IcyeU3Xo085stndQscR2RJaIDRThxCRcG+DK0JDdZtZW+
ngypGQSZns1RjPhbQ9OM1D8hx+Q2AYRF12HKtHDL03RlZ6jeUUz6VNyeuYbiqynA
KeS8mYDO1qebHhGsdkAhp3AVLlWigNHs069gu7TOWDxvqs6QRz+WBmZEXhkhqugJ
a5kJv/L6tIKvMVRNWSap0zI10Ve8M2i2xdWtB+DIwlpLO2uZNBDMYlPXWw3KQgZd
yxY/QfUObaXDsxE5wUjtqdw8V4z7EHk9zJ8WS9XDtLCGwJBvd9ZJE4NqalbmHiOZ
B3fRON0IGDDodGDkRKcg5Ay4R6WB1HlNP347/Wp0tSk7eCy8mg34Pe6n24QuFyCg
eF4tTP6qUsWJfcscw/IjMxgXw7WYZtnDQFx9wod6zXoIwoOgapGPbmONfVkrBRSx
R0bNHO7g4jpTqZdpdpIzmPQ9aIF1k8SYvEe8wo6qDeZfpHiVcZm1eot35Tiy7ePX
LzSH5aJTNhl1Ivz2adw3oWSb1wJMU178FSmZrc9F09muUMqcUSaVC0dIejLWjzYZ
CFjHGI6ye0hK/9g1kzXUn1XrqNVrnuRXabF+eyea0AX+ueDlDxGPVRPiyFGMtTDL
tMUCcznhnjx4vxVlXTkXj7haLVwx5jB+OvInnCMB9Sl6HO2xgwRFPyCZQJbSxRP4
8JxgMObb9oRQ/XRSUB1XUbS3hP7JtjJ6MUA2jymo4nAgeuANa5gTFw076egnJAoP
Jt5HoS8sP56qahrKn4Her6QfUrDlsSIoZWVrgOrcWdO8D4AG/ikdiqjaxz4Ca1kj
IESZaA1s1YQ3Nk2gDzKtjTPL8ETfsTGvlUZ0+wKfE7kISiiyalq5BQ0eOSK4lqbg
fj909wwN8hmhItUMFlyOI8aa3/tTzvp2txM1hp/916Lc8L0JV4EEUSv/24MOxqxg
9mwn+mQjI/zUWHw+pMgCf4b1x/v/TpzZfkXbxh/Mf34ZDqRPwo0SYADNHep1MJ/+
+Rw24nORDBCm+ojEAKrW5mJDahi/ejvbY5w7fxJ6ROeg5WjuFwg3Gthgc3+RSHQY
iOJXkW7eOVRhHjB+RpwXAw9JbHJIzZmC85/6c6FzVkyjy7bgNLFsui8V4xYVgpFx
GkIGKtQoLVRk5WT2yeDElhYSClocHyfdZ585pibz7bKv+MWT8aG38QtCaXmRiJiE
MEiztMX1sP0nhpIDh/ySWxhPmdadWem683vz5RZwqzTD68vXdQVlgeLGift4YFT2
tvhrbVcOpx+nHttRLvFftkwWk0LPHDtc0bDX8TUuN5aNdofvb7kUiwa1SbXaU5Us
FAHJyyxUvSB0tGnzA8Et3VMSPftB1pkXCi5SaISfLxNyvxQvPnlzg3dmfMm7XD45
Lt0ZeDdQOHgmgZgiQ3BJIpPd2W4l0x59S5+ETGlDOBOg8AaVirIP0TWqyZ2Zc/U5
X3sqv9bhDY4oqQg3y1JDNZy5CLpJ/+5nyoI9e2yhBUOs9ap32ZlPWHBEcD0v7pz2
6DMPMjyOXSJg9POkCeEJXZ37xTbf/tal4asssDiwDRS/PnrkmjSQrK9qeen8ZD/p
oxaFboVPFxw/8QjksO82vSGF0vK/bG7EG68iFKwJS6c2LzWh7huwuwAxyvk/hmS3
jpmUCtFhSFZ1wc9wl+k72ao8yZ1jyRK5CDCRSggEueV/SvTI1jJ5/i8Rrk4QOiGD
HT84Ja/qs17JTQ8NFM0rxIHfm7CjtMB5VFjXELinXyrKAxQEkU8KwOA+BB32JUy0
+bd7vgTGGNYGNMACmtAj48qcTyJL7TC6wTXVhk4cxVS/t79jwx71UXj6hfuUXvZ4
VhWcNYAJ6GnJbGSnvoMPSyGN7SyuWkO7wlH5zc/VG5O70OPD1JjWLq/rYN9Hbm3S
KyP19tZJSFw0wjISS9cLMDH9Xesok8gZ0De/RdoB4AJITwnssNr3QKqbNBKXVP8I
YAuxwNzalHljprY3hKIiJfgdkh4Y5dbpUCcqEBFqngucc7zuTP4wtmsCUGKwURb8
+glTSLIJ8JCe+N+dW+A85vJsCoKRhhBiX53mv2+6WQkP4VQcf755XPIl/Zn7Xz8J
6BCYGUt3r+eiGSE92UJN0CI9DTTi09s1v+h/BlL/ef+9YYAD0VLqHjrmTpM+q1As
RygJqwcTxcUCgQ72mVpq4eA3NsyqoXNfU2CdvhH/iM+rG3kjJ5LzTz9710NVyBpw
K8CjJvKYngFfYub6uQ1L+Idf6aBA8/CKwMaDZkl5FcHe3NcnhMOl4PycxBjsBrZz
Bm7sJMkKfVG/NHErUFPvmZQoV8z25j3xKPeJOe9Zshts9Z4boDAKZta3hDIBRn9y
kNGXvqCQz6a2jGDFN8kteicdWdKcgYTxrI8oUKED6NzXvMSdGZzR6IjnRqxP/dh6
OViGVMV7aL/KquaI+iasTxQmgbySseNfBivXFtXNNnPsWzfCvRiefcVes6+AEaZZ
1JoiEfMQENRuGIa2gC8ABt1xp6RYgidSeiuP0DNa07U83E0Q0695bTDoi8CRhYcE
7Yed0t/H478ADH0zQcLXMo3KXnf4bIX4uUWKpQguK/lh2UdWvCHD7bcNzTd/w0S5
0eQWXwcy+bePaegCT/21u64BuRd9OZftTh8tOuzjHGj3R3Y33IhzqoBWYthvqqoz
Lhf1ktA/9NQ/ReimwV8OTT0FoH6vnclCelUxmxBXWItyT1JAI7FnTYg8/yFPq5Vi
I5+6QEV/PP7iBAzyInbF0VD3SB3tDKqDuFTOmlp5KJ8qnisF40eoqR19D9gYIKra
FuXdV6J/u2WCLRFzaEMxhuNCa4ZpB4apexOwKG8M4kiat9zIAwChIp5KcS7AHoVd
/FYbP5ZTG3FGnh9uj8F2m0ud+4V99LiLhS2etR5o2Q/Z/nER+hw8PX3KSEEnQTXi
W/7K9cdGA06Q+SEzFLJIidmcEd5x7GeuDzr+G3QRBPcVGk5X5xljbiYmUkje0c4w
lZ5z2RbcuH+IY94SnD4/wmbuz3AxLINR7+snB9K9nISSaeiZ2p4RP3uDwlvapyeJ
HkD17Vhf0ks/2iGfwc3amTD7CfZA4PHWhtunKZmr0mc1a/m5vRqAwXAhHeGw9nSn
S23m+fsMlrwaXp8QZY+CgGtDCC3Q6P4aoSk2cznbfW0pDOQTL26yMBryjzDcU80f
8PHZ89LwhU4Qb7sFQdfWkpCUGGKTN197xbcNcF7hvoDFaYCqB8dT/6UV3xCKCcou
W+PvosuiSBfngrgQ83sEwlALXyNidC4f+PP3+hfqpT7HvbXa98yp2fNWpCbXnjHx
JSv1SwrGFrNgDvwxVbRALTtFx5T/pbLR/f/Qz662J9Xz5kPsrJ3v54KTY8xnz+gW
m5S9au8uhF86II4ZFuHnIZ25y+oWudbXv1uk2l3M6KU7NFKYsyfSIfBg1HOkYppx
Vn15LWRiiGR2eMtgecReZImdvIhjXYyNRkp/6MpVDZTQ6W7+36N6OwTRlejh20WQ
8Q3eMGFt/WGOJCoJ8oXTP55HG2CFGDXmu57pWN0nHHw1tHkF3Vfzs3481+T3OXIK
oVKDruuio+5lnmxJMS+ycLQu/YRhQiq6wF6fhZg66BJMZHXfoF/5cBQeH7i/kYUp
nNvLxlr8zyCGGbushRNIkUivy+CtBFgMmh8fpJvlN1yQ1shrZOsI0M8KDDhVPUJm
jPjCwOKEqmHlKPyJKcuQf0EwamcPUFxAyJjthrHBpcsmp7PBen9xPvDnKSHdZrQN
7GegpTSSoG88WzE9B2XTuW/0U1N0GxL34t0tQqySP8yN33gpRRjPL4cHS4yVfkJU
PxfUG1p2VCnFsKQS4KTDjqk04He/1EgaG6BfZJz2FysCK9RhXHV3N8v4aVm/vT7b
1oc/HnA22X1H8ohUD6/vaveJYNUHE1R46UUe7oJnGVrdKPzLrN2XWCsjF5pPwF+T
pDs9xr/LVnoq5ZUYQ8yEEVEsStpjE2u4bZ2J+aytpIHTbKtYuVs0OSUlqRppeL2M
56BUwnGcRAVike0/d62RIIbFIcEHDKoUkqGQSFapae6F0mEJD3eT1KuygVHp1xgm
6B4+HPyDEqOk2NiPGg+ciCZn3sAkq9Xi+J2LTYEanypIKZ3xb0uXvJLRl65oNQIJ
46FL4lgQL7IlCwjsZWxG7JGWTdezOQuHGMRd9JmNuvl/8m38PsygMkOx/gsL4bit
z9K3AEfvg2cl4pYnxxc4i98WBizfCSKth8YPqY9FikbJ6p9DuTI0N2RSOKZ/eEP3
Peiiwf3yotZUYtKvKWt++2PXLrj1OLJGL2CDVyX5I3rs2VWtlRE5CY+TAkgLjrXj
RWSxbx2NTbiTT+/sr6PBZYCLeY6faiYqb40V/UyELHrKvCNh0W1xDcoNfCkHxD7F
a2a1hKQTpGDcWF83D9VxvuHBupBVmV5vqI39LiDA1yAUNiXU/4xRu6eVEZ3NMECs
ZRbv0bnkJXFGBubfdvJ9VNbz7ZOxpdSJlIn0oXnVKEh+dnFUObB5ornmipfTVKMX
Bg41p9sCqUWaAN7Y8sw3/FshwO8nkEHOGjF44aUTWUXgUPb41zfnuYJFg+OodHYe
pyLP/V3lWgyJOIOGwUGmCtuazRD3tlCyorttTp7bX8vxtMTsvGd22I1FiMVY+Pgz
XeUTBtP7zzsYhn8SyRdUhkrFYwAJJCBh20NRxKPpmHDr0ALqUAVnhkICeAFqPsks
xTbfxzSJA1CSKGzKIROgIUypug6TNh1gtRAjHJ4QBk00bh6EYjQZXwsULTEkZY6n
ws64VSlL4BHIaDZthrPYYw170jaEZMjdBjgJE7Heeto9h5M/kJyymMRCtEkATXUD
Pv2Qpf/wVXVUNoZROMcvRpPnOwAXLyyIgJ5Qkt23sEqZeYbf0TqOKen0ZE9N59/w
dThXFifnuqtx0VRXmGYudLhAyOJkHHhH/wbWdeU0jOf1ZH1UvWivtcqVIKKnxsj1
uT6uHJTIL3/mTYNPeNB6v162u77fE1OCtI+EXWJ1uAK2dr/ZJTB8/4QtzlkZ2437
36Z7gnu1D7tg3ZxK6t0eqa9oiFeAXUDanlTW2VT0bNpTt/+7OrQo4cot6qjkuPE+
yGC2CiBJviBgxhqBakR8v/QJSfm4e9LuNSA/YmfYdmGtIWBH1HqFkJY1o+UYMsGV
TF2V+N9O/wdMk6yqPdLnkyqaTaYkfKmfozNV2PwUMykdakYWRq92VxNM0iYXwt9D
GFGomT79PLzm4AkhpqibEjJJF255hCXYkP5/MoTKkO/bZmIp6wlLF9BXgWT5iGcb
cWyDPuy1/mtb/ByvQ1Hm98QGViEQVfIB4F+K7r2hmC3+wivrsdX2ZcH4C7XX1/u9
IOyRbkpK4Bj0FiuVX6106bkVeDcAgk/fOwwpTnDzEmFn/q9le26KwEbwE6HcpU8n
78j7WtsYqwZmMjXiNvlujwenQSx8RuZZJ7tlt25bU3JvfwCRsmZA2ce7lEPNjgsE
HQ9A7iDePi5I0RCVxhLN6vXmMg28ThHCsLa6EzFUG5FlNnukPvAch9EG5Nm9Pr1M
26BQ8LdXdlGDgKORXrzh37dN3phlNpML+vW1e3OLiWcJqWM2UJpzYYWHtu9X3U4z
EVxVzVIkQMjDdgSpcNt8IzTTt5/VSgfL+BSE4bxed5Wm971Jr/vAhTNiR3+hQIIm
6BpJiAUsa5j5cqvxFsOgTjWZv1AJS0JnBH98e7v8MBNPlSfxA+JPcFBy/AQERr/D
YMChf5FJa+8IyVoxYaeIkvLXJgSlI07G1K1CD98SLcjI8LEUCJaWCFWwhWuaxhHb
vimWJ+UvXnjhV3RwIcc9OMClyGezFV9TXwfm6MXCk7N4HWgM9+5rNLIu3s4x2r4N
648bhBLuLVcZsmDAk34YkkoyCpWAZI4SyFeUvxbU/x64KI5GmflyQPQqIwd8OdmL
NAGxppCKdsslUkmJoWDqDYM4XhVtuU3o6UGyd4L2Ar5/KiPrSahLPk1DOPJIiWEj
EpzEnG8Q5DSTpU1GrLdm3gxrlZxGxtbiLmPqlQyNTiYF0yksl5i2jEJkRA9f8tpV
yi3njCsROt6547hpeDYxCQGQ1RifhBdVnsi8vkrQSANeS/8/5717cjDxPAtJcSLX
I8dwBh4r2mp9uuO99szes3A1asPK1jz2d+dZH5r5EoDPwRW6EL2JsZ1Wv/M8deGo
jjiFkFDgnmd2zzp5EIHheJcDN5JvvObj/VTMsK9J46b6Lmq3n2PPTQWoLvwkYGuZ
IKetqPsrbJfM6t0i+yumoEOvP5oSTfRdXaTK/31iduhaVQ4dg/GxeHwazvNXegFc
rF+aZyAzYh7Sk7OFJ4W0Xm56oKyM7Id/E2ifW5UQhxITd1WN6+Eq6cNAXVBVbxb8
FbnOiPInd5I5SOODou/sFcmx0zuCgiPQwzltzM3SdqLjC7R5bFOBfC/9efvmCun6
p6udWEMtyYju4+CbXeIbdwacbHTjBahXmvVC7eg4O3fCBvPBdwlHxN7BEEP4AgUi
DqXyUFkoZWAkx2sc/LRGzZXHES0tih5gSdZwUFTT7bdofa98jhZpYZkK+p4ZGNEl
QhgTm4JEqnkGIT352WbyFCdy5xBxY6Czgl9W3qm2DvVHgmf5WFkjgT4GkuJyvdDy
GKg4pmOwjkR4YfwPZp6KaKTqPFFpZhr4TFf9U7Kp0XzkgugkKzlBQ6Z/9ty2qyVE
oR1x8zE49s1GdwVl9AyDeKsv3h225pRKNypBd8UXekmfJFIKauxBWdy3zGJI3ZGw
T3CeB/MtNhxo4owmr8tvt9FL1D3hZCqwrQ01io7SZblA+YN5IR0ncC/iZVkFDqgE
7FdPmPlb0RQm+HETBzQExkVMYJiTZU94CVJyAdv0BbbMt56BUSERCKdI7uQnNNC3
YYhAMsUaN+elu4+EriioQDTfKMU/O62GcLBAKc01FzTSqoorTdnRwwSImWySqo3x
T2tl5dWC0KSbTOLevcVdxrpovRZc8vkKJRD6cRCdc2V9FB6oNIivR8MwCaaac9OR
toQ9H3yyoCR+VitLDIsqfc/SWdzoFsVM0M1ME8Az42Ye3iYne0mbdcmVCf5PMiS/
s7i5AoFySRff12RYtGjXFrHFZgDqb94nOqf47oq637/v4iJuDq+hN6kEivMhqM0M
ldHNO9IBOGNtHWWv1j4ZAGKaf/uiwInl2IKnVqYpGb1KARVYxXCbD6qTz1ZJyHCJ
ldcL+/Akufqi5PwgvUTw7PJQkdBsQB4xk6gflCbi2IJpEyo/iFDKfjjzh35qjJH7
J8CJdR61JNTmrr+CAmDbUSI8WKimJyXXRwxsULTVUjcNF7GDG/NWDbiswNY1AXTJ
gYZ1GqDSAMXPIm060TgE1rjDMIfU76J1Tz/dloVWnkXW30hyhAzK+85++mEW8+Ky
saalAkmB+jql01kG/abcBAF6kOj+QEexi7UpBsDjBln3j5iOlo7YgiTt7SZUUidr
s1+AJD/vcCc1mojKe2j/KPCBAz3W8ISnyOB+pSplaR18dv6j/ECX0LXKLmCdtJ8y
oirfr+2Gemp2IYB6+x3Ot2J220bRkI2WGquUazFUL3qRi9ogNZxRN27ruqSRiUvN
hfZjpGTsFLlc5k+7LVmcc9+Ri//m8pBqankn2Imw1SJqWnwmoyq5dmz0v6og5jFA
p1DEMbiWj98ghFTPp3f1LgmhaIgzhuGtkQE2FuSXW2nGeVZpQH6ax92sR/ubtUsO
8GpfCCwdLnb/+iOmxAq48pUmlvJ/AvULGnfTbbt6Z2uoj+WNuN1kuP2v6F1Xwf41
kTseQlsILwbbKRfD/Sfgfzfm9463WyhH2t6DrEITV0FemjGbqSckAJ3JaR95hFW3
CU7BEecgp434NC1J3a6JjQ6BGsiiPLYD6wlq13q4SGhIOOU1PwIBE0pvryPlsKuG
5704XmfqgNQfHQ7tcd0J8J63JArOrb/tYvAfVnpUJ/J1ZC2cHwO2qHEISG+GxCRL
vNTjeLS6LGRwvtCKOWFtBj1NQzTW+0dRFz+VOQn0gheOv4S4U0eqAr4/vHE55Dx7
w0Yp6bM3CgAPtz8bfMhz5dS3DZTTzZh0ZVT/Zvu7z+IRXmlxFcrK0pYrpsTKgkeU
xk3/jVT0kcO+Hv9DLOrEUJxfkgWWWkOO0L1r/0CVc8+8e9IJhHyaPwndnrj190hZ
0RDl7/ePyANJ6h6JAldT55XF15SgaeEO9o9q4miCNi4jwzadcvC9/bRkrjaylKHD
IXoqXIqvnFTmfYzUbn4651DdnLppijJ+2H0NRaNh1s97mHWT2AWpehQo5qjr6PoD
61Urgd2sFMsjRk4X2NxiNyHFg5NSw0XEhHIhqY6wOrAPa6SrbyPHnTtYlaCr/VKd
fxVXUJa2NeaJJ6jTAbpbT7LaQAKEcnnXXfpEcaMZWHPfEY4vTQ/wSnSN8acfxo8D
WkllyYfSMqHFCbAWW5XPdL8HD2vwXW3vXuh9i7ybI3jVbymegbiuNO2vJqMrwl9s
7Y2zb27cUer53voH7TVVkFeNJvY/rN9VWd31UZz4wq3sRMsJZD3rs6Jwcs7uW26Q
eMS6+9OBE99jyVxCM4D4dnu0WHOcoEfEfNNg9PJv1pDNVeIpz6WpymnFocY1EvqT
kVN2VT6o/hVQMdXnqUbawQzD+ByJUe1x0h8q1Ay3FuagVL9boOf2GLuTkoquXEym
sSYR98yj7X1RxuDnliqFUBcX8BT4gUg0DVvU35em11KchTswklenFPRyJhxSp7o4
EL7MMHHMvGGjuEWDzsBOkKuRoTx6dLhVBQU5MKUKDJL6HdysCoMDQKXd2QfazC78
YBSQYtGV/b5kkcfOsEuFNkZvS49x99VljHcVE4dfJyYRMj4MIhxwVR4UpEQF84C8
VnyNSdJrWroksYJAUI2euIrRzFBfgBKgDrcf6X8XIunjJz87cYMw6v2ex7kTTZOg
ax9F8dDENCGUQxegwcGpguggbkHHfzNIXnjGmagvIHX4uP50HT0XJ8HotWvnJmcQ
itui3tI/hnKQW1vUV/PA3cOxgTF0hKZnQLPrvNQLO+Ub73hKP0NQ9jR7PrSjVIf3
fNPK9/SBk+R7fBPccvqgpnEXzqoGelHtaLIecufSNAOrRP9gIs6togqpevQOcHPo
A5TXKohY1CfEvkc1ZmvW5/HF4WlOBtKieDMfNamFyZ7qp7l1Bz5GenRHbv9R5yJM
I8RL0v4IbGGpV7c6ldb9RijbStP6bOs9xUFs1N2I+GL2yCYKNpuuCDK+UsjWVx/7
C3B1XUh5jc5Qk//7cM4FIR8C9U6duiOzFXaUj6ge02cJs3h1x9F04S30NM8oEUey
sVWu+vn/p0IKjYbf7KsKvNWqVeqVUeRi3Jm+x/u0h4vmoDHydWMDqCSkfqcVW5zV
6CPcuRU6N5EW3DySLIZAyTMpGPzohT3Li9re1jEZ60tFp31qnoeIKIvF/7YfWZoq
fL3jQuTNqogeEei/G/X/dIQcvRcgj/S6joaWDZ81tkHAsY5kwVoVDTfny+6kf7i7
XdvzRrcns6iH0bckFQJx/FaNRP6eFYDhbVqBiGqEULgB7m8AkBr4MLMyX2itCI6B
H8EDhTz/jccDz0caMTXP5ncM4m9dsBAW4+vZEM20p3i8d41qtB0WyPygT+O3So+X
fCNWXJ7M1QtQnPeojCDygYTp0/MMAexcs2Nu8OoW9g1xRsRU+zEdwx9NMmGJS4h5
M8wg63QKyIc7BEz7JIb6bjonQN2O/FIlfWkJEJpT8eV7xarsxP+SyGvRPCczOBZt
legZz6nGZ8h/Dr1nrgzydvZGzWm9eCOBbJKA4xLY+uryE6CneyFb0O4s2qwpFqeG
6btrLzM8dJlfERI7h1opDk9xBTzn88oLeVWRAe3NLBRSPbUPNc5tuEzQLXWJWiHh
PI8l7Y0mcgZ33+4E3sNGlKm5uNtjmRldELHEci+24QTxbrIWPKIIDtX+7F5MOsJE
K0jpzfIeTGYRrKJcwlNMbhT71yPdZ+FP1ngxbiA5x9wbMQKJfYbxJ+WhgvUpdasi
cNdeYqYNvX1T2BdYNtNW69RAAmsgt85lwJ0kW3Bhx4FWeOaXgCqEK2zZu0lzLGYT
HsYnKYAg2cfZW5GOBBPNqsPbVUQmQ9Y77/bDAjbcllhLQ6bWSmgV/g2j6as4Rad3
aXEyLszhg1LVm0z2ebT5s+O73Pk0U679+Te355quy0HluqkNVdK2O+/vfak06oWi
1WR8A+OlSA2V0N3VJ27r4nAWTxM4MlsfRiuz1yg6/LnltFbxityiiO8qiRLDTL6c
WdAZX2YV0qBs800IQ3VzfQkAD8s3D9k77etwZiL3mWGDpQq1Lwj9QZPoOLxSH85l
PfHjTMlSKdHIulte9XaVN6vHILJdGG57QhZ2ydOspG+OGBkWZBzII2QHP4H3M91V
s9PLrWPFobCLnf/s+vOjCz5J6g1LqQLTpMUg30J9jJBoNbszFoU7Z4UAUv6VchHh
dKSKLQaPdklg94YTBdNSS2iXyMR4sMlVp9KZZXE+Rpmcm7YFm/Y/p6K8lKaH1uHc
v/gt6Ks2v7eLwPiAq3jrdTDcLS2pb0BoPdoSooHXrOE/exNQ9mt93iht4VFKEla4
ubbmMTKECYwS9z3g8YCKYPC4tRkcsJgdPazvzviUU4EofYjuY+H0WIBkS+oH/7zu
MjSTeQ+6VR2V08mKnJgDgj7/hKB7xBZxqTIYcMPPZM6rHUo9lNaiBf5MZV9n28i3
IoAaufCt7A1Zcq+xNwgn3Hu+vqAOU2JMIatGRg5/MyPURdgyOwQZMj9U8Ba9s6a/
pjKIA9cR1QkL1p28+JdcnefssvLfxETQjz6OTMG66POyMihA+LoBcAOzsLEOQet/
wUNatoTzc50Y0cu0thXAPRSEJuVQdpRR7oII1sp+5y0hPmPfEA13LxoQxOw0N2b2
lIjmo6S5D7JnS2BXpbHPplsjjoygYIVnrzZetw3Qe48eA/rroa63xmxBxCsgJKJ2
litB03o8uXoNk+1dt5avKg==

`pragma protect end_protected
