// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
JCqzDbTRAXBNYBttH7mXM9487PoyyxBfS3QiksC0QyRPJ/bYjv6tT0JUt95w5EX9
AYcSiDwH0NdgyhxY/9OJQkxi2UWvtTtiE0RmryCFt5t751IhgIAvvmuDqlS4s1FA
Ap4eSKhaD0xxMq1qI12dohgBZAhjikP3A2ESECHhquQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1584 )
`pragma protect data_block
P5whtzKxqc1MEqt5k/gqPVNlizY6iODNtG48JSin+wbkPsoP4WQ80OtMpgBBc4jb
6t665NbiqDSe33p6t6LYSNaevtcx4jh9QTTIO3DopWe6Nsr+dj3qYq1NG/CTM411
2eNvizwbjV5sIMwmHFrmWk+ChDqf7CdCXEWJOqqjSE1+6oKbLJeO1i1gbGLQU1IQ
J+h5aKfrOllB2fZ4EEBO1j0rOrqEfuJOvqVXJkMdrXDXm593NmwV07reAgTjkQpv
xPdseIlxc6JQ/pdVslw34pUyv7fFEP34q4J9O8o89PZBGs7KfHmSm2xYNEdygNc4
KTJvAsITdSSG47FwKm7jI92BNYCQgklWFrjOU8Jv/8bn9pTlmVlCkvyHZ7ICaHHr
A5cZBLjwQZ08V4OdjHDwIkvlyuBmfCCafCAGck5/aBaKFfj/5zdiion20uvyeU0p
4wLmW8gvh6/LMVg0Oij05XEppahmKUxwi2/492+E83SqvJt/rx2o8Xr9hVjK6+AD
HpMvOiYqv3JfqrJt6PeB5v9wL+7YACxRnD+bxj5Ug9qw3vQQDNcLa0gtRg17NITl
xxhB7oh8CpGzQ3w8YQgf7ZkRFSXJAFPoGAh4OS55Za5mueJ/dgUpPy8F1VBMUW5S
xAYgb866JP4ZoiWuE9DwaIr6dk1ZXfw8jHOH7fo+DOFpYmlEBRXNqt1DYqX4dIe8
O6mm8La9zItJpUZCQhLVZuGm3jlM0QOP0o+4j+DCQfzI8B6p1BFPvWuunUQ2+5Ap
zqLLbvuqal3psg1FhWojM3Zeov9xSDpDGe2rgePbXDjOl351dUcxSlXEufdkn9TC
Bo5RrrTPAixdlVHgOXqBbxlC1/tGsdpVFf91oTXM3ypXd8v/iDE9PP+zghgTPaF4
82mliNpfctUgL1TkufLEXjdR9niGAnQNhj7bM0QnyNRU7Wi8x2HI6qgvMfX2Wwlo
pWaQWRi8zS7cX75hDjb2F1gSRfaeDnkuu7EUA28BDLNhKvUDdjt9DMsQr/iK3T8p
j670cqpQbtY7UB/oqT8vLEF+HT+ZQ/D+SlhuR4tom7zOLUQITHmp0BafWWXIy2kw
4J+m785uxmUdJI9BZ3a19R6n7W9KzaPMkqrl3PtYi91LSGMNrXFIxkrVpe063fED
3f1FIsdHBNughvW0FzPr7YS5IyHhhm46nCqPx3PdSjSSYfjJfDXIAoE5WiSU/16Z
WL4N54SHN6MrbqFFZZTIeTdZl87ZabxltytbRkGqDxoWJ1vAlUWXldjeHYIhhuT3
5+XaC1U5rbnuJARrWdHkS0DA2e0fFGGXw0n/LZXDLOSdlbI/r0HTokCw2Nw/FPOK
QsflpoJEMnYs3HFBlE457DazvMVN07iOoyCRgu9YWVV35KKTa1H4LGatEKo23hva
bxRcSrE0HahUJaeAkXwy2HD1w6jjeq/rN6W41hB2JW5Ux3fv/ro1YcxWQS2TuumP
FNOwoCVbeTpk9XnTK2i5dTJ97rjq8fk5mVYzRKKRNIjDWCxzSagktEEOuVaxJcl+
Bj+OUx0tFPX7wD/uUMRPod4vYuGpxFVxW8Xq32V5gfG7qWzJMJKY6Tluk64O70iR
4Rz39G5xdsMUkPcU/utJS6rNB8la9jUPZaq8i6mOM/QeRmNuHsNTMr0M0L6DtfLS
J3FR3P5vaHRRxG/9jxS/CIxEaAMUYm8GiDEJ+T7GjfsbDjkCuvvtZ3hddC3jpEXI
ibqs7rd2Tf/ogTX0sLXbwGFQ8la6Dj7Kl7vvpOMWL6+G5nGqluVenc7HDT1bzek9
WPiwMVyODqus2JGNNPpKEWXS4oMGzif4wdeYHVM8eJ9Hjqq0VtYbhExPOUBUeASM
0vBygZsYvX0yL+bjjx4t2bpP3yvHRsNcemyJcmu6ygLWdu/jWSZClbvam0YCFIgV
j9WjWh0HHG/X77W/Vj6di6V4GlAEoOdfdJyXxd3DAS1AVVmX0fQwYuXBX+nNbxW2
xs9n+xln5hNzVVhKP4a5NwioVmLsVQ68Q2H41UoVFclaTsRQXnGXmjvYbq5L/cp/
/FlUIWNz+3WdJ9TfDLyqMLignH5J6LgtF7/QhwbhA/dfpDkNXzhDILA1czhn0UJe

`pragma protect end_protected
