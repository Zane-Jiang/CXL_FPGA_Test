// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jT1LO1tnc1ei2aH7WBBCCX2XEENbSt9hvtBVt68pgCR1T3VfkjFRLt0aPvW6
RV02n7xAEOdlqKbrhSfoEN4zblH4NtMtQHo+aF2tOmWjUzXfAZYPNZBTVS9x
PpTU0AG5+euktCDgqJYXBaga5XjQ+sF1XrsGMn2J2tcrnOseO9ADjfZ7RVm/
Ml/MBKPSiKOM6pPk789Aghs+5E2PDHreT+ZVKQFtz3MTmj9GlrSuRxF9qoeF
7n/UJrIWFnceA4LE8GKkC941ipAtMl6E5M/hxhrdfmejXbOJ/m9tSF9xYHAZ
PX0Dfjng4aXIeBXCR4q84H+8/TolXlrhppRLBLx7NQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gVdDUzgRtjyGqIopk+qdtRLtcSe6CGN1jnPdYn4B2YFMisDmX/QeSIR2VLXb
EreEPdCK173FbUqwHichqmF/QkGkKLwgmjWKEkQzRKX+X1CtFnAJ8GThu/L1
gyqOejSNLY2T0BrpbSstoonfIv6aE47MfYJpcAxFVuKDEaAru90iuElShmGA
8UI9jcmGvhuz7/k/MU6NxIvm59t7KMbT6HRp/HzmXAPldK4UtJMr8WxCfwl2
kYObH59I/qRoB/LxytGGSiX2SLjsmNWtH1iJ1bPQP+yIDZUy19th/ybvo1iX
5Mxeymdrjo+udb41lUhYSDOYgYbWnLSMpp1ORyIdiA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WLH3gzD/n0m/r3miP9Y4HAuCKg3IAgGV67lkjAphxg+w1ynB/GvEtrvWlYma
9LXxn1RXQO1X4yIvxVQ2gvVCYObbVzgmyDkg54qmQzay9oCcR22Uqu3C1LNx
sfMlw1XmK9aaC/CeXlmNh7Gm5I3Yx7eoGErTr2LD0RohP5ycos9pJt5rm7z1
rQggXE7Hg8Buhgy5ujCH5M/2XKPGcp6qFi2wXJeErVE9sBekPXUgSOJ8xaeI
8iO2mifquNQCSXFr3Os1lIqswHbGJ+3X+qgXWcl5AzF9JSMBmjMvRSvs3RYR
0K64Q/Km49qDGSyWZjUcjl8marmbJI53zq/BvIgaRQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Z8Y/gseR5j5BH9LfQiNpT79/vcZngkeThlrDMh73ZvtldpDSN4yZhi92bvTq
xPVCKJoPYLRc/Jn9MnGps8rpFELuLR7T2aqlVWVJI+sjl4qCf5t2TtCGrJKs
YLia6DP4OTB4pEpcDnE3xAoLC+7VSC1uT6LY2Ys9HmTYokx0E98=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
lG/KTjhjrP5Gwh1BUvJdzy7rDCqrNF6ERn45BijsdgCCt9aFr+tNKMYvRS8d
nVc+LpMdGbciciS2L9C2cdNilpe7Q2cF/m+zA04Wpqp761E/EDjGjdliYrq5
9q8P34vtx39NI59w2Q2blIwX21eyMz3eYNLgujeGakiQsj8hEqZRrDsgEk/r
a0CWg35of4xNEvjpDPm76TdALPoxyp+44rIaOCW+NP8PP5c0mIYClS3g3Pay
23PbTwuhEFhf1rxpvYXuwUIDpk7aRjg9twpmIAhjPh1A2uQGasGSDNbyAX+t
zrCqFjk94NKuUeTDZto2umv7NvQcPcE9opD0OzDmOeE6xQFF5PtyAZbpR0Jh
c5BJB0pb37EP9E4WxS2bKpIZtlYuhvS5RNH3rLWGXErMcGTFeQ4BvdFHzPfJ
Rc+KYt8CLCeAOzGg6XrzeUwImHRgxMzGtMxCyXC0TJQ7l/afTE/MNvyEkM9X
eAq+Bw1qBgv0Fs5KQu6689bh15molUhD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oUSXCw1Wws6rCz8uoh4NWlJFB7jmtRc/M+DTE7/AFzfB1+fs8SdQ9w3SV65v
0Q5Y6zDVv5pITJ2EKoAMcWPvSw0stJpEmR5xvwJuFOBwcOTANoEfAKBgYqak
hwAyJa/E5hZ+1Q5jH+aYZVsaQlzmFMZ63Q8phIoYuZ18QGGsRMs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B46L+vJeDnLRD0diOU9+0CcJ+m4cYNS9tsfoUvKSvF0txk4fw4b7JgtgTysB
didOABNdlXIJtHT84LHKfAdu/bYcWhE3uNXX03tS8TvR0lP77x5Yp6+midur
zBOsf16+PFcQ0+3OdS6vipZeiOkwHTTIwmW/CzqSKC0naVMVT60=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8736)
`pragma protect data_block
fjfwNgnwxlx51766F/NW9HpKdUC7Vp/12lPUE1z+LNdLxKtYMywWQo+xHsXs
Eq6Bds+rxxWXnLZCpCObyVPLStzsM7i+j9U0SUACmVMqNj1VndukvnUWGehp
Xo3u2OwBYt8FlO1JYx7fVQ+c8/59eE+EZQ7w22rA+rK7j2r5H2lUEK8HlRS4
sTB6Y8z9872j53ZVzvx5U2fiMJDwaW9AIQfLpYtkFCy4dT7lcl2iAvimFPkG
XygBXHarYkP9IbRVDbbHLMj1qYXP9Bqwq/f/PbrSx2gZ+d1KVnZYuwAIGMqK
CRjeCia5+PQ6W+4DnSyY7zzi7EETLbIJUxW5ecpywrgAYI/HNqwwG1sxyZ7A
Qm/2LMWrA0i20eJHDYiQe2O5P+mVfGKCIeDZgBXP8RQKxjsLk59UMXAGQMe0
gDBxo6N3NzrB+HaqEw50j0kYHriK+8CTJR8jqfO8akKbHUKKMf+JlJf36CLp
YoNe42EBMd9dCXtcTSQVI+7hqAL2Vix9NsFdeIGgZd2ocIPGIG6PqgWu//uF
2saUup1gcZlmMIGJo1+CYMp2KU3mh9vDbJsdRhLeFF5lD8q3SNNONHqbMTWd
8kRPS6P4L/a1r8TYSeb85PtJk9q8bBwTaJXBzm7WTQBteWk2kRtCwN7wHKac
uP0dD0T7MZQc3zW2kLVy1+qIrWuEoUvFCO0Xlm5LHOBogtUyUgKvki59yXFi
2rBuiz9nROaz5VQWTk4iDZLqU8Qx1tBcSfMARQPu7vbDp+6th3NiczT8C1Et
d8uTaAEKIiEfC3fLO2TYgeU50XUsvakJbawAUVIbjcUJjL/CgNMrwCpJ5e0Y
Mrx5hR5RCF+IqAwEWPyv2AU1tNV44hTWmZK2ytXf5eJ5XS7+nHnMYB7bSn+1
fpb6Ct0ESFRtNnU6QWoX8B1cVsjk1jEbkPShaY3nAsQuGnvWFylh9y3fr4y/
NQ31QCaiY6PLHcqrZF3ksTwOgDe+4F1XqwJ4qv6qvBEnwu1ZwdZChJaCYdQl
7uDfAfgf/dv621jtOouxRyEnEMxTo7mAN8b0zRWBTV0TzC2e8YCh53yyQZnh
ANoy/np8k075NIzEKDmmWy4xPJs74WF3MjGNv3n7FAE8iJ66Sf5sb9y9SeBK
STOT4afW5WKZJngYmuyLQbrjsar5r11MGKI9WcE8Ia5wMmMe3jZkx1h5Xc2P
7MfmrQYVhVI7xSMsjAtEu/xoJxUH0uzU/7LstQ6yxgrQdgbZ7INjVaXBpEx5
GYXx/xop92K4Ze1C4jyP+7Jni0QJ3XIonUdp3csBvdd3dRiS3UxbSmQj8XJJ
FIhsydbnGvzEo0FmC3cjurw+k+bzKLzsV4gkGwFMtFMNdlsdE/AnvgEQ+ac+
iX0Vsl1oIIJWF46tSs5yaD4T+PTc+KZDvZ/DRxKWEctkG53VXygUlapCU/5i
AhOKnr+pE16i2Jk2LSoj0+4Dz1jSwTrX9E5sKr6J/DzjBWciP4vkt8DJPe0r
NqFjmkLrPq2/XeUa5/RQijDVabkQOL+Fo1/LseKPwO7JmpIjyqp7ze4G9jGQ
VmZgPSJgz4ddK/UbQg2RGm0X+ZGlex5IJQlyYwDyUj0zrExhU3PhNsivze9b
GlMJHk5TZoOKFeKpy2/U3w9C04i3EIl0fytThRiJiRozqowrVsY87K6t+lKG
ufncWglfrQJ3JOGXOo1Q80EJSxCgUwfOvafVC6dGAPMAY9vgJr6Wdi46XwLF
d1kfCr/DXf/aTunv1oalNNHUv2GSBRCXJ/DHq/CW3sW9HdPXaENMRobMUtmK
D8IsumHdf80mipg5VaibnI3X8FjMRdTFFqEOh8hJyAAYBwj10bS6+4UC5/B1
IsfKH+utgwbPBmylBlbsTmLRZ1zABUhck61NcNmU65ZPuXbfqLn7f9WPBA2T
nNSAgg7Z4LAJxpRr1s4etqBYlhOZLhCL0Dsqq36ia6oRD4GgW+MlArGVUuhx
SGNVNLQfYEMFcMp5klE4RYjMchLkuAPzwWk6LKCdGsWmpS9f/cwDmCzXfrE+
CE8VyuS2d3TuNAi5hu6coZYqklphXzDyl+K+i6E6DaJYhprhxRb0p+L2KMsz
GW4o9kQyNkoueOjvNLdX46Vpz/r7QmtMUvxeXIIx6TzUQ6Vz/aynkocmqQf6
07I39M8QKHp41bsi39dSM4D7h/6v4wkfEr0ReweuBiuTiVHc4c4+0EoH7ZdD
LOzQSROAnRCeQuq1q4jWPszWjccUis0+d9Lzr327qYDG8EZFvWe/KakArrpa
bPP5U5hRFjc8fGSVoMiarpo3RacRlDhBWAa/zgNPnwBZDDyDrW52XBHByXrP
8GSFA2FkXkxC5SVGo638AQl912cqb4wMl2yT1vQbtyFjoHZh8BOUjC2ZrhYd
jCtaNT5qcBYOTCG/FYt5d8bkEGIpmX14tOCXa/Uz7llG0n600f2idnFuIf9H
tdNWJgoTe+7nmV1pflvICRAzAMtM8tsh7QYvb8VYti/ZszbcYo78EssCInc9
w0MFL5KZtg6zzlWcY8GAYX3sRlaYEtPB61A6V0x6ImxWnWNFCSMhkPMwpSIR
UBS/HpudccGBiC8uFsB4+j+bZ3WX60H9EBNartn8UoOHdKabnXa6NrzFeVvq
E1+E+KmngaeuTti4uWG4PKjDz0aeSbbGV9aXvCVyQWw7CIKSJMuBTKUCeGLU
NRGEZadqKkwlkIIVB3UA4Dzz5Jlt6zHmmME/Wj87DfwOcRBYAcKgUBpTYO1n
2yas0D4B5YkbNjlelCoSTfLAzH328ooMF8WT9Gmf2wE6TEHMOuhW7Zz5OoBF
pu4K7oP1oEVUGzhERVS8pf9CtDUgtVnduCBogr64SCifdB6H431aHbBM+NfB
zHQMexDXhoYcJ71/65yVseUgoK6afNp8tzvkBqEOLx6rAtBnPEhrBs3h0QFc
ODrEdCWhyKqqlyH5zJ+nfyCFd/vlZPbACYUNFddQZxpw1k27yTijziPEvR1s
jAvt/qd0ZlGrpE7JTGTA1K7BDo7tfap+8JwsQF8GIn5xtw5i0fUPQgHuFBVH
5n6t+4X5l8d3/TgQnLGmJLiX+TEOWrhOTIaipZXDiWKSTLpW8YKP+cVv+VZH
0mHqn3Ox6fC07XmQW7exSvvv7kAMxLN6QOQEBN+/fDQHcMMhF4YkA4M/w0T2
vD+GGGokRo5r+W1ZGNep0uuQvyS50PDR9G7+GExF+LMxlCcNPw3w6nXzDM45
EMNaiu24KdGEsOzwkkEqvcRsxzR2B3njIEZQ2dLmOdx8Wlo3GspxcQZj8gKs
FCa0FDEVehwLuWOC7BSxTTBTVxLQJYizgCuW56AMrcl+l2ArlllSI2PAmv9B
MhB3hOdW/EY4BhlRKx527itPzuQ1zlTZO7LjgkfbW+VnQclYRo8PcK0Mb3gt
nlZaaCP3zSQcbUyogP/ald3BsPPOiLtvmSU10dJkxlOUbu/DeaDNHRtNH0ej
7a3SRmAhSsdTM21hHo9eDu7lhGv3fGG14wBYOncCkooKKab6pAegeuCJGKrf
aWF7LMVev//Tmcv0l5Ci+4dzMjIyKQ7o3C3BXGB9u/uiesfZvFp8KhEnxlBi
Im/I9fAG/zOL8B+h7eVJvLO3QFwnHBtMH9IqekDd7sKbsRd+P2C/LswNEnMW
tOJCTGYRt+kFyF2fQAfzHZSVT0c0eOv6cIigYhuwLrGbp7t9xuoSVPdh2Rzq
/7lJ+gYQ172eqLoR8g4rxAlrKgtpPamFBpLxtKp/tgUhnZE/7586vqA2iLuW
Qsfg1bT/zps85IVb/gO7BYl/773B3CCbFW+nvm6LbhDwdAuPTFyi9GlXubaU
AHzRssrcruvBWL/UttnLB5tgI5In0GWfZruGUbiK6wbnCO/pkrUqd51/1kgW
SzOnK+1BahxfqCxjv8UNrM1lGaAkgdBW8/TWUkkKtI+q9cbeXHqRbefShQWD
Mz+2LI2jKkTpqsgqD0WLBDPE6sYpS0lnWhK07iph5OatP/g7lYEYoC915gsm
e/kv6X5RSa2TF6KPoYcqz89Y2cIKp70IwuZNynOncCx5DeTrFlg6/P2IkMPh
ypS/xt5bfQuMqGtK8+EC62ebFPayrfmZbD8EB7j98qN26HsNvXkec3vusNY5
zbIdBdLg78w3ZkqnR3ANDYGtn0tBX7rK+RArQwAKWH5jkoD/QnlnllOM810r
2c3v8BYIrTbSMMJc9WViudT/iuhG7xCBtj8GiugomIGruNUmChsECbfOnn5r
zZZZ7u9pzSNib8AOzej2O64AIyJ9tTgHDkwTgMchlOjQLK34+EMveUdSBoFy
Le+X9gfuZQyCFw/tPAO36qYh67vtirwNGQYaAMUb55jJJ8g7TYwQe365/iFz
PH+jJooNmEddg9b5QlBnq+Ad06TtXmYjTRfyJz0JiLDmmJEsBSXbKb5zQoQ9
p13rfgtxPnqIxOOPF6x5HDTk1yuWDUg57gSqTkq/Be4qcC6JiCfD3uUGLwtY
ZBbGWioEWlf0idEbv14CvMe9p16fFnOKsRVsaTzqTysJaGzRLouYIh4EBPMJ
3Kn4fxAj452Je/WiLv/lFmDbFCu5KUZXhPGgfOYraLKot3UqcdgNS/NYcWgN
yp0l1gmAtjG/6Dmusnlb8JuafTNczmlqDd53sqgiJIQ7i/21MjTKN0LlNYqi
TOa3EtHSrajOB/Zd1KvFCfaE+FeU5xKtxnUnE4RVY/c+IDBn0iPB6GIX1f8n
iHlY7k3DBDH+ei5QctgiJ++HKUeR4dyafoylCsQ94BsmdnKplKSEXLs/JdAc
9F+G573FINxUddqo4KIHQb8+HK38RmpVUO83Q+7mRG3qwr+yvRG0ofs7T5hZ
gOztEGGrzwN9kIYEPiUdCNDextwunnz6keCW1egmuuAoUKg/SMwiKskpVRQz
QbJMcMDDBZ/c0c1gUwt1RIUKudhZ7Fsg2X8CC2VYIK6uosUlQsflrkCogAjk
l2wn343Ih8xGoTvH8+n/2r+eCTI5CgEzjlz330n8nfkUgTqROZZs9fvX8Uh3
gaRbTbeXMm3a9gPZsfMKZcx6OR21utAi6yJaQR7NPp4J4x9o9r+jjIMfgFdx
KevMw3hqWues2vyFvSIhaD+EBAa2cFzeegRCRP8NFEsF6GzzIlCyjhtZ31JC
q33Fs1bQM8YshBRsbyElQmpWfNEExUfJKawmPGMyeRjnRmzfJf+wUcdlVLVz
MVKLbr0r9cM5yjsxRqZcPP5SFRFCd7QksT/x+dAh91NdvAG0Pje3OcUPzVm1
v01AF2qhKqyMfC0sdIwPEiajJQZkb6W5jGGGN9lqUxFHP264v3Whn/O3xVhE
1UkNIQoV93vjRIjt8XysvYOP/4KcfwtSnQl9+Le5ZVYoryn8nnXIA3mte+kS
HbkbnooVltR3dNb1GLMMdC7aAst8+1CFvpc8/M+kUJYC++Y95fgrq8btXogI
vYTfT4j08LwGrKjizXQDtU6MugBvu1xFKn7Cx5rkAaIlJUyXXHWF9uI3Ydpu
Aemi+VEf9tW4nZ5+FnAA6DFpqHv8+hzzjzAJWv0aQB3UZ4eUiX+FBl6/qt4r
g53nibVeaGDNpQav3mduqQki/lM+mrMabYURiAY8USy3tFpveLWORl3TZ2y1
Pp4HawtZLvK6kk2aI9Q9sN+yomZM0rO6nvAJl1QfuS83jF7D2nu3szYwQkc3
evNkKSVhsirrmwk0lhueJQ15SLhh8nZKoB6jRsVpElHDZX7dGCy5L+5dCPz0
FLUggYaPlCEZRfJgfEVG+OWtvfecsZQ0NyQ/41kw40ak03afet+IJdNKuSEY
aCAvK5Yaw/IPdwUWD9ITYQx/VJjUBRucq2JckF3FKxbK4AEzjcV4epCy/MaG
L31wtLqFLtRsarKnkwrhtgXtLJxB8BKpi1kvE+oZxtWVtixOlWt3xXVeuk48
PLmnkrMgDAe7ORMNW6X+UlwS7Welk1q2lMVVP3HRNKnZ/PKqJ3YpkftlniCq
hxMjhjfcFP5RdscR6rsxNAcRXL+4VEv2Nmugflc36jjwk0X91YHty69If6En
wRlXwHy329zy6Sz5MOTvB2kGj4nPrSeUJiR0oEP6iEIleL7aKZ8khfYZ0MUW
yeLV279fUBuTzETrJVEQUORCykZ0yaeLLif3C1Yl3jqIWdg21xUnl7Xpxe14
cMoK0TsTZ98DdBvCznAiLG9+WadUJ0ypIat4KWV7x04JdZWTWP80O4rdXAms
2dB/Oh+NDqiHRaAgy/mYUd6GsOH1HcUXqkLg5uLh9iils+fPIESt8ZKnXjvc
KRaXD97kBfHuU5p6ZDnnwWO0qGG+B1OsT+NRtB1vFZ4GWCFm5klBy557oWEm
xohVMFJw07wCWF/s19zTAzLGKrbNQlyhdBCFp8eLm2TsGg2obmGSBMU7ziaq
NIk9UDfBUPpni/8SiYTpLz1/hZZnTzlRq7UVQVSpFUzFF58WQEge1OGqRtM/
mlKmv+N4Tx+JWWChCbSPzTtYe5BTuUWgHadxzOlvNNZPzdQPYNWksivd4Bfp
6CTS8hCBvXAi7gfzsRBR8ADCAQboQoGZzSI57xm7eLVUSkVH5KAZ3NSY+obt
OKOvwElWjEkxV+j6U076moxjMVKirx8QHyK7uMI+XTQrVkrT539ko3lXMWaZ
i/iqWKB0bPJY5gwOCiM3fDNdO9qliHJIWB34zg5ZnjTN9SOUlyd/Jxvv9DVp
UdrwJSNmFN+HDF4a4IIy/6kbTGWoO7Hnq5g97ATTqcq6KoIDWO2naEENccLU
Vksd31ipp8ihZtGNFEGn/p8LH328Et8rsqvXCIlvMCQTFegJFE/xKu3W91wS
/SF+5jQ6k2MGOlU77U+jtnCzb9S2L1kIo2dYF22wG1wRZuERJg8jshXdgFhX
nB7uUX7CRX3UnQLC8/UAR8nZxLMRAQEaztnKuXCXeTcz5znIWshjAWiYbJEY
444x2aorQ5Q6IQYlsiMjqfX+dM4eEl79x46lKTGyCbRAq+D2cdp5Nc1T3wE6
Ej+gTWY2UslwG/kiX2RtMCwp40znmxgrnOP0bVqBt7uEmt1a3HFsJAASAQNS
U0w6RkOi9RAR9fiyumkE3zPiX+ljXNQeKaa1sNVFPMnNwdZIEFlS5gWyw/V2
vwQ2eGJDgSf1ts7518LDzaBVmPoOcUKl0q1wPUgPT6Al06Nst7GTRVp3/+57
9VQfLIW/VFtzlE+qsEvQMwN6JaqbcGFxaxbWU2zHanldcp0S3+rekbJMBGai
83O6tHjYJAHxLGWonV6OduSY/bfCPGZIERpmSPpv6WPnngAhR8EEaRtqMK/B
jMMV/8WNlgrmWeg6n6PTji9bWibXG2/X5u+KnbJcCBsMFXzU5Hm0g5zUXxdM
20WB3vgSpzq/A6Ow/NQzsQDNKTnp1RjO5HRI4dxbNkCEcT7JLJsfeB6uM1sn
kYar3LkP8OdFicE1zjAyr0YOiT79xVBiQEUlBppwMdNbTk52ZC06MG6Z6zqx
JHok69loz8GT7Zy/PoPKql1l1JOcVturAZEv1KO63DiNs59MhseQl968pRJf
W+p8osL39oKrKzBNunxshaFsYy5sd/Pp+TEcNSMWz01KDLxuar3QodirGZnO
db5v8iokYEirQH04LYnaptqZ8X9OX86/2p///NoXaZ7ablTUOfJm6uqZjLT4
b54K+qGiqOiuU+9XfuWxK7CjRZ9+aHRxzwwjIt9nyKLy6Wyq8B0qHXAhDj87
V1NjKEyP0NkOyj4InLfIW2Gsy2+QIyDqlxaCU22rqom2Z9ce/qO5DZhO0svO
sRoKT006Xg+QNUG+w979XAMnJI320mv44waZXjEKCTDsW/Qvs6o5UJ1V9O8O
U9/a+iHXIFmr1njAf6wx+ALqU3WwskrEVi7qShM1cKks/SkA2uDF1HSIH5LW
zN6yvreIxU1hMi9exj0ebhvQ0qxTKNj55/zaxgTF9uYCs7NB1+qBhlfnXy7K
RNt13AF391sUTZ8aGtfvZPY5WteD9U/sU9kT3ITYukKc4ATEAB2f0JpcBukI
m+9BXz02vSTs9lfiJ3tgxUizhzmu3gr1WIV/+GOzy1yQC9Br8A8ZUfLO/BiN
XAlLUg1tgViIfKKbw4+QzeN/nMvLSe+7NZJ2uigVDdxnxsi8urclbenR4W+d
zIPNcz7sUBbzjJILLqQljI4vaqBITv1IekczSk7HjHeRTXJNNsyxtH+5I1X1
jUqlBxvK/0phOSWpwojC8YcTmR094iwHJXwbWtOr1EhPXda8aHkRWH17ugl4
Vk3pN+zZwg52OrEgG/qzEzKSA/HuzkbUocMmW0Mqpej1i+lkP1rFQo2fNtEk
Y9zoPpfVIGcqqXL4HAN03ok1HS+cih0LUR9uGXaRb1ptOmisc4wERmCmTA9R
4GLzFA42vfWSZ+AkUmQQHUTX1SXOk7c1oo/Sh4OJGpXDLCLKGhKiIFgJsiDT
onwnWRyGtCWtpTNGBaJvVMl/hUu9PzufUUlrTeP2yYRni4NUKliK6aOJu11n
uFheQOkv+taMPbqkjAFxt8cUXJKmjh4RliB5vnrgekCnNrLB+tFzHGoSMyFZ
P79poqBI36KG5Q1WGL5B81BYbbiYZ4Y0v2gif+loVnReuE/BpIuO6jEWpgkl
kud5KVN1aybhwU9a1XRdUQPoYHZwgE5Yzmzz7xcJtqqf/Wh5ymn1gXYRcfze
aCR5Xx2iEAe2CIrk1xXkUL7R+ATjO+FT70xGoxGDWZxtXlR2hDOoQtOvNl3E
AMEMC/I07UEY4afRXXMxF9V2/JooNdauF4REpnmjKGwsoSuRk45T+PL7jCCj
YpbiuezvdbMonDOauVO2nuYOGc5HuZlX/cAPSVtjObcUHjwPgTnndh2TqWs1
MUh+6ruHyt3isQ7mnATcXB6DCnsDtks61VhUPU2qF2/Htp0UTsOY6h4JXFpy
gGlyAAj+eunP82ol0th7KeehWTIWGp4uFGhSSXr7os5fT41pDC9jsAi77f+7
zXLlbUS/xbUmhVq5Fepb7aHmiOJOYGeZ1hVwk9TzmVMmYDKqdSsTYSa2Lcss
nJf9U+27vzvv63/AJO5c448xcU174ZOExKOxPDi7Gh+Yfr42z+neIspS2+c0
WeF1YSBHixMizDlB0YVKPjBSIV1xFB9B2DV4GVqq97pP3G/pHYwRjP2XzT1b
zsOUaqqbN7q8Rz09hoOw9YiAuNrGTE+oZ0Ot92DemXneF7C/zQxPvbmJJMzU
KVqSXjZLnpU1Oz0UeJD4O8V2tlwqaMPMYydHeX8O4XJADqSc4ODZMqGf6RPr
aL8kAiHr9Z6QtOelgI1SsRYDMikqFC2oLlT2bS7xpENh8lDJz1UmPBVCFIxJ
jRx/ctZKMXFFeQzxChnF8THv08cbb/hH3WEPVLa+S9TXRAJYkKyxSNmae6bD
LShoREZMi163pGsfOLCM7WHMiSUVnO1YyfVJufa/sMkzIScMs5yMyTZzOcoL
CvdQ5g47N/oLuXzJ2tMILJ1RnShXoyevqeE0I4IgR+gCUOYcH5Jt22kn/0NV
U4UcgyEtbsiu8vvqgDyUhLoCjdG1H10OsX1/HgNPFaprFheV7VE4YvOgjqef
GiCoQSFPfWGcNEQQMzurqdjTIw5gHNKWdYTHY6B2UGfqZ4VNaGwo5I9lcUew
9jDNpTuP6eVUTLax7XI9ChNQpvgfsmdmVsMCIkv/r3kbL/gfS11S+zwfAKlT
RBJ7txV259n7uEwpJU9SHmLvm+xymSTjb4a4Eo7HpdarJBQ1psbmO/S3WUyX
8iWQXdqntfCxnMv9GH3LwfF6bxcsJQ2ddfqHpWyX6LLa56Lcmebok0WTMten
SJZBXy+SPQ3Nhgi0H7INLv+0R46ZOdzwIcw8TeSz7cUy88NwkKvU/Vty1+LC
cSR4eVmthTzFgfudgcaPgV/LG3Lov8RRC07SpVaARriZHvlz85v8OsQ7+r++
+XS97hkED9yMTa1Y1ygXt9Omkt8sR0YTPS6iMEvN+QI+TiKr7qBV3IY9LZsN
aoaYY+/LuSTiCpzwPu6kWFNn8V7P8pey43ounjf+175Im7Rw0QFyDF6tqVdq
gBSXyevVIoMVj6Eezk9O+9GETVvf15SAc8ll5YR6gUdZ483/IwSvDC4kr4mp
1kTLMbDkBZm4JXoWhjwys1iFJ/hpnO1dlkXK28xT8mJuysE5YeLQ7SJiT6pI
jDgJ+YlYlHeBEMY0o5ndvB150naHTM7GVSLsRKeMy2XKyl+W23/2iTIYxUev
jeq1f32HUTtr4E0BXglEje7A+BfiUyLKLw724eLJm0vLuxEBkW0ZyyN+g+H9
FAADA+JCwkAYrPcGhcZtBeee/Bk76D/vFymOP0Q9t280rifSycPAovk1SOK/
szxs8nUHUGUiXGG7xifvkni4ocyREIvir/oh8G8nI7fWOLLHdv4LPg+7NHXT
vifEdUscL0FCcW0jkZM2DCoxuRxUwZXXTeqqqKPh3kd7PyP0bGpjkXC+ad33
V/JaC5yDDDyTV1aSe+23HsQ95OOOW9D4d7HjcJmDMsmIpAcAuCP1+T3sxSJl
K2NjexfM4bjMckG78WFXmojR7XGIXMPQ4EpcGbHJCOKjnjub+af+JYjFJVOv
SGGXf/HQcjyuewm8gk+dwGkfZtzYDkOsK9hx2hh6AK3Z4FhMaXuqySToGf8v
GKdZhEc4Th905K5bx6Q7beBhSD5S81kTtyl3LblIQK96gjvW1SrwkBZINshF
M3kzEMGUIXxTMItmPWLvbKIKiuv6PwFduPHUUhA8Nbdy0hlMjbm6QgSmGHR5
VknivcAuyup6sx2aOtcMq0q9aGg98e+VcWqGhtgtelMWjHxyv1RIiPhhyS5q
gKoqbXXnlFVuCVpRykGvZ7iQ2ddRbeajY0e+Ga2VJ8LYsK/zFRhQClHZxheW
UvizpIJO7KS5AucnpwyEd3ErA6raaJ4xj1bnHdx2NpkypvC16kk232BYLQP7
ZVvolFuRiaj7dGHJO0IqKLjlaUOFpJRmJp0Y1GmZuFj5nnyDI9c5AtCl1MKP
WWn/97/LtlMyu/2Ns4KP4CTHFzQT/R4SYZN32IRII3zpsvPYy6w8mtKgglWg
+cdzdGxmya8V5j6RjW73GsJilQl77J1m7KQDyBz+mtLxhI2CT3k8s1YGQIrg
hp3VzfnPWf2ICGmy7DyDHdPS+iMOXaTchuq+LI0GQM2+GtCpomSUdreopqsU
rL7yE8q71ICyiLHj8pc+z/QaGp7CMKAAWkdozhdrzf0cWi9beC6KqkMNaV+7
oazjiuaHb26XCUszqkWQEmjzBGb1YspnzxoHDa6aIIOIQ3WgrjNJDw+ZFDEO
7ihrtIKjG2uhjkYmwXU50flrnzSpwUHmWSRFHvkzKnPXjjTjCDvaE2q87jZA
z8BVVwNRR8LVnFrLh33vnQ3lNGdXoCdPMLuGYJHNVaBngDeC5BTLh5UrQABV
74r7lWWuifhgvadwQRKMd29Yw5SBf6d2DfYoOSRijMX9gkQ6rRv4p+yJJug2
TzVcvngTnyxDUkGUiUhC/Z789Z6fT0J+TMEGHEydDzh+n5ont/h2aq9zaezk
IFeDIZQ2GnuRCeL8b9bA2Q79FykgpOrAmqBSKkDqUHSuNCXdU2PVa4pqycXI
c/yMJP8X

`pragma protect end_protected
