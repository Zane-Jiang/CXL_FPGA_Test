// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NrSYWthCSf5jA01PQv24mIbG6zpcK2/ykZHWZFAJtrcfmqRjfI8wsp+KHtxz
WW1lgyHr3npkm0wWQmxKkPt8EgSPY19h0WgA33tqVOcYDN8adQ+SYzCyKi/I
kHxQ/bsl6wodWnrQQgRFngSXsR8UrNHMj8f9vNV501lUEtdOBU1nBH1dbpVL
kLChtvELeEnAC3THeqG6j7l2m6ohI4PVVYsdxcMOOhptvKAIOitL6feG0Fc+
gcxHfhGIZ+QAN1SjhZkU7BNgYNQHFvx3bPGrLWJ+Yy33MYUAVKCe10tyHYGL
p5vvar+5pij1LXWQfCYJUX3B0fEWB+Zf2QKvBjOH4w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BYmXcyE7ccEEKAafkNvLKFQ4xDLuxLLDG8MRIU2t1J5baIjXM2erHnrjnm6n
GIypMBba2yD45uQvcISgZ8aqgu1GMJQwJeIOkLiQd+FgV7/pLKq6xeEKkXn+
iYT4NpTD4YBUhYoz02D5M2qjXlcfaAm9f3A2ZbBCyfN/A/7koMKVzLIJ/4Nk
4r7x6Ca+mA4i+vqXRFx003+mWmZhCRHU/KoIQqCjpbeHGnZ0l+s3OiWKWZ54
FrHIphKMtkBcvBptB3QjDCnGGwKEB6ONt7gE5XwPqfh0bUNczbzGe6YXkklk
nj5MTo7mvpKvuIQpe3qR6Ep2k/11FhfrVT3lToaw4g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AtFigGStPdHwsTWdBjgnctTIX/a64y69HT2OXdZMoQHDYeRx8EJIYY1M0ruq
x0figp1pB4siIvc7s6i0WvWkvvY9q+XWh7eG5gJjv2LyzFtmuq31foh4dAg9
jEXiyLddjO8nBYpQId8+0FhXJpvdz47o9gnGS3+1QTbM8ucKm1Td9fBjngc+
+xTlg3bSnbzICmTeoZo76GGUweTUED9SMmp9ppJqgU+Wvx3B6bKuADcndOVp
mlT//LFgnMOfD57M69KAwbL91gU+xDDGhdeRcVb4sDPz4ZmSkPkuu/tw8LWh
O53C7HRrjQpStEfIYtr8mSKHWV7Qmc+quZt4gfKHDA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
We8ig8LeUf8bc4sxZYuPYZLwcqb3cmuhtP7mLHkawo3MwcYBKhTJOen/R/Ig
Qrqh6Dbab0qhvk0WyVjyTmvpIyDh+r38oyHKmknTxXFpNmhLz5NHWHxrO+ag
5lmtzo2Cy0aNg4FP+Wo9/vK2IgOUkl9HbqA6qO4FLhMQsJFGV8M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
M1v4SU8L8n4wPn2VPomkz8YJvVtniY4CdB9GkAyC8cgvJyI7QVMJn6E+wwMq
wpkYmsWr4iKtuSXwaNx5kyu7Wdo0z3tvyfuanjxoxODjddlD1+0qq/H8IF8m
VzhSGn1DoT32WUxy9btEghsRcvEiPGU8bW8S2x//wjcF/O63tYDatmOE5CT/
iQibsXRSld+R8L1K0yUw2CIHslNUJizQIechh0zSPjur40FRW1KWkn4knxVl
h1+3YeR4MXYnO7BaD4cRXQOxTP70XlJcrZlPVOUS04rQXXQgkDvrYLRfXU0Z
T6tYOqfH4XfwVeG4kR6PanJpypXOuK2CpgoNV0pO502VITirHbNjroNyqIKk
wTiqaQtWgb5W8bhHV10l9SsRwzkHs8RZeiKYUxY5QDYNEuuGUxdLxiEc3YN6
cBnRz/ydHubzpXYKRf4nzLndgULbXmdv3HFmssNhIZkXryIpTwpAtt7WfvC6
AzKPPk6UDQEV0rtiMSmWr72uG5aF4Jn5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KSrHA5i6cIBva5vqcjS9WoCiZxCTgGD8OySytHr71B81E/OoGbqbBIGDINmn
NIz1ZxMF1X+TtoallVuA6V7K7yx8EMdO28xtnCHaia6QjJTxjmWAVnM+3/a5
Xk6NhVLR3iu0rPiIc8q5o84cY61oB/lt4NVGqMjoXxVQDLuyKBY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Gh5dHbje2mQR3S5qyX6nMmQpSY75twmGfdQPlWLU12eT508gQL6G0WHxCr+f
9DC4R14E1e35AgZR7PSxZntyTJJnqub5mDgBWIIXzhjwELONU1L+gLiwxWVP
xbTBLmhtf82TYr62usD7UwF+LE7VD5gPJG41IQPRIYkmCiH7bQw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1008)
`pragma protect data_block
+dwYOM8jQEnIrZ2ulJwweNtiH6czIo05DSms/dX5PvrILiapmPlLGT/M2ei6
dW+qFZoddI6PpNTSj+Dw2SDnm7/ioERyrJE4VT1p4Zy6oEMKuyhkMR+uRQUK
NmVrFbFqqaSHWG0B5uIieW9eQocqP18SeSUbmd+m3Zkm5flil+9unEYS12Zc
SYfw3EqEUeGo0HtDhf/2EPBRu/CfTLawCnkmDaK5W49Kq9grQfJl0wVehZsH
FxGS1UUapm2I8+8ms+8sA/YRt8RewHB/6O006iLRUTdIxGHVxYx1NrC97bDL
61HSdGXtTbU6nDkPcgOeSRFZZzfoAx6FPAzOVjCjrVZpCkmzLzTyPmzEoJA3
q99ZotMBSDmFL1GAUJ0NcdRdELgKEnBWq6I7csTCzGzCGCQY3fcDeRIVAmvN
y0u2ZZgGsdHH/hYKDnI4DlpzQAIrQdvi2OBMLXFxlNfTnklAB4snFWZDQegn
Jjpvyo1QeYCdOgT96zUxONbTvM5UqRNzFVqKw9fGvw47fZGdCMa2Y3OXiikv
oR1Dn3e/GJ6RHzCbsQ+wJH+hJ2PTtgi1vw5al0ownD8Q0zeXKTk6PVPxihG0
YegUBFnpPdFXfVDw/9XoCc5cAjvgx49Ru31rVSLK5QhmrAmbZCEM14j2GEV2
WRuVCGWQvgHBiBRj5OCr1bHmATVjG6gTOkdOhgxfKvlYOvN9fJXTUjhtmgTU
nleVodMr1MPmuA8HPnfouIaO4UzAf4iuYI8Qyf2Kx0sBs6EbSrntDzkJrK/w
nBxwa8DGE1ENzCThJ2S9DMJJPI6sld+HShN9LJVGFb52KyOTZd03Kg0xkk/7
dFkzMI3DDi/wD2hHq3X3TNzgrFmn+SN70u/hTOHDn5Sa6DqKYjupP6FjStdL
GZtR+JolCebe/RZQDmSxjyAWIRIS3W+Cr0OyCrFa9dl6wl8sk5RoqlFkHaZ4
fkIMuLdno/UgTPrwBji9PWuXexp0U9Hmj/ARHeXuM1JF640hD49oi+DuCFX+
QDdC3svdr54XwZBTjkqFRuU6n8xABj43QMKcZpArrA+wXMs1tqm4aWlEzc/y
L1QfPi9KP9s+g2gSCB45Zu4M5RANk2KscjRtR45PilJJR93Np4xC3itnWrmj
6S/uYX3UlttPnYyKaR/VDdU+pTz7xpccNEWe1pB+WN7J7ufmkWP3rbER9JLU
mXCJc6ljxQgmFCits21t6rQYPqosQ7x4lEiJ+EdloWHh0eTUYlxiZALcpBac
ALd5QrKT9AuOlfP8cXQTaCZXgT6wow4DgWHi63qTpaMKGCOeqt1p2Gp8IEJT
lMhllDNbiEEL5O7XvAQu7Uhf

`pragma protect end_protected
