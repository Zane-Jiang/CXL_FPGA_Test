// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jpqw2ObzsvYiWrb0fCkdGeqDdoJ5eXMqD5gYtTIKb+2q8cU8cnoOndYmhb+q
JQr72KJTobuVLTBExBy8lkV7WB2NBWcKNe9fdXr0uwsoSfhskoNiiQbN0s6o
SOXdTx+lRF9LY1M/A1V6A0djx5pkxNvJzUKrzm7O1p79XOyoCvPdHcVu4SZ2
jH/Y/t14iTqQKXDbp1ihFXJOguZkVsnI8rXQTQhJXAcMhSN+cJ8KZyCEft2K
IeFh4FvDU/pGFzhRHKgsM0jhq8Gi0uXQwV+ozdM9xOWe4XSWemn0BE24HSfG
JllrohxZuDlO1KS1WH0w1qbuWE92l95WoEtTuaRsXA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WgLqb77mQc2xU3b8mElg4beH9UQr3kziPQBUZPWF8Axt989QX3VfS5z5wDzh
2311uzmrqTSO80aVMX4bhDKlAozjiy9A5ZrmsFMM4idv1J8Yv97WrnyhTlZX
3dDsLTHtVYw8nRVufq2kt5E7sDX9BQnOUmZgHYL1Bwji3QJQGzbLLc2HZTnD
xDpi3AtEFf3biiuJ0hyAGrx+TvoAcS5v7SP/BIL7HMnAItF438RzJkdqM4dw
aG7LgdtJq1QxrRICCQUOyhMiQ4ZrHzsjMnY6ArJIUBt7m2AIEL1sK5+HXI/F
CWUI5eUqC4pGgZWavZqKoiUVKis31xtD9xqKGUD9sg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XQZCq+Zajijcq9BGjyI56mKIuhKB8ylkew9nNQlR7foWN9G7YVbCS+DPqNIu
Zt6HuEX1Gci4poV2uF+nhoHG8YpXWpP8Wc5jsPtSyFfB0E3LRl3JS4I1SpU5
q2++p9aVUq17vYHludtbv+/23c3D1C7RqJPqmr8AYQZHZdRA++E09wBqlc1K
RziiRQuMWqBRpKFyqLNUZlySPNOFcw/HSDocarf84A4Ckhu30QX8M2aNbE+O
bpPTAuvCYlbqP14X7B/aJeZ4pG9XS6C0a450CYWwHtIWHZdaoXHxV0tnB1tp
ohaQ/8cFZNKPOKYzBuzdbA2Cgu1vH7w99r4DPf1G3Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
U7zbzLFoCinwz5fU+jqz4jCi/4Ua9mpI96znBq7SgEcVjX9fUugJFJJCwTcb
nos4rIIXrisqdHTgACD33cth2RULAv/hLjxnIuAtRF7cWtzhRN9IEUaQmJ/D
YLLETToiMC8Z5TgGj8AknRAQ6fYmOphCaHVnBD27DFqcbxGpnlc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GimFhHsN6eHoE1D3xrfzoooNx3WU261rNcAKXPtZHx+8c00/8zUmrZCBWFqL
waOyk0fU5T84l6uw74kfSQqq8D/08pC8q4DMNferaEezhvkpn5XOPmR+Tl8T
8b4xvjnqKOTMhg6zqI8CoxZ7qXboXAUTiwhockVjvMmuaNfRML1j5FgtnQNY
lWv3j/QrrYjwCaELKd/03DulrKpC74j5Q5L1frAbKP4FOB1WkdQ1qOuYjU4k
StKusGPwce4Fu+KZByWZXMSyKseBfv2w3Vujhtk4Egx6lwxnRS5jQBsFNUhd
Di1nn/Apl2P30vVQhkIuxQ+epR+Q9dd0qG86rY5Up8G235nW8mcpDOAoxjum
WZ7CawgWf+kJZ43bgz0cVhIrGaECHYAfEmxVEKxn/Xox/SwhS49q6OHqMOuh
YyrHTXuZ4kLeGMY3In0aFCCEMLQcmALJR8EhBUWEDoRPPD2h2C4pXAFXHvBv
CPSedLjzu+psXdH7pMtgMMPlYM3HQmR1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
b1DeqHi9ztZ7hmNFV0+9gi+ICks6kePin7AV6b9eCTmYd9+oGryD3smbamOO
LSsuD2Jcq7FziInjKZBJELRKnRZjVjDSNYSzxF4QxYIA3ty2WYhlmUoHzgFL
s9JrncHTS0r3N4he0KbHeJ4TYIELT97KUHjUxBcSQoyZPpRd9jI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
c9LT+q24f61QbMssQEvWEHsvN9TnIov9DixdogGQAQsGAOOkWUNENeN8FBFj
bIYiIvPY4ZIFF05xRzFK1OCnivSTrjmoPvJaWsDpnxuT1Dja2BMB0IK1n4au
e7RSZUSxpJ40qa+bAoSWPGEQFOa+iQrGweZ5jbiMS/hdzDhXcs4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7872)
`pragma protect data_block
EAnJ8EFo9KcbHxAO7dSIeDmL3u9pfANWjIrbmbSMyCYQ/fjKyO21zK32w8AW
oAgCp6qXptuy/51Z4GntdaR5mrL7rJmChVdkiHSlN7AJHkJQLkM0ApTBBnV7
qxko/zAcM5+eVgET1aOdNpVWyDA5uvVZmG9wfckJPp0iUyds8YXvDHAa54pc
d24n1U6srZEdiSF/xMNf66BMIKsklWTzsErzsclt0jAoVNwXirwhI3OVVD4r
Z/P5SSS62Jh+swlTBRPlZ5sEVj61hF41pp4JlgoLf0mScJEQ2IxVLeyJvL7e
+KUF8Y80xB3y6f4mPkQ6Xg6Kc3bQFAc+n3ukQQzokiYr/fgfcnhyudBaxIJI
M4FTtyOZ+I4z4aySO6FvI2KuRrjecb1jXZjEE3OKwuA2UZcqy+G3jsupVcL6
hdix7fEU3qtQ3P5VASeYOMdrGx3fUN8P34KSOY9mlgMZfqT2TONGvjp1DJrt
wtEQO9R+MvLPndssuyLnaZuMftrCDKIgw7LzXTOEe+IBbnjE7iDhPMtl7Xgy
RRJhywirMuA3mQQ1hi2ERH7cif7FCYFuj9GG2oYfh3HVuNAEKzMhyXeRgZMj
D6jDdyNT+uQAV8FHB28IZRyhE53FOziNaDUAcC5a9/fuMdSOmJith/0xflTS
c1eckyrgtNPd/cVwwcnyAl10mm8WBllXk8TI01bENz2rI14yoYi/hFgv1dit
NqGQYtg+r/fKs8Jj/SGlcBpgf2pp6ALLNldpiMiKjZqFfsTj+fy7Q68h7z3P
6a4+/y8nVXLMFBNaC3oekvi4+EVCNg1lJyG8Ds7vgtCbQ1hVH60PZyA6BcQH
RGOWDY6Flwx/txFGJa1yv9TnHFfle7O5wUxIgFIuquFNx+GmCeh49jwuP/AF
/BUQ78Cjm84V6h4fPP0XoMhKCysHTKw5iyPigayyxi+k1MmGiO9iiYBbJbev
hFV9hI6yiSRsU1sZ9LjWDscjeFvY7OzUk5IYZS/8MkD4i6dLEP3h6CrGXaLz
gRJH8xHNTW4fvT31W/ELxNnJ9o5jy1CDWVHHfyL8S4+JzEHpK9v58rGPFYfJ
fiMqeBk81Fe+KTlZWWtwhp/8HXmt20wC0IpinMMNK6uJSOl5IbjpELV/O5nY
VFFtFHSM4NLPjn4raPrVJezL1X/9XMc1TVrwo7/cZAU5T3rmjsaivosQ8vyP
LQdNqBxlctCy4Zt5fvBBVsoOBYE2Aiglo8D41IgZpvQpcA2ZWhdESs3cDna0
LopD/aHqwIWY7IztAjNDGRO4EpZY2dVugtToMAtRCqHwTQS1QCZq1Buf6vd5
NWuQTx3T21qw2lZ8Rdiz8eQZ5c6JOdStagFahsGHyrlvqueciyLN0eScu50b
laWPc1LzF2sTKnemf66UNScozbO7y2rz6z1dPcuJzMXvbX7KLofzBo3bDjot
ceAwc4JLC+bIGRhL5b45z9TvlFyTHvHM1Tf+ksTsjpc4gwrtIex3bLcO3MtV
hjZPcXIWRjIbCApRItsgGEqsuD66ZtrAXSUnnrA+RcdeWfp+EjvXOJQXP1sa
ix98u4LQy3M6Ez9HRqR8eXFii2ZXKxSsK/GXSk+SKbabczylvZyvWq2fAda+
ZWAIBqFBTuMGT0zti3oohxCUUXwOmS4LlDqbUyvUxbalTlnVfbaDD8zidwr6
M0jobPz1Y8rIvKpIenf2MotKmiTfkKDCIHjdnRdhW+/NmKwKCO8Lr127hyA5
YHQ/+WFmTcpb37F9kFFCjiSWCVMrZIeBJcP8p0evAp+eDGEIzFdwolBHu7KX
gD2T99Bng0sLzaGKN13YmHd901KgrAxtXefrbvvZEDrirqpWL3zlF6b/H93M
Bzkdu1ug6Z8mjPjS2vanXocr0K36tNnL5vz7FF8IRqSFXjGZSdZXgOZy6WWd
aBpD5tcRakvHdOe5LcrymxWBL0TZGejzq7XXjhxkLLdKwuqtvwl/P2mB/HHU
f+N88BKOSJ4sQefoRlhvT/66ZJyeLgSxGvGPgEXuhS/EH5K8xIhVsiWImpaN
UZ8go01jX+D8KczNAa0EB3SOgheemcWvA4lmDsbK3Juu2Sax2Pg4W6dmRVRv
DHCMqPCc2zvAPCE4bgv7sz9pEGJuBxw25uCHIA7NIb7Vc3opX02MePQSt0V2
CFbW1uhYe2Q9GiESe8LmQBv+T519ZIUTcunnK6gUSJXYl/jsDZwi9bdbivnE
8D+AN7EZJtI3i8RKOmtvcpRJi3s956U60FvWYp7xOqk1iyf2PRIvi9ehKucW
AjGaxsBgonDK97tgH4lY9YJowVPKWOPZUVKhFepl1sM6Nb6XvMsLFDsY820e
o1+Nu/dATSi6fBXU1yMqomH7/nkVDtF3Cn3TJsabJ030EWgrh9RdDAP9wr9Q
2wOVK0gZMUdppNJI0kor0von93NyTVbsneYTiU2LvE8FSGom4N6l3o/uhAhr
QSRpn+GBnziGLR3yH99DE3+6uvqG3InE8dxHdjQ1g2hGej9jm0XQKzcu4dNk
aoAw5s4HUa8dngtDN5pJYWdN+Hvu5a4wy3bhW41mlTiuLAHZFKr4ThC6d5ik
JnnN+EQJ90heLTpVBCgB8mTQKDyacKRD/JIXkIVQ5SQyMxyksphQPqEncWkC
soVvbqoK1nnAlkWEG4NMSF3iMRbQkzu+X8RG29Ndbb0JI2MHPYzL39l8XJ0Y
krNWBWpFRLT/lYv+iHXP9mI0MQY1++jMdIAsLm4Y42/aJFjFTTXyAQy7LnJj
u0C/hmoM+q2hjUDaYQPhidSF4i46M0bfluzx8qG/Oo48Q6SakNR1vlZ9r9Yp
9y3W9UWES4AiRBl/V+r31Mv90JPDVfzVVKHs4Qz9s5Zz6P6GhMk+Zh8QFFs0
nB219Z5CoAxwA/paKDRwUX8fRcUayY59WY+0aw2ByzaQP5AUAND8UGFau27p
i+L65VBvsfx6SolAp8GC/Xi8GC7fv0u66kU6AubLqCgfcfYEgfS2o3od2C/z
LHFGG945qVqI/sMu/tCGiW24giXxAVsKvD8GDubwJ4TzGm7oTLMYzQID8eW7
N7kc3uakAHU+roVcBPWYzRuNbJ3QwhcJja9xInE0w8jhUa1annDtqN34K717
Hv+83V8sXBLPf2ohdNT+nrJLbb47W8ttvPC4DrGtGtLnbZPtozZ/qceyQ8WO
P2yOJUVqPhp9KyulparBtaNRyxE5Wxy3r+BUHDdkJTJ96k52PN2qhbLQ0V/C
bKrOS3mMM4Pu56T/2jrv7dq2q9RPD+GD/IBFgQQ70u+CTaDdLI3wHMyNUsav
ReA6cYIXN0NnoI5TAUgBKeB7oSC6cCT5OjxE5xzIFQUkbF6vuK3UXkkltp/N
BWMC6dqBmQGvzVvYmlG807EEqrhA7KIAtUCDGrpgAJo3UNCUAfFJLMvUCJK2
ZVcnZ87KD7ZNdInwXiBAZxuX7/Tm0dcaSlUniRn4d7/pE60lF32cPcW1zPqg
eGvmKp/F0AitwH0wAtbAzLOCPdZJbain6jmtdQuDcH3YhYysM25fewUSMwwS
EiCW4VTLaSXrMSzQGAqJ+Ilzl7oLImpNq/ya/ZuDCDy9Bnbq9pc2P6FrzzBH
iEgXRAwOVOhDYWQ1dmqYXjqi/LwTjZvbUz9vdmUE3l7JnAKsRGpprMuL+oUP
ramEoI95QfTxgZhMNqs9hYRTEflTPqo0St5uH96dpfycRHMTrpNNpu66gEUc
R2hFqZKj4VeJnyBk9RID/3A83yWx8H4f3L7m6AoAWcnwWYZRNeW2cup4NQzK
5GiEpGenQjfyNL/COBMPsFLHMAAIXieJ7HddvBu/XCrNepRAT2ekzK2qSTcz
MSpXP2lnXS0QMJfm4f2bmyGFHK2lUKyuvh7cm7wXJCVOx3dqG/q1VdfBgXCr
mYf86dA4p0hg2HYvdZzbHpzQiHyjIZcyynmhcpvIOzsX7X5PNG58Jmhqo9oj
xpwckl5oCx17gTJLCWCPWH6ps7cbUqkZVKBaCVghCFWdpSr0+qpuqSKU8UxI
t69NvX37IIpSE4n+n5lVvC6bJtCJtXgKr+o+R5EhodZWO5yZABYkqLtOdnFG
buN6cS49uYSUEWRtpIQven/J6EzdSknRMsyQWkf9TbMf4JHMiFRBciPv4OcO
RNSANScHAkS0JfDvvvCHtL++5fpBK2unSeItr+ci1534zZGCcZRPaBFycMdq
pERtFABF9FK4jy17HQjb/Lf9Han37aM/50GthjE3DP+AKDkVuBKXJnAtgS0y
QwCgrRvSG8rmgdLR5+JNx09fK/HJUZd0cK9GPy3qeZk9dMpuLbJyVC6bsrxL
SZ6doA0dy/8yG4DGgXVXY0W9eaAYbZT17zlEBxYVtvXiKBzjpetYm0Y2t7oE
oFqFQ8RuvuSCuiTze6WvuRND/BlAOLpKqqAswwWhIItqybifHnOkJT8CfwH5
HniefeKnc2mA7EhfPXJ+gfC5MbcPKbAzdUtiUHxx6bQ0Qo3NtwlOZp7t6CYy
3xb74fK5NxPfviKkxF4G7CSxHn75ZZa/rG+0ufFOFUrMbA2J5NVtLpsEtPYz
G4PW80LI8FbFt1XZ9LxquWkwWzNSTss6NtjR10/9S4azDRqnsJm7RPeyyzGJ
0uwwZVyg1SMlbupynvziBPIXJkkma3mUt0g7U/iLKUowZaivlPL8G4aRBDru
9GPTRjiGMVpMWeCPmBGRJ0dKlQiAhZRUTOQ0cFDs3muavjkty3L4NA8SYUXe
P5q8wsMqE4ft3KRFRRGRgxG6RdTFW8byd448+M7IWR45TIdpt1DYSOkCYyoC
1oLNROCnSAJpGE64M8V1yt9EtDl8CiXRDg41lapwpg8W5nDcg75wbIyJ9dxf
rO8TqO+mtiYo7x8xWh+86ifVI09X0T5NRQ7dEqjiXhonpCIBCzFGYMhYLn9S
JBqAWxI8bz1kIVY7WBy6wcCwYOwi7/LZOmHCadzk8HANOT3xzfTvTEVqzGsC
KoI6//rMNt7gAHXiFjW9yOmuna2xw1rYIgszE/G3uJaMv1DNlofbN4tAUnns
eO7n0kD5P6scjne8j+wtFWufPby5T46q8f7/DQc1XtWtQ2ZhR+GfHYRCILBE
7OzfoNeUhxspIy6dqfg2CQernBBBcTOxRt2gcBK5Kmb3s7wYgZHnoa5dpmcW
FCGdBN3IjT/SwucgJCKLKhsKPpp0QGB33fySq3BA/0X9o3xAlDQJsCGO6Q+0
3F95rIkeLRPYEvaejE3Z1nKnlaunZTNI8vWgdIOvwpCXCmgVT5asx+YPf+V6
eVGvEQOiLtiiuvOi72AJt1ogVxU9Vr+2wc0ogWK5Kn7qbZP9zOWZ6CB9cEYE
KyOi4zzWM4W0T8CTHpetSq99YHa9vDZtGo/it7SKr3s3oYxRKP2XqBeotsM2
O6udmVxQnuAh1JwMsHmIAjzReHItg9o/idWa3SpPCxfUppkJA0V6z79Vhw91
0RBbJGSbBWueUI07iacHKs7Dr5vGXuAXeIQoshP59dAVpOOe4Zv4Q7SlcgBE
RyuARt4KB4JQehkq58eI2InKnblgw7KaHtcotzGMKvsQn0prL4uKaRZRIyT3
N9gCXRVAnl9hlAAXhHtjrdkwTXD6KKLNUizGB6urKg8W8MU2xUuknCxlJU4b
rnJ1H08WTlwVgj0x0Hdo2BU4QEQA/gVlM04IPNG31NkaKL0HvKmLQkuItBzt
vMchKyke3nh1DBrAb+Q9lUwW0/b9+/XVL0tzNeNjnLMG8vhoyWig57Sf0AhQ
HfMXge89rVaanKV2/jorGBUJ8/0SzLKbHuBcK53s8JrdAOq5EVAs5NmaG723
XSr+g0L3IR3Hhye1fxCLIU2wyOk1UhC3I8IqJSDYJuIAGM4l+ZCpqAHPKBKz
iJxihVXPLPZ2v6zOjYVPqVZ8g6iujGeZAtGngMkXgekEZYPVESOPJlJN/Ag/
60/BqkeOfHDZ67wODmZBQGMG2ZdOix+O9zDZGB39kIvPX16Gq1SuOXy5383u
JUWv7qT+g0vfLq0oVMFvyxpSO1B8ZTcmArS/mlaBuKmNBzXWJXp+Btk3Sn6b
xK3Tf9RVgqOQDDnLhQcj5cE8XkIe29NTXjZoNtMcT1B8VRznDQPbN0w6txaD
O7RyPRBOWsU/2Q9cP1tEtnOSsjUoVTiq3jzcBffKCC7yAt3fM2Wo2+7SN21W
NIWqppSZy37iiEiesp9yAzdwlwyTLKfamTfVmFft2qHL239oUOyrSTe267yq
a0yVhBgJUyjbnAzGjUI1FlKu3MvHA6hUGUDWSNb9mWpKZ372eEzH5dBpDWUV
rAZq/qeHhCZBiIQO0XauOguWm1nltltCGlrapPVtmku07TtE/An2X2eUoyi6
fUkQHhJkM0l2Af8w6FWjWIu5748LbrKL2/ODGImQbfCZhvCdgbgQvyCUm7LE
zdqFqNTY3CCUW+7bXqhMgs98P0QRY6UFxgvALhF+HnIpcGP9J05klFG8rpZx
MrK8k/GHxVAR4lWT+z9gSa7lBF0p0j4cWMYZLhs3sQV8NrXLDz+48aenLLNP
zwYPDcdyWz3QbiXHaJU0EL4UU9jZO4Or5uqZP24PEHdKscAVy/v9LbOCZWa1
eB0wZ/DmJpVBp/Cgi+KcGBSU2RkJ5mlppBM2J6LGMkgJ5kWt3zo/Cmj5yObJ
6BX5RJM8KS7YY3U2uxfeb8Z7Idfx2XQ2kut++nBNr69uXhv2bJ3wDM0+QY5C
WGokabmoXB50xFBxR8q1K8gyBvUG7tcWqYo9FDPRmWw90DxwjMHuI4KrgP7a
0vn/GgmxA8KYRGqyhvK3HGTDDkHE/UWT5yplVmEUIjr8jd9WDvWub/NbPc+B
ef9WGyC4HUlAAZHsTPJ8oDNs1B9M9eWcq8u0N4xbxwQYmVksxzVf4qo6gZ0R
GRRT4tgxSljfbE0tLZ4Gyu1ttsuxKVhVgf/Vs5cmjsqV5yWKtsvD8yXv337P
gQJG21ApbNdwrsHHaa4VdakMrqrclxWjFOFv48IFLelQ0c+yIjJKGBH9dBxB
1E6yKEQFjLR1IsSEof1fAdSXe2UIecHxXZFo9S49JFrqNvzkluoU/OBVHUFI
g7dfl2lmNPrsiEPYwJ1deO4xnKfui4+ntM0p+UddnjfJFGZuyF+4O9nfanOA
ps4rEfKcC/xy8kyT5G3b8osqYD/0TEnKIYdriuluF8M8CbqM37nQXiZgRUN2
hcIPRgdxD5mW2KJORMUJtDqhsXhJt1zAn1lg7FU/Q6oCqJsJmCnxYVkhPmoD
K8APcGRYpXO3NevGzwZDulzU4vGX3izB5opCaZ0/Eaae8+oEyEF8SNUDYsCR
yseJTzxZBI+q8KI4SyePcFSmI6eGWSB1shiVUlWSLdmVoEX3kJpkEkoU6cZV
kXF7bvC8jvSCmwMljgjFg/m0iK14FXwHCkw4s1TMhZ9v2+8EIb1pUnLudpjp
dVypWsYoxGcmjC5EbVFnH8rVjX1//6htX9ULp8MW2MGhu3wGEIwLVlM/Pfaf
hEYD3yk7X/4c1EfpghzNHzvqy9UdmLxFBCKXBrHPxM/yd3TJMYBciJiiTDzL
7jeOwXi1Uc1RRB1ZvbAgijk4HrBRvAAy8vXYO9kE2yZAonZ4g2HnB/cgg4Tf
NJhU/ciGu5DU3ZAv/tNsiL+ypluqqi6Cm7h22NBKDspwSXM8ZS73zUTLs7z2
RLE+dskV6OTqI7SvmF13QeaBWZ2WTwSQE0w8FKITnXhSkbol+uvKbUr3Z20v
AkMQkMPLlIjmAvzLkeWw2QEXzSWrGy+F6bHpUQWTTfIWN1U4vNjWFDJ/uQsN
QJdr/MTKJjEQGAOp/WofzuqM0/7P3u6djYxD9nsRBWcyWCQZybPMQYn9HJ0d
r+gwNnY+ZGKURbtIWkJUBNfe7288oJcPW1GrdGSjBDlRSpXaZcHuzDAeKJF9
IuYEkp1IDcJCP6ZbWdmzjDqdImZHe9fxNtxErRBwSsDDznAxsOHA1npWj05p
K1veT2CdddVozLgVcLd/bo1/cL0BBSIUYNfvGqzi879kxXgABJ+Yv1Ibbvw6
UaJSlLWGD3y1vDnSSw2WfS9fVBc3g51Y3A5ptZSzMVwvResndHiODmD1KAE8
64Q17OuuzmQxsFGNXw6fMLfTsr7+9kw8KX6sH1UPN9htNKolaB4kgJRHEX9i
UGhuXiw3vC4AWtvDudQNVqqGYrd4TU1T0/I9ldVM34FTjZWdOHR6D0AgQyW2
T4Rj+c11A0DS7B+lFNm4GE+9s3MnawSFvXgTJX3vZYMeBnuQywVXLFPNPUf9
P9pJMDXhv5Bor0uu6Oi1KPbisAy2DYx3+U8eEYdufWSuZplVmjwtB8DRBMkX
HNQyrS1ikQfS7Nssx5UsPLoI7HGA9U5b920qDP5zPZXEFh1i7lUgdwiFVa/e
jeVJeJu8+RjVNIAOmsneAnwUapvnkEuMC7KVEPZUwBef38vuR7EZjDg4AnUo
CrTew7ugqgkqc81RA2WjMht4/krdlsFlvdkvWoan1HTY8iUswnvLcLTodwQn
4/gg3SHYoAx0VvZHLH3ePMZhdJ1NR/lkxRNaimwDTtSVBHPeFAr2CG022EfC
nz5iMBTynarx2QtZ+gvtFEqD7J9IUcxH71GOUl765tG3pSQjzX8tO14Qyrm9
9Ct8xLzEVsUnzMofN3SIEMZPPMqyeHS9tIIoU0gmIzQycKKcdLLzpwKhWakT
PM2NxHSoIbYU1FhRygn8WXfFNDwa7U87Oy9CqGVardeYECwsRg0iok8c0KKH
Z9aO2r7z4s1ORDz3a/nPv9+1tn4S5mo/JsQH+r/F65WDXc1XQgUpOZrPqCFb
dtodj7w4+dVg4se2FN00TGNHapsW1bfdEzK9BwYYN2wmmgrDdcp1VkkOgSht
y5+cFKwBzASmdUFnL6Lv/F/uEY4dSykh+lhD65hbmuLT5O0NCzy82+fuynrK
5AthswSKP09+vWSTGAJCYFRqXVe2hTUTZVEAecbPDQkFi9zOAv6CVCvNaQFZ
sCMNxs9p4EptkSTtfKRRuH7XPEIdQrB+uy8hVvGEErWNFAEKcuIxQ/FyIplS
PayXMBhAcrkT4Y1i1aIYXdGGvKEFoUiXxX7p5/Q5yq3ZhfWzo8zw9CprmZP/
hqhCnIMCufZpohBOLf1aUGjBA73378ectqtTchulvhpdHu6faqFW+RypAlbT
XkcII1G3vFZP8PQXzRhKF/yPYjseqQ5Ns79N1a9IoHUfnK24NXAU1p78Pplc
4C76rKyo10lYucvK02u3KvbudZw5AQm/A+Q+zIn+6NQNGRP0sGvxXqsJTYmH
9JWK0mTKxpsVJWA7bz2gUsLSOj7Sgwe3jZhRPfRhO+Leh6Ay9tHLrNARmSs8
Rig9oruMp8BTAxdYDHKtXK3wbmLYWUhgSpW7z+mzRdc4zTYC8fDIZPrtVVeg
zQe46WVSfXiHhF7X/H248fL3i4KetLPVCkwhRoW72fyXuqXJVlMVD6g5yfex
nb1k9ykWDaAxQakO0uUjv4WLh1wFImmEtP2TNwnM4NvwxYUC9mzOwSg+o9s3
MPQBcuG1wxgClo2kowmBcALhreJMEA0ndBlY5ekNVx7mYOoFGc2uGZ7jMDQ0
1sPI+bb7Mi/UsyZpz/wY5GByuZUz3WwYXjB5GuRN3JDbxJbkudzt0QAOVfmZ
Cp9SXWIkeM/cWrgvFTYitbR5/4c17T/Xvz2v8/ywZEPe55yVrMqmZkzSY9Z3
ML3SoMyr26Xk9kAa5HgWzi/jtXuTvBInK5bqB/0rdEc46fH6WwRIG3OobyqM
oA5B7kg1yUWlBDbi1dCbVTBfJknlqRJSt9vCQz5qp8vB8qiiz/+oQNSCymoR
DTYWIqiGDRZK0Q+XPBXgU4gBczGiiSsjqeGS9oWrBENErYL2PZN+/o0iholH
YlcOJ8Wyt3kNV3ylDL0KSYuzi6l7OFNMloAQv02NLosaPTRid/qaCE35RkvY
1IctVu+wS+lKYCyvbE9ksnYG5xnIzla5pAOGHdAo5IK38yxYrtvDQzo3r/fg
ESRKULniAy9UZSG8YgP1WXMHr2YH7SNPLMOpivm75k4HqcxWH/f/UPDIomTT
N9i0IgGr+sTPVlxBlW4oF5gnOkVhYaAXgoTRwXBvFxbZfmUpBf1wKpw57/hW
Db240yON2oQIZZKOnN1mY2PHDTk8If9S3c9u+qTIfV9ThmxhDZ87HrdtBtOS
plxQ+qbrQakl2WALospAEymt6ouplPVet/EFTBxtE94ATgOpnjYOabej2AiU
dpFvykQ1hYimLipEOD9XLHiD3sy6fbWoq2/xijH74SV64sWLZsh1xy8m2urT
UGioaeRL1J+4+YcJVuvgizLA7xeaQ4F89f2ctsgvr222mUXT0yT7TvHoXUM1
D27PVMIu/PbLID2NPAY6rLK6PzSKFw3IfBnQXMW7Oeb3XdUeKeqGiXRbHDkk
67BwSlfKEiSxSMPxzSKRi/cACtyE4r8ZQFEtuC9rs5/mL52S7f97YLbf

`pragma protect end_protected
