// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Yokw2l+PE6PdsTvFbf5ln9svQk3hEKtW1+JphgVHEcL2vrl3se3cGZn65zdnw8fU
m7ducrwqDbw42AmAZwVm0xx72Cf9E7LU+IK+xhSxV2b25coSM4TF3YVka2ZwzZDu
E47x8Ut2CHECZyO5IydVSCtJ1uywv7y8bPaRQaFogEs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 28640 )
`pragma protect data_block
GVUbGXMKTPcyclc8QOW2bOApu6Uk1Ad7cAK2JIuLZ3fkAJcUfg7Z4RExLZlV+9V5
b0XEGOFMzO9Th9dgpg9QxAGtjU9nTNePl/HZE09ooIkwUYWE5PZTLo36DMHvSaRA
fQ8MsKUpqSURvKjUbXr68MOl6lv0pE/nD1RQuvGUBFvuiQWoASpDbHDFpE+rIVGq
FhsrkoYu1WATxOdMOtCWO/UZ4+p8DVPiTgWINe/Gh9q8obrVdwiWV5241jLcQ0Nx
259roohx0J86Sv4BVAllx5t5sUEQeRaFhzfMtOpzkVGS+td7lzhhowb8gI7pSinE
nY82HXjYrWzfxA7a8TgUl8b1YvZyN31GCucnqrqxUGbRx7kKMLE9q8XuiDIAAUaJ
U0VUvNmdI6L2O7jTaMDyg5ZZANm5QfKWX/5GHMnSx8Nd5PIIW3gZ0Rcx+XMXOw3e
jKWsIKWGhCm0+h+JRY409vA5JNbjlPYqV/esQ0LeNun5pV+hmavCw/4hTZLz2apL
nafyrp4I7oFM2Z5ITh7AND7T3msZcmOmJejcYnxiGYDX7ArW7QHwLDKeSPSu/Q3w
GzWpuhMaccvlGLGGB/aDj402TtBuf4X35rtlxj+g1F+EEHwmr54/0fV0WleqXmyA
T5WjBRqZPkMDnPXQ/qthCMViV7uOOega45ev54KN3fPy/WvguWx/P1Ndwl6K/rK9
bL/6ffZWlOy72+CsOVGFTxNHsX33dUkkZxawQShiya801syDA9Z75dwCCPCB2Iqo
+X9SV9ft6Is9kzOMTjgUWtKA3tEJ2vhxKaZ2r6oq8k0ts67eePcgtYmWdADYNCOi
4J9fR9c0xnM7PT1CwlygJ61iNcOBja2X6PqTxO+3E1pAKJxIxMiNhOS3s6wPT1Ne
VE1vuE7pQsdJAJ0VmLHpe54qGr4dprs5r4Dztc/NiAz/RDGg77VTvnAUghv+LMOx
rgvYr7M3JxFpmnv6SbPkFnbrI9SHgee1oBDpVnJG2Dz3w+i1jdtV6npIaTS8oSzP
7QqsuGClm8hhtcHq1+TjJRM0MKA3aivwGybgkl7dNNTn3wmnCmtbV6lje2/AnCf0
Jg1HoQShLfw8kq5oi0vDm/tKMDfwkobsbJNoT0kEaW8620CTT/55q2kqeFPRss8+
vaOkGDGLuNd+7gggkSUFXxQgw+hRU4vBtoIPUQ9xAAEfTNqSLfCcJb2oKUS2+Ena
hAWQdBgSpdWBIZeeixyCCk0wgGg7wGq+KizMsFnOV6rQ0B+pqpcS616C0QrY9YT5
qHQg6QMzmd5efq2hvHW+m5EOU2BkYOqqHJkD8LSOv4zfw6HFfQeRUT8vM9KIavDl
t3cWGlvTB7vFRafxacRIsRAfTHnTb8jk53CzubUxlEqxzq+3VwjvvpQJu0bb+RV8
Mmww6Qke/uJpJn3Fuh29Qosd0r49UUcUr5kLqrWWufHLDvm/lc543GoXWC+M8TyA
frnDiKvErUs5Sm9xMNCTofkFMInkWacaGy8fxyt5v/lok6Z/zELyhFLIipmKAqRd
2JWRwPVw0JYrbNnxA1c2N4WdvyGjazswx9Y1m39xd5TgMtywOVkFNE22MO/vuecW
FAatwhWh6gw1bGiNb3Pa9yIvzqOWiqBWWY9v3jdq6IhIhoC4KwB+6YIEoVpGihaH
G1nUJslxs/gFeTb4dC5cDSPCW5PIV14nanq/Thh/cRSdAk+KxceHqNfZBHl7Pdg/
kGXF46YSRRjWLwrOYH/Ab8vA0SKJyR+H052iVstVqxEBBCvPXObUQZkbSBrDRdIj
dForqK9tmEMkzoqkCiUS5tE6qniV7aZwmlZ+NjqUbFkSLKrBw8zKW9yRG5MiSjqV
ZmNG0wLa7fThkOvRVdoviHAG9LhW7K9Qahv9N/Tzg9q2X6qaMpLfh+Zrafsw51d4
8tqdey/2OwE45CT4psEdixUuSwQ1AkZNV6gguiFQfRH3qiLCxPYbKrCoQ2+HT73W
OXjTsammNCc+Pd7w2BuGQ8mwuMFnKhiHnLrgbWOpd43hLQOyUuvtZjaTlm1QBygq
n0RcpKQWuX8Y/E07iHnJxiA04PoQlQNaK9Wuc49D8gzabNtgG15s1WROpR2b3+hg
gGW7UdoQPzgO2FagvNuw2baDvOVcsRreND5eOh1m2E4c8G/Jge+BybYVtJRBGTsA
E1YQgc88vJiOCte4T6ejEjMPKRlHW93hBSvwUa2rh/fpi485a5vWIyKTFVWPqwtQ
co/Blxe4hoepNyIprjWZ4jpb9obahhefe+LVn5REzGN2BZX8ezhARhykcaAUBjVp
k2v4KeQiPR7Chqq8ipVhQLDjrYKGQr/bwrSzfZdhrar5LgCLMq90PbqwU0H24XVj
E166XbgtiscxYn1bHSjBsVOHIrknBSo2d+tWF8wn3xFsAXRiSArZD/OmKnluE/7l
CyRoe9mA3Cojod3vu1yVufAVE+8tdpsziaunOqmzwLdNk3ylieFWLsh1+BkxosTL
bnr2EkQhQLiephwW00edHvZYRKjgWdROUf6PQx66yog1ZLuapXWc/v/KZhIHfcEv
UxowFX7GcsgIBe47hbPwaaws+IqlvXbsolxHIae3DGn9ECXoFN6+r2DGwQdx0r02
NewBOZsTXiDkSrj+oj/Dd+sZS/QlA0ntrakFINLwIoI9PDDtpXJ/mrdpNaYyDQfV
dgyjnd19TwX3HFhC6Ae4X5tS1aRFRbK9RiUazBpbra9XaFcFlLpffYgm46S30fXx
yVYxsLnY3PBCEvggJ2q6BTrjQQyVt1gQwu0xj4JO4Ywj98osbGrQ9ztWNeaKR6SE
BRXMG+iv3eNH/9nsRzdHOnvFsF2ePfQhsjutn3t5x5tZ3H6VxXP5UYVx3CahT5/r
S5h0LcyUuh8AVa6NsCdOH3Xz/3l4P2BaTjDI4lzZZKR2El7j1/14r7bh3R3QFcEh
wuuz5+xhOuGVDTIfhnlrj+EwNbS2cJr5zChN0zZKEpOL8sgHi1lb+1FngBIApZgF
tp5WEwAlgP6BgitD3KKPhx6FBPwc326O0UPRoQO6ec5KIXHlaMTIlwr8OahT6Gm8
IsuKmiISyw3yKv6XmwDafqxaqqzvEEOIdEq7Jp8PP9JiGXt5G8VjnrspY5VZDJhX
Z3xGSZ4vK6ShmsCo6ZkhDQCu3SprGInM9Yhu4d9VHbftTdPuiF2rwErxosk7kHj7
ne2V2hWXUAoX6yM5Kyn6zajgBrNkrfOWikiR/HrhKNUkb/Pk9GNxBt7MI1+raLhJ
+6SgDZRgaPetfaEqYcQG08zWRzYmIHY6oudZmhMgxExSrlMyw17R1PsUJtTr3t0h
wbUkylL6g6HYmJa4lw89AMRPXhT6ZU1HzpjlgjdAe8CBZ+WcAe6ksL2bjte2yhAc
pwzgZq2R8QDe9cMyzRLSv6S0gNF04A4UzAytKTWuUMs7mGxyQiZqVQSNco5ZuRN3
Wso9dJQHypSF75A/rkZQi97O/wXF5zVi/vwLfnCmd6yHoBw9dBD7w3GNe82V+lL5
kgll/gJCrOciNUc81I0Ar7RDwtE3wGxAz6QcDH7sJpIbJcyN72dwuHA2L7h1soTx
9s8gBw7sH1WRC/yV8pa/5p3AAKWgCkbkU6Zmdnqjh9W78GT0uMJuNL0utlGZGP34
6/9YJpKLwqXjEZ5Z5RVjfg0YRcdDYzRx2DxZOKEAScRYwShmi+hHtyfT7JE2vTBa
tSM3eneZdlVJ1yG3cqR9J9afaEDUjlv8Pg7qKWzpZv1PxgpdyOSFdxbqG04MLtUw
/dRmxLHGH1KdhwT0TvM4ZbycMFKcHy+JhW1Iy4nOq5WJY6EO7MIcWkVxv+rBgYL6
zSy7u+M85VSfvEdywiQcRzII6Nzksk+oLesOJMzzEE9R4+/C+UK6hTgRBSka7aNr
qOj+wujL6XOYaDfT4rn+Mmm8PUH2HmhLuwzWNl6PcCK2xdWA1KqtrEQ+1yT/F2tL
3utigaoxFKqJ6Hd7JyKTka43kIcKMUcPKkmQMVAHD6AhPT+b3xs3+YIQFcAp+giR
3SnPO0zzEPTUSyR11gb7fSCi9uvNf3A4B5ETPrilGy85g5x3OljOlEpZBcUwSycV
nK8TfSe+iJACoveSYORiC6b0D11qf0xza5neZLXHrdvv2m1VD1fX3ex5calg5hvO
v+ecSuY2H7DKFfvkEMdoqbxggnNLvOFQGqSMXMN53dgLLT5ZGpHUK2e2a0dkpq/D
WuP27hVqnQzfeayapOEQwaCTIvsrGj0WFE0JSkuQ/09TOohmlpjefLwMD0Xt2fTZ
eshllDjUYMcdAC+ZysT+PADh0t+iz4wBq6kOQWaMDNbPWRI8w2APxpg0DsAxI1rJ
3CxzxXe0PPjLcT2e63a5OPJBKfa3u+/ZPkR/+Yi0Q3K3CcopMR/EJtGMmjBwW04W
bQcghuEHAM5OkfccWiuTmVxQxeMBZrT9hMuM5Irrshg0EDryIFxem/9MOYPDOFbS
dPrx2RwqFpn+1agjsce2/kKaDcLm/r5anf37eSSrNZMCX5c/7xarfWzywkLK1Qru
61I1jKaQgqK7u2dASxc871ySxWLs8MS14piT6wCOS33AxF0ZTrHQVwk7E2dX+v9Q
9LrZmbiA9hIeLUxR84jH2vXDXMTdU/hu5K22OGuR3bI8d9vVzhn0SIoIdiPuV11a
2f1CrwV5DCGnT1I5aF3w+due6AwpY8st/gU0jjTuymWRq4Rp4b1StYjf3PteFneX
cd3pSFL4g5DfuC1zDhjjPDt4l0C8Y5Rr4kXNPCPR8AhIB36Oyp5WYsX25N6t3rKM
q2bOMC4W3U4YShy8lcLXq1vZf5L9buLgaBCFBki17OhWR77s0mamUn3iT4kTU/9P
HrWl4fbDNb23Y98LQsdzeFYekJcETJUvDS3EUBimUZ9YYPmoaIEDWnmVfrQUzooo
oDKbicau/W1bVaOMPwG31oUIfjuGpeVRfq1u7HA/6ZDt6DpiiBTGJ0VIHocyMnB1
R1tQo6ggiVwrVvVcCnnBaVbFY21p3nh61sS1a8d5F/sMS9iE+0+SaU+caISrQbrZ
jMTpyvLB9W1lARJ+Qre0VrfxZvkeCuyX61z9e5wL+UEExNwlDakVqSeJrTJkml+h
WJZXQl9O+p0SiJcHnTmu1973b3SdCfMgwfcmrIfsB7O7P8j1CnD0dA9vR3kqO9/T
wUeaxtHcHhITyOieJ+wNlUcPnEvHKdxoVFBrwV6GZxSMO7HrNO0fmKuqP48kPjck
WgFcp1HhKpFAzmEsJQ5FWpTXSHukknlDfQPRpcIr0z6Ho4zddrRh1nlwOQtEaT3+
yhPM3owLYnE0f/+5tnJA7bHnkLSuuFtsp35IhMG7pyXnDQe8z0aA5U/dkc5ANIIC
J1OTL9YJ81A9a3qg38j7lGcLu+dvcP2HBMPIvU4HVddCJ3ZDh+XcDOS9TebaX2+M
Kc162CZhSQ7ZjJiAfSeOfN6//9kkMXP+0ygTlUsCKAinMHg0VwroeoME2HFJ72rQ
dLMx7XHLlmfK/a9QY5xD2iF9wXQnzfWq0ZdsMP2Zno0HYGjgKDVTt26b0uVDNZJF
qWlEGHqilQOE9LSRz6JSfsdpXGH8XRhjb/jnlwlqDg5mle7EipDHElmjdIiS3HAa
8LV8Nq30EX/HNIy10Oj1WS8nCxWAeE0bh8Wfin33utYMMkzxvSfz9LhWbWzT3ZiE
ElF7/RgmstsqCvEKpQO+YV0vsNCO0TH0ERFZbj5d5ag9BQ00AHBhGeUImTej1Sqy
yQ0nXyigTZABPoNZ5rkbeL7YYQp8ayDR6J0JjGnHyh8MurUlAowTxI7LKozPNfhe
MSsAonomMQ0lEwLuF2ubrjPUbssI2r1zF+85qvf7PLD3r6IXI9ty99/eU8+qi6a9
RAifRmVaudY5TflC7/i7SMfb731INQezOyq2zR4Z45xX+BxNQVgmE/g56lliUM5M
oCeeNaAl8y3GQwfcGpbvgYwZVb736B7GQeo0y9viZBUnHikDE+LM0M1YTowUCqxd
hVBgTrRPzFMgioSCd4TAGAidiu+o/UboI0VyCgioQduympE/FdlhN2Mna5LvHVtx
8Vv/gFElaRX2caVv3kzYLRGP7rvQrNldk9E0eA9CgRp1ASfa1+fyeMD/PcwxVjFB
E9XiKZ7mzLADXtmCkMh1GtN6LHWuxYTTZYKYpDLvzqQK3L/01UlxOj9Lx9aIL6Pe
JBgffI3m6NzByjX+c6OsOxIFE5kdhehrfIffMs/L5tHX4PuleuYo6xQ6LS3cvt3o
pB3qba91PQ6OTa5jSKhgtlab4tU+deRYX2ke9UnMQ4A5V12f7Gj1QR9GdZKND0bR
G+DbgKyuxIoJTYMMKi0q1ge9yd8l1qTeIvPqOPkOnMycd2c0prOxQMfPgf8utzY2
TP7f/zEJSLZN6Wjl8dwxaDC54TwIagBUQX09v8hv9SLKnieYFvUf2XcF8COYvIUV
ALL37hMYb7jA0GKdORgWpR15xc3e1xj6L8nin4WzRRDyUlhQ7yIHUXWdqtEsbbrd
/wlQymScGVU3fU2HqgbJCQ9Ow5TdGQGjhp6uV6udHNY/QN97rV/PA18AParNrWAY
+Z7B5VaPV3LXAeQT8FB6Jkm+MabRwAbtB5KLIA1HK/eA8bq1u3gpDJsQ108hDQxY
GEHhWa8pzXaNVaJqnsVju2XkjCKKURCOJyr/L9MOUQ/6lX8Qlg8kXzpgyf+xAbaS
pvmM7s0QIhVP2FyMlDCFVOgftgEvQIjLK7YasNAqFa21cCEoGnffAhDR4ZiqThDZ
nF0kyNrjODV+iNmg6VfNQt7CHHnYTuXJWGMqtQMNqlD8iL2mATIcFE32RUWapWtY
fBjlHhlt2T5z5MMwFtclEuf9HCdD/KRDOJ1roFS75fehPFStl7lPYB5GlfnWVByy
0KkXkuwuzuHa4cyTU7l0tuQsY4gQQilsUC5EM21rL9OvdfwT9149vLTXuV8HIEnm
e+iyzqZIOealtsc2CO5k6Tkz87m84ux9laENGAXpEiOllUUuP4ji1YF0FsZGpmkH
Qn96ZRwxn9dfkkqvwdD0I7JZyyLiWBrSmNmV6Aeuy6k9DUKo3QObw4RqwMN5wScr
lHkCqpsb1hdj7Dbt98WUsqN7ZzteaPJr7sCzGF/DKzZKk1tv7+R6KwLPJGD47jPB
Eca3dmC0L+WTjpUiIipQinHEEvvXYvm/ITef3Gbk72mznKab/lHBM+KbpVAu2B2S
cQA87nEUNRlV0iKN+xNRNPTIYyAC161ElntIWVRkgilA5kxma4nafHPmXvdnpr2S
2huUEfv1lUrC7vDX6UwML70cu1hMEBNaGa+3dNCH6VHJsL7Hermy9rLeXub0fNnq
S1nXkY2g7hDnyNB+97nC5KFnw0zN6RjmATxi3PeOYeTx4xbuodUSoXx2GQeHhG4D
H8fNEzso4E0Vz8HC7v6iR3UqZxsu6VtfmuRTe47DVlGYIsiDIdXPJcJ34/I5ILb0
NnJM7C3bVQtG2rBme1aeyOf2eqBIWWlKjIaxj6sK6glf8DP0rYZBl08gmT8/o2DY
EN5Md+HQzlzzCsvDcZFNk1RgFXreRdvSmo3gjMGJXUJDsz19Osw0LWDAY8xaH2DV
61pfDSP/CmrkQo1dR1NVeTJuUtpmP1G4yoNI92SLVnhMu7FxuDUuUxrfYRqDOba1
78NkrB3t6zbifNCQzKp+4Ako1vXYVyzFHYZ0uxmUocmmiDj470dcMT9wXeua3xFT
GCOmjHWHMxOVuYpUmsXMQq18a4G2zOIniFgz0X+VZixxa9JfiSb1E9ZeBmL1uI6+
Jdnnb9lpPcUkBEWR5BrmLaBJimsieXDgVKngDzpyN9MxIDBERCjAkkjF8FP0NeUx
YiC4LkrWOfZ0dcpWKYEF2JhnoWp9cWZQaA4+ICNn9sO+f6N8Bd7Tq1dCK3bonReg
yJxdB77OKI9Nuoo7GlnnXBDZUkmtIQ1o8Lh0ZKAVoJGOLeOH4nnxKShAaNJWVWPd
t5ADUfJuIFeGkyzfErqG0qVO0qZoxnQT/KZhwGaka0MCRkM0/cQFQ6hk+DY7krkE
T6TMuYzRgp/7IDTr/tkTAP68lhWK/HKulaFIrY8x9w/17NS+Xcjx8rsYx/j/8luG
2UxQCbNyK4hjpVKfTVwKBi++/kt//c5Z7mbQ+at4R/kdF0GQF/a589Va/GWASxTd
f3264T60/cWyWxLGTHn/JWx5S0lnVrfKiU2PWFOaPk5QQg1FZaXp3E+y4Arq5zzE
s69JSs1bs13pP1cw2yXK8TZDrURhx+XfZld/wgC1hCWwWAle2wTkn8MF8v/Yrl87
eoIAM1MGoRuvGrxWo8GPeimUw/5B2Tpt6ltdH3XzdgnGWBfjVobbnSi2WtVdFwFF
9Ypgi3NZ43IBMaKVTnpjHu6VysDWSf2tDa1MhzA60qWVPwybwr1ccI3xzZAHeUzY
4bv4lAUEujtkNlGqNbe9StWOBzEC1fNYXaH/qsg2MbyqpAEK09UU9z1+onQVFoqb
w2vWOIgJvTxZFsMPVa1R5kULFE2Z/IvHB6wH+TXSY2u4Fb4X/GPk6LQtSEcppXiF
P6mGHB7EOFn19SluBhS6eTnMjGlR+/RveefeIg5/qJCeOxxutHvzjbCOX/dAHktv
8ceWwIizF9NJfA0ywPwkCm2nl6Md0ihxIWlz1F/7qOZtmrmZnnfomY6A0CfWCEKk
LJ6WU1JswIlz9RltXWYx8IcACfCthPP6B6FWEjXk1bV/EfCtK1IpAQKcF8lXTFHV
q78oprKhz31p3w8sLS4y+ynKQEE56MUlAYsP944DnXGmiNB9b8MgApXBUqlKNUty
w9eZ3I8nRMCP0sdwPbbxtkiwgBwmI8st2S7bjFYmmI7OVTcv6Uz5gD2cdCYIOxyi
QJ1RoHBYDpldLzDoZmILhdibFCI27AYsvkjwsqU821EYnajj8rVtwz9L8FMVXG4P
wZ6ELRh6BodbtssZ4AIIkmaV+yqIdzodQGTpr7uRvMJLbpD7KOl4Z/9aZCPbfQuI
dNk9Hxk+mMdumr8R46JcblAQ19rRoYSrwTXe32mjBZ1fNb3vgEbDxerVAf8oYhQK
lG8FmC12eTFoyOgBQGOJ+YB4ky1CTU3cOVaEVcFB/rb5obG3BYxk/nko294gxmEB
Ful296Z9M/KrIwq84isnb/qzGgu/5QZ4RY6hJpd3pc/rYlMn4Py3UtKGdELf4Cni
5njk21BFen+A3QUu4gENoVhdAkYnszEzP7xObDEqBQevC0TkqmBOSRaDdiurx4nD
UV/31jhSDS499YAiLHB0lxlPw7QZOrtEq0OyW1ew2l1paEnm83Gbmtu4Hr859l0v
AAYJdKHPq0dnOkFUPj7e38ryLhGY+5MZl3gbUGeHs3lojX7l5Lf2OPUY6jaBrUul
hSVY1IDMg2YQMSWRdL+rJqCrz/Ss3+ZemSWoWvVJqe6wrhsS1DAoDz9T+kqDT/HB
c0Tyg8+IWNnCzHCorpKDxsX7qje3L5X0hQo9jD4N2aNgE3QnDjfB/8Hw055XZwr+
7FoKVc5e3fFlk7Pr5wQNF0KsE2n6LXXmcsZN4X+Un7G+Zxi7QchXLbgjJK3A/4bO
9OY03iAVIXOjILtbfFJerOBVocNlVpl+a6rLiAdjUH3BvjoRwJSKyhaGTycsQ9PK
CA+PJxMnpuza2wNfKdxB3jnNOR4hYhHtQZ8MmsCr1wlvflUBFSct78sjqQ58WLQc
M272K3xSC+cwV/PQ7X8RizZkHxMzxhsrebslNmzny9uV/YUZEYf1CWr9MkjBQOSV
54A+qwV/veicCEcvpakSZVgRZNwgpbj5kKe0llHx7NMvopSqCQbncGr66VbIKSyW
SdLaoHaFXSESgP/Ps2nmXlThYaMCK8fPGFvvNyJ9GfbSuMCQKKQIfRkAg4nB0Iui
UV3syjNUKX3UcBe0leyHuCH/7/A0ca6BXNfo1yWKLppbbzMCwSLGrjU37zql+x41
cXqqtErDmLQ5H3NRQEOJ8Gj5ww4HvjqWLA+0sPkP6fYbypVdo1yqm9cPuYmNzQE2
HCsMW/Sm4Hg/hBUHE28dqnGfmzSZgEYsn3CagRhsVKobkdcfTSh/8U/jczrdtPcy
FnRLXdhVHHxQIJSCrqLn1agTZP9p175elNax48BSfnH8RfYfT4QACzcSOYSn9nqF
Upq7VpS8YMl00XwpKa2Ui86ro2um8uKZkZBOUDfA+HnXsD1Nb7glirV4J6FTnHKS
O3Xz0ikYiSxvcDETQSPBCItzxjlsgLcEAJ82okRH4TUCer23VJvRKAnP+POEns8p
JbvGq3AyVnsWD35Lg0ozfYh7+gczupsPaQWNn7y3i9imunOv4gTHgXU+vvh+I4+I
etKyCd+UlcOJm3pEo0Ix0fhlEVTW3zd19H44fTPiZDRvy+horx52begesNJkwsP2
GSGO2DhznrfM5Kew46lL6OgDXvepmBlmqykAAp6ZbYUWlfKVq1xkYaxELI0o000r
uWgqiY7K6Abmye3Sq3TkI+kZI0Vc7A8VETuaBHmt2CcXR62Aa3AU1qO8FdqV/q9h
qw6RYx5waLHuhPfiAdrVQGiR8SQ27QGR7QqoxhatWazDsx62CTGjakVWPOKUQdgC
rYYCRilqoyvyamgktBcFyv15kWJ7Ol9yvHOzgSTh2nh+O7kf7BJEGnOyvOtjpYym
qmNuYUEWJ/ZBEfJg5M7m4BYekPCdEtMBRNEkpRpIFb9n4dlrOkVMHB63gnZr8H5X
iBwzuDl2caaijwvkSfj+HcZihfeeJ8GQgMNRa6F6DJbXV4OH8kBAuDI9E3rr5e7I
W3uEn+CuuVdQnJyZOlbsr0TuOlUu6nVb58nAgsS6P9Z/0e4466YI9tdew2ovInqP
Lwt7yQGy8s/DYlK00R0V4NhDE/phP7SmgTtC/XXCqFryhnsqkIM27HiCgx+tqaxv
2Fg+3ZJs6OUPwp/6muVOjFnYkd3OrWUCncODbN4dGPaVpWRgm+1eVPl+i+nlpYPp
aXqgqiinEyBP7WpDs2bMCf0lcYeSeuqK1K+Gxhsgx/xkk77BBUIi+xc/Vcfrg2PP
JNNhbq+7IwSgniaO2LIjSn0TojDwXmvm1ck1ci/mptch9bnyV6UMb1XRwR/vUE16
SUXl9gdHyB1Dw/WvdAw6QeyD2ynodFarsMbjegWg2NNiCGDXVYWIQ87vV29sKryD
TcyPQYHb9CTqx6YkW8CUh0d3ov6qnTbtrIWczeqK4Aiy+N/KuDjXM4BoBRFva6JM
bCvzWgvTxqzlafPTneeeeTngsZQ4yRXKA4RnXnig93P77c5dkByQYdusyD7bDyUs
a57/h3O24FrK9yN6oauQARIicdh7VY4Wh3LEp3LjqrVK1V8d09hxmsw+cN+VzDAh
SZRcO5qI0kE1zJL7wAzbQO7YNcNps7QfrsJLs0mjGpr5jTS7WO9sYUys5xzXHsNT
kDEKf/Rvim0OJ+3JNjOPJExl+kU885PF/H9YljSXUrXpxfNUYz5gkLrs9Izh9eWr
xKanOUMbTQXODv+YP7IOlmdr9NixXSJrdegcABDXIqZnZdBx5kXuxHDHaeJRE8gz
32uV5PJtc4jQllUFPaaKbiKyrvUuQqW8tdhWcSl+77u/+KxVNWxY3DQYta+1xDUw
cVFwyY2+FuSRe1LFvt6XyOi0Xfl4b3rSUHsElaPGPAhSEBIda49ezsLyFwTZmVAf
IGfk9RSOievl3GiZ37x/JD3d7k94ZkBm+L/shtSVqmXqQx8G2CD1FJsjQpVTE0iN
p6IOZZwfpHgZXJuuBVpbMz7io+K3fBYpAc+Y2LKPYrSpgAfqhO7fwbsrmbj7Qzvn
36Tz+LzzM85VXv0SGNynWyR0s8BYcSErgDC0M3Tc22n4c2JeGfINApB3fRvGrHy7
TAvaK+adjOyMYBCVuzaG3JkuqZv2x9jKesc1vbbRV5GkbYJoR3hUhRwUai6hDfTb
dKUeyZeJQ3hBlf51FvsxtIgfqKaoXXp6d1JpAonB9qEj3je2eDVHAReKemNymD1E
do4G7qLBJ7jshc6w5WH8W8nkGgRAiBZ5327q2aEHEQpOLVxTSfd+rPNDU3smnOya
nPslRCYqo6OFLGUsJed0lun/W2OLpWtJSpefgZpd+29Rf4AU+ypKJaNl6GxLWOQH
prXyZ3vxDrbcQwgDam7nez/npLcjkVyCjbeIexueuV/m9rYQ62kNcso1aaf4NdKe
G7tWun4XS4jMevuQbtlArrRlfW/pwrgOM5OLzD1Of2dyZXnokbPNsrpS+sZ+/DiZ
w09JtBfS3uFw4YhClWpUYZw/S349Dg2iQ0GhMLeGvUnoFH1RmL7LS84JLm4LFZ8y
2XZ6tipSnpz873LwOp2Z1FyhEVw/LWVZAaX3G6vaUIVUbsrrxtIkdsSZMr3uQbSE
vdpNYCpEiHO1aAnMxqQKDd2QI1NQwv1/xZVyOZj/w62r+MEMeOaY+sG4WR9zh4+u
egJ5t8Lz+EJXwmXUiOfm3mQmwbMU45qsDmYQBIWymcWSNh2PqAt93376mrTProTo
xmGMnMpGbjINXu/pCGHhvuV4/Bopa6DDO35Y21sMICW6/nT9t2gCIZ5AIEJtwrEp
c/Pd3AukGogWqqSAibq8EDx7dEbgmWVGqhcmkPYN8A9fjHdAFCYQsrNr33ItYsd5
fWLOyct5CbjSx5t9E/FpHxJ9t9KnWAlz87aqF5acYLQK/CmbzFcKyNqrdB6mzMRK
1cNvX0/Y4Cp4QJpkZHqeVufdiW/c0/z5pblD9NVxNVSXcJclc+zwJrwXO6w/Cg3r
m8xtNx7EAo1pnD1RHqvLjggAke68stVs5m3jCtpYwW4HlDUrVqnQb4sll4N0mKuC
naxsJipqmXjsCwx3BQ6qoK84G9z9l1I/yi/f4XBVPdNmRXBg18ts0oujWnD6cU8t
kw81+JtZoA3EZ1A42k4wA/LHJBneefubrrXl4zlj6pjMkEyEk+s54ScYjFuTBgP8
ri8y2TPFSz6bzxpdq8xOy1lrDTqp7JzyqH1OjMMt9TeeYp/ArUqdLbyLt64DPlc1
2iSheFOhfa2ChUbF2ja9hGmsxqpymYZETM48lI4qJafvCrMRKvqXNFy4R3XhmJvf
GW6As6zW/Sup7ceQn6YFq0iLOMasiMAF1WSx4D6B8RArunUSbKULS94C5ngsWmLG
hRUKauBaygWyUDRjZYdXYMaJHoMy+fPTyKAw9YEq+6267TNEAGmlvZfIp2wLCTBH
6Ban5p6/wXL1lgUijcXuJBdws8EUafjwt1SrXUDwSq8dINJe1AawEUvYMEwhjWl3
olaGK+DihYtGSqT0BNVbSmMCBIr6Q0+2yqX8W2RZMoASckK+BAjULjJVimRnyGZv
BfitgsZdzR9TtOR+caVA+7lG9Kc8KG3Mtp++cH4G0KxSIxO/MekvjFCOkF3kvWrV
wXGh6pZGTPUiS9VmT0HQeT0OPy1nmQz0M84W4Lr78khBjCrSr+pvIeUMIjJ8znLB
SSD9MKxgCLWZo9YKlAPMMjrkDI63kbZEnQ0DjT+ThTl7Yi5/SlDuPmyK/lvpgmGj
fny0sYwQMXPh4MCPV663VlB3nFqgvnE9dbv4cscWcg1lVuJb8XJps9ebDr2o0kE1
+Mq27cVPoQJ+ImHf4AfnHxxjwc8lDoWA+w9hzuws8Hj69sNQUCU5TXk0eKfb9W+B
qs6Gyx4j2JLXcIdtNDSMEXRSwuaoBzFebt3t3A02RS5pde5zAX04I9eEeNiW7Z12
+nQDSphmamHtSJ0OhWKIDnoMPduURVVE3O6anulvbYvMFwTeBfCU8XtmqfQG94ae
b4+Qu+t1bNh9emS8I4rlw68hNa0rVEUid3LDl8KAtkYAGdKmjEfF+pZTFRZI3hEL
ywkfzH2Q8oeh6B9HByRu8snmXYKSyt/qzryHyqSHXgoJRxtvxK1mhSeWmYHgCiWQ
JhIsKK79qsVYwwJPNUcBR3t9gfr2ycVeTGG1Y/maAJA77HCvYqUi2i2D6uHaT1uL
SSrzgeNAFH0g6fgQxcsnVr20jEHAfF925toovCZ4ALpTK6rEcD8PkFpvrARjKHCL
214ac5JZziOBQmOUkB8cD7pwTkXK1CV+5Yru6ZnQUwPD7ty0pgA8odvyGlGzR9aH
mdepbdDc49qA5Jj2zLgKpowruomzd7LjuC0L9sv6IhhBr9JaG8TFbib3Tpc1/w6W
aRY8RM50opBjQUIVIhw+SZSjfcFN7uUh9eecTsRqegVn9QzS0Ww+ihqCCNtWutXl
ZYv4f5WgzqEzXhKjJXDo3t8J+ZhangN6rTusX1OCuvaNODuqwY73ebRhgUDLxQ32
Ti7kMrZt8QTxo3eAnjxfJzPTDxAsVLFDtKDAViTkQybuoR0NL53Z+mmY83c/ve6R
NNMVTpdIoC7ByNeIfeFWZYoTEIZ8sfMvT9rGoP3HNWI9+KCW3cSNdC6TSaZyPmXg
YOCfW3hrfssE6QTUobX3oFiz91yYJ4yP6KCSEsOjXKeSxXnB1pgPWffEfhQamdrx
s3K92e7pUouyJu/Bt2u/PK1hP0vXCO8D9B6YN2bnZ3g0MmlGdKTTpNUqcq77/IAP
334muboE6PLKRXFGvbCO/+lBAxveu+d9Bzd5Gy/fg8aJPna6crWc1OZ46OZqilV8
DfNi9oc3t+TZabLBmMbSyXdxg63CKiuPH41la5OlbNYGNes5kfDb5Wv/dawz9iFL
+qSSMWSGZNHfy49N1CP7HxNSwnOGWhtStSFB2u42EXixa7ITEsYo6EpwmlTDKdEf
sU6AbPYwDzn7IIqyO85ULVxVtnfBMvwvzeQrP6P3jWXP/GpqelF2wUMOJcBHTXZI
3wX0BqDDgC89xRWuCYSu2Nno5gn16rHeVCDe45kXgYPIo5gOChmizaD2nwdLfVf4
BhwiDzR5n7/cS+aWnZl1wwrdicu0wbDGgDDlLzHhYV+omm1jDMrZO/Jtjh8K+nkG
aUxiXGQeBSdEjdJOE03CHRLq9dBGJDe2q7VZfUSAJExEFZGvDiuZs2XS8Q6nU5do
BOFZgkj1IiR14kFY3/Edy++qC/EZQuOak4WJXGFuiGdjY4wf6ZpFCgDu34xXgYeE
UnsCOKwBaF80i2CpUF/+tB4osCFjRILnMrM48RHhBGCWF15nNo1F7FUg46Qt2Ozn
iwkPHfHHsZnczKItHzRh0Q8CV7Jg1rx357ZL15CZaWrEbu4sqIFGK8NobAGrF4/x
oP1gN1X2/VQoyBJGAwUkZJG9uimg+y9M0n7NBm7sSq99MWEiNYuVaeVNxrzkuEMB
gXCA0IQxSGSiCfrmwDGX34IZtO3ba5NAV2AHde36TCheDXg0qGW+9du5iMv0829p
92UPuG60iINyMDsh6af5hwMX3OxiXE1YUv5iPhQnAD2JkkqF8oFFH7r+JKNZXo0A
yJ65yHmpVZHidUOnt5Bt2eNbBBW+RrT/tUyxGDqJf96jQcfPs3WFQA7c7H4Ay3BQ
JYQFNSxEX7UYl7I8732UaLXDUCTiZK1vB3RmtVMYzDKGJtcqqMLI+YUKz6kGsm+T
Ld9brmmTQDvu4Y+adA1KR6Q8pT3szJpojkLaI9ej9YI5G02VTFFsW2ENsxJ4fRP5
AUyAMZNPg4MsQ1QBNLJYcKQmX/43Z7AalC8BijSMiTn35/YWs3jhjBld/FZqgcJc
0BuahjWdrdS/TzP9x9hA2ptaFA4P45HUMtVchzjjJUgjvLaqi3gk6fl0ELgUuEJL
muMXWIWK46uVuvbLwr6adJ6WJj2r98D4DgYz4ZHvZgPXONy5UTadI8j4dIcWB2KT
YK0+DOeAyFRscDdicbhlCO/qYesQ+snxtky629YAfv2JJ+srxecOq5re2Dj5+j67
rqmEhXwNUdhZMbfYaT+9gRtRcHxJvG3G+thB7KaRmmsQ3izacoBjO8BA9+kIzLdw
wHFiLrfBOosZ/VUsQJPOHWFtHRUttaGAs+kV4FyNbsSSSN8Cp4RvoJmbzT33tBY6
7W1cCeSveaDJr5E+6eTcOxIILtaRl7J83f3eatCVjeAyyhhEfKTpuRMtCKl5hi4G
1LK1bVnFID2pPDYxdVKU+mr2QSeHyWQKdKRABd+MHJxp0giceRXEaG/Fpd/8gRGX
pSQbxDHHmw/Q78Zcsc0MFScRy0E8nvRObGQv0tcK56pjbVwpwsdNT35BNvxJOCAp
vfWtIpYvE3haYXFNWtHuaNLGy70TTMjnAJ+DQMvyBSwEbMCBYFhHYUqMO4GWA4b2
dGNahnQXW93GtDMzxgRtjzC5T049TLgzVkDpCqN1pBEQd2Vagpt0hB4NwWiCKLCf
lDozMSjHmznXMDD3d9XBvILcTt1CZxkHbMbEjP9BImNHHMdcRCbBWZAkDdBZiZFo
NIW7tBPO+WWuVeaZjBY671jv6GhHHLITSZ9BpLA8oAjSjxCt/QK64TAJ4aE298Mx
unJKVHvW46su9Xx+0p8nG24YP+1sjIpBx3xqn5EYHh3gVMeniLcHjGOvi/ygCkEF
cpJaGgYKXrJsfS6Rd6ob5/9UfwPYZWKPaWMgndZVb0CPFCUyHPSDJfTfNLBtfMrw
QStZ8jtZDlH5dMZwvMyt37ESkxmOmThT1iFb2+mGaaRmH39+pmJR0BWa4GvsQFSu
8c00WaN7Sk8Ua3sW1cAz8TcGviqli23aMDPPwMpcaX1JFN3SxLfMRbGseX2mjXII
ZHIgeu7+9Qv/lrpEuFjeP9h/h5l0X8bF94wx5kij4Ajz66wtdOl/lAZyogHDTt8C
aIQCohLvwfKtiX5nWzEb6MRGUyAipsk5sDA3/7pdhQfGgnWI1OMik1aqoyXaUb54
LoZ+CB+YyJcEu3WdwLr8rqsRFvcdhlxOsa2qZQfGdmRr1jJV5os5EQwJux6skgOe
3hToW8vxTA+tsxQOkR9FpM9E7kV5XO+L+Z0AmfjO34nKdJAZSJURSZmxhS2Z2sIh
BRhEkamh7eT3Y4Am96XewV+P+6kcDpOINNDDrFRQvT04AzaV8Ux+N+t78D0dKS1D
JbqgGNPTqSiihZGKktKnGYvf7B2isvlVZd90hoHCmRGoL7oZlaI/5k11njEwCuOI
3LxAtW+GqxUIqIfjaE+K7RxwYVBQtpsJVwc7aeV1WRdBDHfhLFnp0URM/QkSZ0fQ
+irNZX4qW5+TFFjeq9uRo0f/SB4QZtcz9/5BiJUuKSjx1AwuY1l8CdD54jADc5A7
1Czmhd0NloOCVHrVKHuQYOlwOxotmVPDO38naxeQAcOq43XxaXHYUbjhlXUfiSub
/TyV4dBNS805ZhcXjZPkbwapC/L5X8L4fqr4rCEmf541kwP/a0mUlT1C8lVykU0S
VMnWr/aE/S6GAXyloq5tA2aS2vw9RY3rWsjOWvx4FAfey8HP3kYGh0/sSrwfDWSg
xIB+uhAT1ukMebMb6wRVDB5NEEVmF0CVO7QpS0cWRrskltkW4DfMQq3wj2atpusD
HDxdfG3ZQIT/KvpQVCxY877Hmx78Z2+olHTMfRrWqoyFKZh3Nu89P7FRepEgpqSB
M8LuDBpntgcPm0yhv8ydvR1t+JGGuBY602+JbZw9ozt9b0+WkoqPTlVBejlsDNDa
cFrQLBIrfgvRrWSJoq179FkPeX3sQFPLF6qs6EqooMYM1lV3KhZ1+J5p3PScTqvh
UbCTgTcwJn12Y+STGJptej2fsJHgiexgjJYHXKThL5DBe6+QqBbifZJ+ruarK1bv
plfaztni0Hnm2/bHZMy+RBqcpsyr4Z2ExQ+Ritm/BeoJFTklu/+yRv6xtJpTXn/5
zZT+RBsTD+KpI391L43lWz7xWZDjxzt+0B8jUx0YUbjRUoVuoZtBgfp1RhwIUsyJ
JdYVF7Ifs50GP+nRSypElN44q8D9msMxd46dIouVSjS2IC0AFyDwDKnSPFTHJWQS
0xPEm7S9XMby5u5yn7O3A8uZEVpztDGK3TQf/tWRway5EIMFLfVqcU4Wna/SbZ+b
a1l5Kw5c4Cl7LuMGFECganPzOYYMK/zwbj86ln/xCzqv1bP5SWwU67swj8q/71vH
7jCkXg35SLOk+NYzh4YxIlyR2mfmHNNd8C5skrp6CAnxjCOL2u8qZrFeQHjzIA8g
YmMCXRV4EGpwetiaS5XNvoLW0mwGjk8ADOf65RW0J3PWZWdTLDnk94DbFdQo/2sZ
5+QyPZsTtXD5FOVPI1MrQco2R6F6+Y29x1yhRigJryzEj5lROqdOLQKA//yQn53x
pC+LLWVsSUmG8peK+VpFDf7KjciL/DXrNQiJ4L8uXvZDY2rlLctORPVL2XPRiyva
q3H5rLrLAGQstWye6reULp7502E5ZuFF89aE7ff6kT4YaUVUbfAUaosbjqWTIXSg
JYObzmqdmwIClaKVRqyMiWIGG904ZrN2Q69PXuSscxeLNDavus/9RirP5A/pG2GR
y4aHY/tNAe7rgIo8mLEiZVSoDxHYnfDTnFP8tUTmTYIbKkHNjhq3u+SKSLo0MuQl
yMpn9/Zi4uTK7BN9kmWWraIsr6z+6RzbyLsiAU3Hkakkz9IRWdj80QL5V4MtXHjO
5MmotYKWGK4WXXzmldtLFF308WY9KbK289BUL2VYsba9hd/XoFfXtViC7vZs4oEB
NcALVePmZs0sfX7zYuZ2Zj+Fzg1kZ7tWr7Dm9mHOXuoCrMbbwuXSpT94znu+Lb1r
h+BYqUMtgaKDT48lG85eCFXFc7AYYEVfsFGDmu91p9LAH+tkFiMPNiqWowcPIm0Y
3cyzMWhCu/QrA+MIfmPjWMay2jgbaiUQHCyfTw0tN0sxyMvlTvp+Nb9L0E2vBut1
aNd7j0iDujS5v7CdPkN9pP/KXr4mjP3L3Z2RpsUIL98jHrksjyYP+eF4YbyE1BcJ
S0HUClv+PzenHd218ewC0Wa68QinQFABzrB4qHT7uRGOdrw6cyYebuvYqOxuwgYV
/Tg6uajEJK4kV0hcb146o0kMfj4WPXcuqctFzPc1bW0wJmmfDaI7fcc93un52rub
WZ9v8pbyO5tZ2n+65eVPpWwCiMlUI2bmYM5gYGS5BvCmhxH5Zd9LDV+/WNrZaJag
pjVQhbUxrfS/ejLVuYZgGBZXkby7ay9JIdMbTJhq5XRLdPiorIsg9MddDtGt0BXf
p4587uPgF6DhlO9GFknLGwDgv7Xgz7UrtMT52lyhoRGLMllbwZHupluK6gaEjnUb
9UVIDs5SJ0Hdl6o1qFxdZxt4fQC6Mg7HQTD2cVtnZyg3JYRpbRpM2j2awEC7aw1c
vVgr9Y0EoItBiRbMMshpTEliTDdvW+6AOhGYW6sbAE3stY+CmJTkbUR/zrwGIYcQ
J3Qo64ZbnwtsxSoKlpPGn51c1FIt39uaKWSroEkZ7vpNRW+dbb0rzA2ecy3IeM9d
5XUQq1ieBW+DAo2c+morAEmI8CVLsL/XCPPlo4oPJ6lFlychSE0thMXz5H73nnVX
yqPDvcFoi/2sJ4MofnoyrOLUTHzVvAmcd6q2RO2naxYh6Zb/p6XJcjnkiPXD6eGX
KNKxKx2nbLFtk467w+uRBVfFY7wjSUmjsEUAh9XB2C5d3Jsv+7YeBGglGIRpUbsh
F+AB0YYuM0w4SzHjIgojrqphLB3Oi2G22u/VS0DL21EUf4lhqjEleASBoMpcwq14
+w+HzOsGEqGydp0nEbaj2AvyhpanyZldrADYYjKWBGXFXGDH7Rki+NoEeYsG64gy
FtrgwlmjgnQrbN9y0ptRD41DRV6ly6GspqQJOE1RSg4mKFt/0YHz6EQyUEWWcFdB
J1TIW74uDvRUA2zZ0SQDjqL35N5wd/uznawpEQZ94f7q0EHv53oZwyQYbw2gWSup
HS/ehnWxvQg7z0ldnzU1c2TFSI34Kp9oOTJPoW/axIKoyZiLMr6Yw7B4cPqL4rtm
P294Nv5FXUUll664ZHx4yeQo3/YDn+vI2zSU8TAZDRChjRZEd/9gQG3FxN4UOurx
VCNb3isKrFkZKpT5lW3kF1eBALQ/OHdbCJHrDuWKxFUQnJvtMWZXaDF9LLLj+66N
zM98cgYIbl2PKhIqFwpr25KnYxoUtDSW2hJXcw4T4Wzqp0Dud3eFtjCNngPqT/Ne
DCaawWMuq4iYok1R4HDLmdcWAcsX4ZVQZjrf/xJGrrNa0vNxl4+qROI1dLMf+2nm
y+aBv6hmqhLITRgMLPFpEUormGlMGtDYa5iJPjY0N1Fjvc9rsMk1ii8sbEXfLY/+
DAY7iXFxTN6fwfLEbP5l3kR8BFOvUQj+HpgTVupYJMp7NeRUsQ8PXqjj8TDvG7g/
oqcmLJgoSvxtgDhbAtNY9uFDPKPrX+roiRr4eDhLc9ctxEFlyJJsu/cBlFZD/QNs
fOEgK73Gzcd0FiTqfyveIbNJf/8pD8ARbAKIU6ccYMzUVpDPHFc+UsnEYiPfNWAL
x8NGjBVz7Gjl0zzZ1TgSSCxGrKNTzj7kkEAj3c7PHJ37C6T0uM28kvTKo5CqPexl
LqmgowGqzIkK8n+Snf4g/lF6WUqhggSbefvpTnBR/KSTONj8OyeZ6vrIMpM7dGae
6rF/fENmfFVdOfOdxjljpzazYI2cIcyqEGmyVR7sKTQCkEnnbTcvqQY/UkjmQ6rr
Vb3vsIi6t7LP8OiRH2y/6HQoF/FDLk0wPDPkncARHcXicGQrJ1M0TuOhhIIY92yX
5zSqOQOIrun8c/T6CMVo3L4lMQ2gyRVv5ylLXStFZs0/H75aOgEe5KALwjB82+Ib
m3cH/J28BM9ztKKG/SwY0IfENtii2dxQ0/JOeR5WrV5/gStlghh8wr+sCV/W3LjU
5bFCMjSBd+xPT6Cj9ci3Qq9ZAyflTpcqubcpkNCgrEn6eAHxohu0bTUfHjqWSDSt
f7+eiAEBzjIK4yPgKLhRIwZ2vSrJnYdvrpiISXi2pmr8n2yJF4Jsa6CdCYZNYsjO
/OkosewN3817ODmJ374MPLTyc5P28YvepqGgVjkdHa0ixa3GNKWD61AcpeAFa9ET
IyrFyrVFSEtNb4uyYBlWyHGsQUWcrKHpJoprXJq8O9pBDBOgrXQAllQkZN6zMNvw
y6l+5adD9E3uTz0eX5oT+d5whqBuomEW/8GZYCokafVnokRThtxqilE0EgsOKSqr
JBd+kKcwvcLqE4Fkp5U4g44NQN9f4QkDKgSmaA64wkM8nv4yFACBz8GFzpxkBakj
JLT5Xyxp0AYzZuk+nF2Ab4NwnwdgWvGUyrgYBTehPodU0qrZ+pYo4OtqCqoJQHjz
IxeilUlHdIUln3XnqJw57fGflwzl7KTDZ+ZN1vMEN7ga2+nu1B1SChZNrhsRSQaC
xvcCtTyAH3daD2xz0Dwf8goLvhBWsro/HB7zG4+7Ke3luN32Xr3vysGR28u43W1A
ahnSYzQkCYWWc9zRum44UcX9wYG4SsM9liTx+WJzToAIE+QESfTrsu7O0LKux7Dg
Rvz/74SwEU0+lIvvs4QcxOj9+hSFqxYTM+693fZGMOVaBdIgpng4kq2vLPEbcNhE
Tq9JvbQVgcUscqML8lyrnRbCfEd1A+obnC4qy7bzDdsZ/YzVd2pnHk+1TVjlI0nn
rU2l0MGdsE7XkuribqAG/vgghZI0WYKQFKTehE54eFfeTfWN1uEyzHfidOPD9R7e
E5NO1ZErBoNd1vBmKqb/DCqaxQE+46QRlC39lNlMAbtXnsBqFWknTrizzDaUx6yk
FI2Olw0fVweZAQmGBn7ZgYGtrDnA67lNbjiHiBHh4O/h4PvVfW1TggcvZsEgCiGH
b1PwW+61W0NiT+7KZkmQC8Yn7991WyQRhjg920UMRxPLx92lpXZVYouQxWDofO61
CTYwkwLmbLCmPH5Zl34qgucKZJRWuhgTTvKwNws+oIQlM3p1qLPhDzGLS+n+WwRi
wyoX4Y5XIMh7gDiGNCsG31Md5abBO60eT3Zas+9+UhAmsHzB0Lzx0O7qM5ftT+dL
WNVx6u9Odzi8LFTp0FFXfOYd2UMTVIcW3wdXoZwz5bPZAdEizVIQPJgDP/GB9Boi
SZBlPJ42HbGSKpjMFbsWXjOCdbuJ0QSwQ3zFjJlrfwVMyUwjMlIauukMaF73TF+v
D3rB6pyWza3H3lGgvLqzh0G+4ItSDrKp04lU9J9WruDmx5emlWsXXNrnsv389naa
Mns+k1OritDpmeRNr6gh5tI0My57+21uq1TMIa4RRc5YJVJUkqRxvNtElgcghLTn
OInIkz+miD8wQiUmfxZk5uC1ubHrjxm1Id+aiML0RNuETbkWZpSkJjx9vpS/gHfS
QIll87xNYN/JjuIOG/QHQ/A5yobgSuPT/h1z/DG3T99IOjuattmrgQFCrxmCLr+r
nxOEWiR5KRvWkEYFzseA1DwteJkOK0vEfMblUh5h2KRGR1GNPN1HlpKRaFts5DUl
RjgRfxD+5HSR+B2eWWPxP9uWQrWtwTbySJdcgPIyjGjVgbPNdItd4D28BJFBV351
C6vWiM0oMm4cShkQBElfbhCz6ZDembj/KpT10CiU9OWE+2E+9bZbzCg3IlAvkDYx
I4GmNdRFFIiMsUTXGRjSs4/xSQWee0mj0+dKWw9T0a8YZaLZdNqFzgsqDr1DnEq5
xSjr90WNZQR+g5wrVZ35LhE2hTXT7WEXIGtXAUs99tzuqGWX65UCDgsAOaC0aMaJ
pxCLDYK2kWd2t/KtnCNO/7m2kUWTgerMAanLY7bpDVEtZFkDvDdmKDy2rNp6M8TY
yYZLsNwEBqK0r2wA1bc/3YqCOrzfSih4theky63qBF6DIvqvubsiA6VWdKHKN+PX
cWXWKpwlswGCNn+GB0af9OrIvySMzw/rte2YvppM4m4tO+mJ53vco1zbnYcuU6nv
x5ba3hN0x1Dzwkyy9ueN+iUOfWgBCBolsihsbQHdv4I82fNjN+KZiviw6uyaD3ZA
HlLpEnZ/L/DslxratgMmCvrTTyFGfQD+37rGOlLmfcx6KCNij8/astA/oPvmjyvP
t+Evd9dmdjrbwbrGLHaKd/Qbx5rH0bmFmXVo/9rUp6xaOoxRvEcnUlspK/SdsE2D
5rXe4gc4m6gRBrhcC0XCzVz77XAhNuFXAE6YCh+bt4+QiIW/tseigrL1H4FdCnoA
vRW4/tbnUUhiP6PaJA4p5qeZnY7jeVVF+aznlPHrRz4iIR6e8a0o83tr7EpH34gv
BWkmuDgywlrA8kUaDRDt4hTdT2X0g2PFtkyBH7k8tTRRsXAio1IbujREz4FXGJR4
fNTj6JvHpGFoetNC12veh18XvQeqvEsBOrU5N2U/XeWCFkC4tc8zNOOSAEZao74k
Rme6qt0Oz/tVirZHD6CN0VKhnBD8MxOW2rPMGowOo1PdQtqVqOLX8aCliThxgvk2
ZGrpwvI6wPby2ibkIc3iXxy58VaygFMVRz4VAyFHx5WlMTU/bfhdb0mnDPpnT27v
w+/ZIFOFxMN2hHcf01170gvLPrj+l3OD5qzYLZF5JMCUHhNVekQh4GOnfTFV1cWp
coGCcJsoRSKDUyuIVMEXuzMgfUpLLP9bToefWho/bHzGBYM5bhf2sorWmgbXRRpu
j6iFn3gsLYscbp4ciNc9NKE+BcgH3ckFppclYgHKcd/RZCcIsCwq5QVelTeT0Qf4
CeMWhK4+GC6hKf+o4lUy0SlN4qDNsOIwP1DroxPsW1/XF9c4fWvV10CK3SsWFH6H
Xdetd3jelqOP6SlB6SowLNFtGQchk7yNNilW30oVhoWzKva/PlkKj/SuI9vWbDNw
3Je0ezrC1zfo5JrAwIF0jVVVHwTT3fio5uL4cyjH2TkAkWfLPWEPsgORp6GRFwei
me5xFtnNZ8YycVB7lXurT1CHfDT8ziwBviofPyb2OrQinlSunA0IJsVrIdpgd171
5wk+/PmQ9kWLG3m8kz6LIgSEXoEPmGNbziO0lP+r1AtoXZ3Dxvqrn1/Ra92N3Zzh
AQvbbqhf6fzvEBvTaW9LU0lkAGW0rV9sdATUOxLiHI9fJAdGcURuubreiGieRA2w
A58uV9ZmU5NAE1QFu5f+lMmB5V6mlvKp6H9MW+fPfe5IOBNkkdOnO5ZqZK0PVAmy
15yGr57PxlduEKesQM1a1g8mcqG2StU36LD/fMMooEBP5+zzT8EfvZSi1VOtUqsU
R6J0hP5GqwXZKcPPIzPaq82l/MrGtCQUSkbYXBms+hmL30ctFw1Bd/2FCwB+315Q
3+gLkEYtFyjRWp/+0updkTNee0FfoOPD8zZy7I8yfbIvT5dDRiHfla+cHhaPq1Rd
4j3KZhEI9BEgsUp3KtMBLm+QvcPM8fYg74Df+8cFQVg2Udv7TQvRygJImdlq+G2w
nlz0yWZilj5JzY2nA2KPO6iufLCkXEjrFnjW41okEknasgTHMsbbxqHHTEZb2Qyi
p8qXybJ/D4BAv4cO4OuGsGlgAdYmM1gHjoX8stPZ4Ofvk7pgs5OvpKxu+7zP1pNU
zCg8/LVw/49iLV1IXyNdYsRMTzfRdfSXRSNV8swHaRHnleOPx0+KpZcn99PftWXJ
206YS7QpsjhSusiXZhSpWWfMNw6DdFdAWIapNC1PfHUhY8Rp6j9/7W/fBivmy+G2
CTZaBU0uWO8onmrqqZ/5fFaBui8J4EmTTddYrMXYWi9BLGR8vKKPOEAu9h4bru1A
6Dz3atkfY7NfoVdIMySsJHxkVwwlXqisXkyKu2mpkFBDQvQZ7sf24xmuYEK9lBlY
vGPNvPfGS17gudT3AfINZmwbB7GVelEAXdQYIUUS2npqT+VVCU7LVGwX3ev9wapC
zQlzQDxgU5krJrOMBsZZDrVrIng8Ianj7t1TAAPVXkz/TLvNqpyPK7jofFIDJJzD
4f8Yxfon7L8lraDvlMbkLdXWJ00jr1uy1n7QcOhKzWEFMXmEFoVlp6KvSTCD1dIQ
4nmTHaonnJjZhGkQ4c3MtAG4/KRxE9BFitGVQVggBw2HafIAGTpjN5pYIDmUcfIq
bibSwhx0fmRpD53U+meVP+2Nx/g0L17250pkQLW/ZImHkQcE/wK72yQZ3QLyN4cl
ZW67Y2XID8mzxYVXHdmlHKCXY9NBRcevPpBCasGXwINR9KDxpXfF2CbdpJWAwY5a
bUtrMzybTqsb016vMf4XwYF832ck92ESx09vz8IAYWlZP6sGir6+XM92BjWQy/c9
e/TWyxdAsCDvBaAdDKRuaV9bOcIfXGRIUhrR0zVkdfMoOfORSgBs2ju7ZxcQzTxF
qJjaI0aXfeS+1i26u3L+1WFEfiF09rpGUHxMGMgo6CZcji7Zq6zbBc8BJx8mAEHD
vtRGGuFkwLe+NHfxjyb1TbL1PHqKJFI3E8+zDsYRHWglsTrnu5qjSRbtNDyUi2mJ
R5P7oSQaQuj8jhMRbsOGX/j++6TmVJ4xjqMry3BUL+iEJVdvgr4K7G/pxgCLKCU4
W6BQiD8iZFaOtWjE5sQf1Uh0x8ijvIbumh1oObxy1cRDabkoKT5tjDq8uBQlA5K8
E+w2ageBXpRSgEHnZzDwDAsLvF6y6P4NBg1lcBksf0lKbWQoHURMtvnCkFpDWO3I
l8ljEVMsTzXxQcKoEdFQ9zVcctHV1r0SMZd/PPyD3rFWXr3Yi8TmGgym8xbMbZIq
NUzUv8sFlWstEZxe9fHUz5KYY4SFa2hsoFIb1FBTrGLchQB6LAvdO8mH68Zk97//
NtDt9h4tTVCS9hhiUAfHQLHqupdovn9mnt1p7zokKqqYCfOPCcUoXghM53sCcWex
rUfFsf9eXB329vUfTEExbHtYicmNaMWGK42N5c/sa1u3/SZOjfvXqNVXi50+VXxK
BV/LFdTGvXs8sqcvwWTNuHMyOQnrWVzgusQYMkjg5DkOrGs5it/yjW4NOsjhl97y
cMr928c41Q1jtHGcD2DkzOmMRhmFCTYoVqnenaG+G74VVfjP6DMIhZu8g3p1r6Dy
6nGwTGL3mfVHl/yUYb1D8enuZFnqKBU2+cr4rewCQ/wpvS4ApCPOFDWPrQowHd9x
yugNX52LXRaHfCTb05bbYbR6OOn+5y6wo2vgpbNgJCLmJKfw9W0FBZurMYtzyr+r
O9QhrTExHIgwPMwgLGSCDSI/hly+4g7+/8AQCka/Gw0UjfgaroeAJchq7nMBlDDW
mBNvReFa8BlD/XHbvdc8b7Baze+nJ+6/2i0pa3kQPavezJrNIm5f01nmSDv+wifB
uu869lNRe7mLLMJ/cbF5+lPgAYWL2hw3V8V68NoPEccEr9krvy46F0NN7PQ/lIse
4J8LO/wY4ZnYiqhDFMac09JYLWMI2WNH5tbZs6eQZL0xmamFsICEwPVyAYyh4wKP
l+4OubjgRAn7OiNOV3eJbyZ+dpKQeRy64jSm7gXTG+fcROUvO7pWn06uXJ6gB8jY
juuUyXvFWG2AmsINpweJ7IPAthU5HZ13x3uYpjc8ZA+NOel7yaGzSjaiqdNXfM4s
6iXiH/T8G6MzMICNP3CmI+6VxSRxfyHFKSMEo6I7eMHgrwDes/zygwbLIdbCsneK
oaZ7xP+dEQFWt8nREBEWVrWOCZk7ISxHUq+A+eQjO3klp3FZ/EmQPDIjDmZRqoG7
hfN5bFzUxY+cb6K6e0x7K1UZl6pjzrOrXvZCsN17Nmq61LpCANjP9aeA1u9cPQJj
wlc1LjMkJbFK38QtxjcVomKhrTGSoLaiZUp35kR0o4GDk8GuYDVRPoYTHtvMLEea
wWwbnie6Hq8qZfyLA8ZZmrLrrxCG9yAPC+zMvM2QS5oFzFEApseYhyoCFcnvt6sm
GoXVaD/U3tCR8Y0qOWuwW+mdyWePvfcEz5GKjWpJ/mJUU7bW48RdIIDqlZS+C52J
2wsydsvCLkSSZOUT/3V/QdbYXMu+q0XRSCkHsc0SAbMDIryjF7jL/m2gDSsGGqML
p8lUlg+fNd5tskaZVUHNTZgva87lCZH8IbYjgQ8P3yasliPZrmgx2bMpqfJG9vcD
FIXKk8NqO5aCKRWJFTx68yVzIfiZRiIdXL2RIj2m8oV33mUeRTdn/tj3Qtw8YWg4
UfQYaJfNJvhckcFSYVTBUfVMGZ/i6ykoMOQKnTtVgamLE4r7BYW1I47Bvqz+zqAn
4qfdo0oNuPOND0AB/0ama5n5cfyOOv33SVQQfbozG8QqrFq508JB7MvZ12I1h3nb
vSSPQABPFNW/eEJMkLTcajmPqBrWdyuzYx5L9NBEGVHYmXz6VGCVDrK91LvgJZFe
qmt/tnzpJ35WZ1nCHm8wxbVxZWjmCfotLnWf4HhVFmjCZ5nxELFs+ZZZmBPoJQ9q
6BnMOvKrRsYxymR+SW5f3xwyzejn/EdbbH+AENJZ2mBDyYCjpnQHUXYHdfS9JtdQ
PwQQ3U76JvKA98724Xe+0ruwmaNN3iLSfo10mpQgc8RoV7IxqFMifQJ8uWgrPw4t
XrvSHzecJd8OjwvGLcLVSdE3nkW7/HZtEyHiqTlAUrDRZtPViM6deTD3Vd2q1vpF
ekKXJ+lCIidHzYSFH2HoDYhqIh3x+ofgbguRpOvFBkhyQmqiidJ2Jxww2HvvjHvl
8Tte8q2QhmJMJ+ZxhAUjVrxUn3PiGIQx/ho2e+nKB2H11U3V8eS6HPCXlINUWGMa
vaekJSm4ZwOEXS3E6DF0Z5esQBOaG8PPxxM/9AVcJo6ZrMKn0Py2wUN4eZD8nQ2j
/8E8PorK39vM/BGIWaFq0X+JhBlU0eyryVrWXrEQMD9ry42pO8SOdoJW6yWPLphC
Dd+3AW2z1ySIj2sUHwqtuG/maUW86AhPSR8xRzYhV7E78EMuVLQe528KP/iXsV6C
33Wcqs/lnBr1+JJUUf659GkGIkck+43ZIQV8uKqEH42HD+Ts9kMsu0UtJNutt+1U
CVYPL043dD3ofxtaWZtS9qyl5g6ehW/Ei9clDP2DOY0czP6vir6Niq1gbUYTyqFK
Adn28Ocone0YQGQzVzfSXeFuqKEgprmDNHmhTCpngKQFThz3afeMmY5eE+LxBQZ8
E2eFkjjejuhJGAuptJxGYlWXlaKS76JsV1YTzSOPErAHKBxlstAi1gUgHxh7K7q5
gu19kZX598V/yb82rx/b0/j8BW9e6rLxt7IC1L+7lbNSgLIlwhdVR5yoAm2J9DjZ
i2w7AWANqL0uy7MyWU0b07I4heQfSNvV7zknq9MPmfG9V+aooczXxYCMfOLR0Kkr
bImYSWgkw0tna3E0CZZ03C1RC9Bh9mb7a5yfk15FPaqIjt86CYOw40yDgALSFD7W
xE45qmBdkf385DmlbVw358MzzHGj36T3QyIBY+YqN/CZb1/iktOSMsLEa7vSI/FX
/DYa4c4g1yRvB7/q06huGhi3FnKJY+pE16srHy+DKCPe6kC/lnB77onoHxjmviU3
CU3rYKBq198mOGuPZ/Sb6kyt5hDVWQNIy0lXBTbkn/qaNVC7RVO7ToGUiLrN4PHH
iOvnZNQsTvPESMzd05L+e4nI7DT5pKBkUY6D/eFtZqdrnMDmaJ1iPYI+7KMf8JH/
1kUSzW8XVn1yT3O03Np2f8n1XhgGlGx1nqe8UGmtXnhNtX13C/fhy3GquE6mSWSQ
JVoHLNxy13wGuRB90EKiv/55CkJLPxr/YfljSG4uVBMwWkXWfy7ARJ/naEZQbOLa
8RocEo5SiYN7J6+d5As9MqGunp6rdD2OWkUlsKWXuzRsWbzKiOnYR4nl2VXnWtko
6cGSKijjeNVo+W9486uO+sF9iTgIvSgU60fBLfwiKFYrqjF6CyjVhT1KSvvj5NjD
V2nFnkgNTRc1KDbdsS4N87rzdBYZb3OzUtEbFvXEEg2HMCpfvkCmcPH3tUC1ofZl
QxQTZK2vS8XbiHvXveNB2aV0GaexqgJI/eGGDo+oT/NpqzqICQ8e1aItMBN9pT7u
taG0zZBcIZjFtS86/iC9+ddXx7FHrdeW/HT7jOtWpgjVgbRxjD67ezqpzaDxKE8W
E6eBaSvdzczDpVnVvFRRhGXQajdvPJvojM3y5JSsQEgvv6m9bjWFSew7zeQeVYui
aRXdS60t1un4WgPMZq/B95m+PID5rxrVqbZ9YhNMpixp5paG6mmfgdJH1AV4MPsB
NodRqTXAPiplPAD0Jw+Zly6kqEGcXoNxboZRqIAxp2fD32EhaoI2I9GuqNGDBzy2
E0NRZr3I1eDguzaOvJCy3N1ctEKnYmLglI9+mSzgrCgsa70KU9IoTJ33+SMX5BTO
bNmz6txUdwD6XXx+jwz/mcWgA4qcHqAdtpWej/m6rH58hk+p6Q5LzR8dozkz9pJh
kDwy+CwilfwRfAXrbjSQWWxyDAubQPNfeYWmCu0KnrpbyCGgV5ghukJmQik9a43v
7vkYkZ3CQXu26XAemqumc7/lw7tgA4o7JfwlyhRwZrlGvjt3wWbPYCenws6MtP6M
i7wn0qTqPk6S/DGhYr8uKGWNdtx18XiS5H3FGFae7Hp2aDmmTzg6BTGdlYDrL2EW
Z9iQKP6aW7q1Ms7B75wWdc0IfynzTdbsFC5iWcbKsUpz1yQnOQ/aexkqGSJ2i9qz
xDmERH5n7XQbaWqiYSJLfihGiSkpn0Uq8PzuLEeN5q45bCtYTVOAYf3xtXs5vdUE
hThDbzUjp7PuW2M/2BQZLgddSl58q/u635Va9tfsXPqb/6789pbBqVSWG8WGerP0
qFWORMdgwc3SnqoqiFqPuxqmDnFsbF7flQ2jSUYS+a4vFStB6OJ0qGsLe1vnL6Wz
PogJMpjC6hS1Sio7Ew0cnNqIEok9JHda+z3oW1czgYoxIpQmzDMLOU/A1tBRScRr
OAhpuv3jmMxrs2papJp9KbXdRxlafBhI20A0PgCitidR1JURUh1SlbrMw53w1o8l
OdjCCcn+bsZDtH4WovyQRM/NDIeFdwN6uvjtCWVhD8h2U2yZWW78yrHK5ve7y35M
JL8auabw6eehlr28WY0JmSR7KmR1hI6SfqBd4zQeqnf2gW/7/OcGS2NFRlabn7qX
jYPe5qohKVcgkZSFKkMhTHnUEB4OaapeP2OIcSZ0GM6dU+zu8Swd+eHafZsG/86Y
TbHZy88Yylc5pBCzJrlN98wiw3uHnT9oT4qHpMpCB+wFjnz90xbeHIL+YPlEW3OK
Nhv5M6FilwYYKJ5xic8s3JiEk8lzoHjvmCRsBbPDw0NENCBMCgMVgBjR19UIxtBo
3GxGWgnr1LeaLmt6Q/oLySvIHxp5skkg22m0LbKzNN8fg2luz72a6+5WgYstWxwZ
AdDUfmSgAD50gYZnqiYyt8/tqsokFL/Uye7XjgflXn8JZfVOtfY2rvXvj6Vs9DnU
CKBnYap/bS6B5d6FWjx6WqFKln7vNnWnoehvqYpvYv4r5tTk760Uo6o6A8h8np8n
BY6LJpO+ALpl0afCpxH7r6M1wyzSMsBBCgT7cxtbKSWtSfTih/NUlL0y1XDIelTI
/ujEkUXH1qaVdL1blxnDvmbFuTeT3dPWaxciVRmnKMJbuAj/ebJyWKYbvZ2yzCeP
QhkKmk+rmenI79bE4B8DfvJtL6foJy34QXdKjdg9rJYsFpgatH+iVVGeYWnyrff2
WwIwZoPPWNUvVvjhI6sICEQ3Ffuy8C+ptPT46xywUGN3lorAHA9x3AdgYR5+ux+0
zpk6GQro2SLEKBD9uONuTyXXUEN6Sb2xWI+1wGKoamYTqxwdmS4WT9g38CI0MANW
r3PiKMA98U8RxQEID+A4dxS6hrHzCVdDpXkO80fs00Hf1SRhIfxMXz1jiivN7ukC
ki28vdfa5nP50Ok68PhpvGVp53AfJI0OF6XDdXiN0dKgFJcw1kYJWN+mjSWVutJ0
NqF9JMekD4jB5F6Go+Wuxd+lwZHqEj2yeP34Pj/h3QZ1L56h4zp1y0HOOYsBFIhY
N+lXgHmYZXsYy9P94U7dJ3kU8D5saeXjwHiCwQj9/nCB5p05lcGvhKZbGM1jL2By
/ehOrz5xhwckdGbWUh1g8cGI9iQYdTjp8z/vXpJKVT9ZL6H/geHy7HjlvGPm6Ckz
kd7OsK/iy2QVACc021rvYvfPRHPZXfxqYX1BIXRxv0S7hJgtTyaXwjUDRwrrqorD
KkJ1bbAIM2YqnGLogTfqsV5M1et6D8kXH5OsFhg59GNmqNzQS/XqlxHNE5jYOlUC
AaxmR4Ju548DH/UuLb3N0DVsngRtgGHvnrOMfTqF4p0gpeXvBjhMHz4vPJBZZAVX
PioBCliIP9shOIQAvXW2vcCOkd7Rti5umqGn9cDXpETHTN5S4Im0Go6NppO4OWi0
kWdFzucNyNgy1t2ybepLdyN+9ReqIVtWNdpKs792oIhshEHXp1dlDQAUw6j/DaDP
WQ35LtYGNay/wWuxiCed+HtXEe4gvCd/Z89lMpmSali0VABBQWJQZGCxHmpH8BSH
1dpp18aR2ZNaSBMYqf7LHVlAoFmK6aP7QGACsBpGwnv4++tt9iMHb3U80d5BxqDD
+dDkDo4Kf34mApVQ1oCClP/LhVnrCHHhNBiuON4suQDznfQuAFbtEi4uK6ML8yGA
xnHJmZ7+nJbiLBWip5IDSf8g5wYmPzEYfaNxWRizfbddqb36w0rx79g0yy226qjk
ZqL/e75lHK79pfuk6ZV0tU24g2zUfRFEH367WRY2JJ8s3gfS3I3jYI7NpCLNvwy+
GnduDZP7/1qF6OeOxiDMPY9J6w5SweuuNvwDAvKBBwSVaxYHFDqiBfiLRirAruvu
ubLlOjMJnJLHTbZm8+mDHKA74ODliq7F9DbQg6lIFJ3Yps4qnHMN/jFxVunN7ILW
Fba56DHxR9Xbf67EdD7ZhyToKqeho/DWH2eihCMbpwSE4XlsW/GGqoUU58YlUbjN
CSV/YEs+9pGbHI/MaZyd+24deKF3f+lC+zhv+Co2Y9uaco6muXos8GB9r3ZdR/Y1
uggHvm2yRu+QGWkpjkv2PKFmudP9diYhDHF2crmgp3VOfJ6Lugt3oUWUfa+qTrmK
x0iu/CM3VyeeO5E3wor7ZYNE/OsCW/zBGIG07EKuTY3RRjP+Fv4ppxg1xczRIJAr
6wFL+vyZD4XdYKxjjwibzAZJnbGpsFs0O9SiyHnJZj7fZPA2lppjYCWmfAAFCVc6
frgtHRXDiDD3AnOw7rmHHKgfjV/tsJuJUCWIBx+/KNw1RUocoLBmUDmEt2qXJsgB
NJOZ2p+Vno3D9WeUXjMZm/DHBTKox4vJ3X4keKGC/XFP9tjPc4tqLpAlzC/G292L
PJnRBvu+o/zdF5Iiex9tDM8nvbh1iaKC7yrHuMSO2kHweGbynhd1NQVy3rc1iI7P
aNpKaMbhkTOANP2niWRB65mzoLZCJLdqGEPtZzbXwuu9yeYSSRRv8oKTyaFQr0wx
Kd2uXRVH9O75I97NDBHiFlCMbyRSmSLblQNZig/ojpPO/XZTHRN584OuXA8zaLmZ
YoQrnUc+8bvlTn/IMAzJAxDo2SdHgvjEUb4xd88gCauzG5iTeCuIvnUhK2gBoBeJ
Ai/tRvEHftpRdOAFNNzVkHYX37lbjpIY7BpkGc4loke3OCTdSyoIFNaTxUUa0skd
KRAcz8hblpcPz62DpE0ROSU1CQOzYwKrLXpzzvT+i8TgpteetGHKV7lowuUTJ9c7
UtAWwJDTL/jOgcc37wbuHiPZ0z8cBW1Xa38uR0GPgww+XXBWVYdQYrSDSf+DFi4A
rWBdFe9JEZmX2Dgd0S4Sbr5UriXduzLdmdbt9J9fGVsGkyYO2XDqDbC0dHpy8DfL
xunzqttE6y/ekCysj/wf/pZqPkzwz3znwLTRhYtTOQj0or+VhvtVmB+j9lQZ3s7J
pToITaKOsoH7EkvqoYl8rNzqLGuMf9z7aLYBit6nZev91vd9HDVieK6RKMEICKtj
Z+UBp+fN/0g+dSxRDBrZrjXOXa7JFkuJiZn89dctss4X+2lckGM7WEpzKC9PuTW0
ugp6H+iXophHezC2odUiwEACSyjE7x5hshZU3yqj9F6QyfNjn0ETPo1LC54k9b6Y
BPN5yF1ObGzRUXYWcPwWeC1qcdNbjH9Ehwdv1+/vJLX33doRkW9/AS5vGNIaLmHH
uNprC+o68WV6mc5rDkDvKR9S76ryCTZ2IQDzA5NYuDHUVHwd/Wh7Hh480i6G+WaR
W4dF/hMOnDzalgJFXRSVsMJZn2XMaOo3JvDDdi223LOVmHMi3QkTtDSG21h1SZ0K
PkW5SvdpIu6/v7QFUNdEQpFnccl1zlvIHfIUAcaQkdZSfwtMkyA/kwrNFadSNoSf
gjoRPE1qILq8lKgdlSKMdmOiAhR+vp5xE1jNr4rFSDKY5DqJteUaquolquKQQuJT
noGRzvrPwzbaMeu9Og8EKh2SrdOmDLmazxnib/R3FRFv0OU6My9JQibAZScbXAv6
VITwPZIlURb7sQ2MUm9Lvw28ip8jsrVzdhrhWAropZBWJnBh/icj9Q3YSxr2gqSl
5cbEGPhwSaYIr2KMh45VCNf8gqNaFuUJ7x+ACvzWJqpk8lMw+eqUl8iXpxH5L1CY
aq7q+xWBfHvCzE4S+ZWnXdM32MIBTBSjqhN+Ia+sBxLFOmN5FAGpG5xJWdrEhn9C
46qS+QHQzy+AZEpkNDZ4MdPlRtP6Nba99IEkSoS7XevPKmpnXQDhrhJkOQ+p1IsY
ayWe8h+d8Ecdn3RfN7oU4mlgk7wtSZh4M8MElh9cUC0RtoX+od4ETRhqPUBQBNQl
5y0RQyHbeVhTkqwQYzwdR9dpt9lmF3ws1p1VdlONNVOYSRMNOm6LpKH9KsebJdVi
MjIYJvLtDz5ZqA04AIvGXJdA/vMrqzjBQhhGmfG265YsMvweppPm9OYjYSDNYrPv
gWubfcKlWwfFE7saI0a0venHgQIYgRJE7vSpmlSu3OZ7ch+WCJ4tGD6wOYF9WFG5
VTRvhXFnPtBRcjEhKjo0k7RjfGQsxa5SfYAiGPGfAKZpZfJ91D/bI806GPX4IrkY
52dD5lfFlnHSmfLW/sdGjER9jIKXN4RvrsFoTkLlkxhOu6l2ObttDuc2p/ov4wqX
YnQaP9jheF/1iXcHhdH+0L2BoPSdwzp0U1pOjJr5ZXVGQxs1Lc3FCZyooaFx/si2
Mau6p99r9bwwu/VWGAy0F0OXUZ/8J+Tz283jZwP6nS/thcGeW184/IYsm12n2E9c
axPxx6KLE8aVmkzNOb+jB57UcRlCJ5izOpEAGO9fM0QkOi5M1+Jd7dmWrq8N1fUM
XAlHEblPbyP+meAZEktBjaQ/KY8VIf1CxgxudPFDM94o63/oHZGCXBSEpVIOWIBU
noiCTpiG6LFzoRkSzx9nUkTBbGdFZEJGq2nYqUJzvE77wwthSmasF7d/svMs94sD
SLSkDSBhOBbpUEnT5T287kl3cCzQ7T9LGmqILxQonmCqY1tiIVVYHmRct4ZIDoMr
QShmXIwDL7/86Sv539da05LT2l0wXbzwpepsB6XnXdkct+2Lz5FHU/rexPzBnY9j
2GZ9yIEIE6hnIvRKq3Nt8R4UPPxJawzce6lzS76xpXeh2dfEAE9pI4BAtVPrMOXV
vAGmKwqDLdoMgUnBZf0t+NxDh40wFFN7gT1tKqjUOT9kfz+9l0Kigu4b5nURsw1z
FazbLqmf7E4Bvxi5fzixJwa5Sgo3BRZe1NFefFEgkhGZ2nbDDmdkkzKXMUjeomC7
xQyn52kJCJGqWh2PIU9dt9VczsUDNzW6NwKUdYzflZ+6JyvFx8jFG+X5DhsOcQSW
U61SE9w8bWNC6ut9DFUEBuXsVFHoW4mla4KRywX47yqCQJltQHBFvBdRL7XLO+QQ
6ohsyt+4050va2R8k5skfhetplXf5MeA5DsZYI+x1w69plZOgeA/XjIliNKkoBB1
sV+Utscudg8X9MVyGu2eMZKt4dMTkpiSCK3X1cSWNgrRtBKCJMMNXSkfKoiGdi7D
iM9YbeGCu8HrkjSfwaaDIKySFrZ552uspMnedGUyFLLCyc1hNsJxXY44E5km5qjT
M79PvVW8vb6YWvRsux+KB/0vI7bI7m7ApPx1mc10vAOmIcHDpd6eStbDYQq27sd9
mnMhFsDs5oTPdw/C+QvRakzI/Q3Ifx8NAGud5g+xhLdrbQ6rGkap5zWnwz9tIimM
64Ih06uUe6uTlu4lNX6UrTiWbLJ2FHBPe2emPkcayz0W6TCwa2as1h39hOqkgmEB
8m3eX4FC5vB4p4yZ+GCqmz1KTY0U6hrVRl8QhrGrtRxwr7Zhj4wW2+yl0+mgqmm/
HYOe45DVfA0xmTQj4Sq786OQGV10xCCH43pW0QBtjyg23SzgH4V0Q9Ob20VxaMv9
hVUUR9axVoR4wejoTOM7KbAbhk6ROhGniv7uE5BDNTZ4gV2W0qD5aK3GLOJQtbc6
RHYwDlLcTgm+/oyDvwwr1LlkJPFSvSCwPBf2mua9517F5Q19zikg24Jj8hJ99nYp
q1kK+Ic7EyAN8cCUKNTlwh2tnKbU7tQ5YFsRBMJp7alb0pquv+CJQZqxgaQ3Iz4X
nsKyoTYi9nSLh1EAArC4dUjrWF32+PxbaZQmPCo/PhUtnydBMF6p5zHGXpx0NFcm
0CWEDOuuLec0ZtvqSTsID0ndChJv/h0kIWJvruE6KLQkGh5/VlqLiRId6EwoNdec
ZjjiQhHPJ4O5cd+TY9h8zYg0CIdstoZ6PDv6tIAVgaYl1G51YYfQOjH7Md5GDQ8p
1xsv5FdaXAgPPNbky63oo/zk3IiODpAxQLfggQk7xe6KJGXvAJDBxRdXWzFhKR8Q
cMmIsVfscWxRYqBFdP3Tf4/boCA0sdAwUqov3W33TPDR4QUH3exX8fbKijYd6fh+
3gSZsPQ69MmrCrfsWVt29Lou4Cd4CB8B6GlUv4WMWMli9lCz5lIH64yS4sCG3NZk
AyyqEVZgFs53mZsUEuH7quWCmPZDs8NtV9lDThCwomBAculfC6/vdzLP/MuKnoCD
Yvz19n0/tHRIyA0yXwFB0mdm1XoD43M/y8N2X7WY+6U4dQJCkFh1mYJZICVLaGBn
QGMj25/VWq6r8joe4hdpLQV+/mFJDlFe5dKPLRBQJ4ucQAx7DvX3TOKeS/qXmgA4
dNibepGetbD4G3JN8bXIx3cews1ThzdjBRvqog1h1B2i+HJnYAN8Ftk6fsvWtUmo
ydnThjVg3G9QG8DqyykOZ88mz3ByFooxeQklHBfp6kaodGiXShRvFmS7SHTM9kmR
ldeLcpFqKzGDnlWCQSqvp71nnn3YMDVjwkFNw+AI/KSqz5EYskh/PFzDpMtTvunY
NmVKWYbLYOK9Iz0z6FTokdKTPD7e9jKtSnciRIV/c+yc2LagUYqA1pXPwDODr9fD
/SXmHqiqHviGSclZCsKqjy1B/JK3Wkk8w9Azl0qbns6aKvPYzKm9SUwVihHyGEsH
ToWvreKQmIXvpPz33V1+k1Khmihe957RheljIXIo4yS+VowJQ7GdL4v847UkUMVk
cqKbdSWmRQ2HVnf3/IzBf1Ofu9tV2H6wxo6uU2OkYRFy1hb3JtGfmiFx7WMqsoOr
JykuzurIkCC2SFu16G20edLAjAxhsVvKJbOXG8VpnPOPbxZjBKGuvit0D5LB68KR
j6lqXvLZK3ulL7iOVpPx/p2JX+OykbFEIEuEqMoI0JHvtuhkakCjxAXf4ayfa8s/
vTLJV15LqnFywAwl5GWW3k3l1FNoyZ4/RK72Xm0ejS6lyoqme6dr41lIrAbtaSVK
JlDeLgoB+zrw0r8dR9fl0WhQPCwy5dvBxvtYb9LPMp2r4LbNmv+wuSyj7pB3p1H1
YqUp1F3N9iQlYtYaXMQ59pgQuh+YeKGs5o8GjeI1fXDeqMKn7OAGv4z+1+xRb3Gn
GnxR1Hv1l58O+GYrFjMV/rOKoX7iuhtDCt5DFuPA/fAq4d8ywoxI5oXQSTYpM0+e
87RKaudUbkkgMBEyOPEtA+p1QKYs8nHl8CJqdkFzrp/aiflGQEdExZkkFolJBbG2
gz7xwbKrTQxxNnDki8aOIBV8TCIg+wXSM4eMkE0/D+2fO9O2ZFNePNLxpa3a7c+h
LIsD/ixu7lccIopkAWtmxPI1lEROWiX3zugDS4yBp55fqxM+CES/1+oL1L/I/8ev
EOuxH51nCGzPMkGj8p/aAyqFCHs72d0H5DfNqOCBO1ODRHMb9IQ7lqv6x2w5x1cg
O/RcLPSVKMz4JQE2qe9LU7yTwCSuaZSFUL8+u0gXc9O7brT3yoRN2oby+V0EF6Kd
7j4lNki3VZ9o1nqYW1b9XZ5Np4q/Mx/+EXBp+VwKFKGdm8kXCIlLfN1iDLAthGIL
M4DS5CZhI9MmipGKLxVgboxqaw8sdrNkUuZkp0Mj+jhtkMPEg9NOxocPAGS51RPv
EHtODBNeD/Hjy7PEVSziBI6cmQfWEZJIW29z+AqVM6oxl8FrJdty80Z8/11Ft6cA
KsgIJer8uKR+om+K8kOiy3T0vwniFp5QvSIds5QKUfmbDEursscttlg/l8ch9drX
kPtKEtxMrHMAx10djz5V6v/uhtYDRALLv6DwREY/dMTJchel8f1fby2EXzcQ8YG3
mS9O3tkjN7E5gkmKu5eAYA/Es77OdNo2tCPlG/Pb8/dXyHYbHYjC+RbBp3t181k+
tCPd8OPM7iM6pWneQECFqijPm5smJKp4pGKSBMYGIM1xidp9vx3NCBamVLmOzIFg
uDcWil9ZiQatjIrP8Vb38CUYW5PIR/+GYVkebdd6AznzGP1TcrayfniBIrpGD7yB
lY95i2thpWg/+l9sG2l+2pxvPt2c0k5XD6nKAatXw/3wcgxSWWdSV6ammEq5i43U
Gi/QvbFym8KkqcG4jHH5z4SL63hNdZVJYhkAGhal9iERRjxQNDxQV1s1EX/4dYsR
G1TVJ4GJLMhTjVaaGzaJLeD2gPjz59rtn2+w8Ze7iQh+Az8eolbtRC6fI1xkZ2mO
TBWAvwg8qfx3r9yxEVDs4x9Gz7v6KEO37zJDVvhjmErIUNmG6Kl+ot4cb7FGJdR8
xE9tZE2G/zHYnqQdH4/APpIcqeLxd1SBL12biqqocoTN+B9qQJelvEvxljhOZHHJ
LYsood/bzhafa63Cnwu//bqjSepJ/IJja35xfIzp3ToOhmUkrce80Foa014W5cs0
YghgNOOYmrZhdDKoQfaRG3N07wIeKjEDOPp4ZjyJ4J8ZhLs5gFtyIofPKaXGvgCA
Q/mratcud/lSCeCKQmBmrogPtTMilfqRzVhyO4G1f3Y=

`pragma protect end_protected
