// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
IeOdTG7n/G94GG8bYnWhV/d1lW+enBuNiN/BE8pWeEKfwVgl0728IxuCDBtfrRWk
Glll0TawYiBF/XFo7zO8YI++N4Gc7z4ZZ2aK1Tzyipd6nVmogYlufEuRExYjLBsp
PUmMN5KCbLABLPxmRZTCXhqc0DFZG1iGRps90YazRQQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5312 )
`pragma protect data_block
UL9EpozCi9kuHjDKWV8eNRboVKx8eCn4sDfB48CdTgfRJ5JzTSaoK5zpUyMPsg5o
4+rwIlTV+ra/BGlChxoemd3kDJ8xZaS5Qh16kTcFNpYfHN1t+J+SDtlD+hhKAwRc
8OFBqQoLYxCTp3N72BwRkRCAhvy99VPtsizLC0CSStuNJoJJ9uuj+jpL66Cx8rBj
LL53g5gYwRPL50wZYUa/61V1CEA/y33FiL0OFqi23eU/swy/fQQ8Mu/Mv/vhE7n3
EVcPWh7u/XRlj6WBug0f0ZKZ1sxMQrzJb15GZKG/1AC2n0ietasaO/RKqw9cYAqp
Fh6FokiB+N8XXV4fQO+ko82TSO96ASUFQUBavHSQQiUlFGd3NHVly9peJE3FT6wO
j44wkKpbpgf+ZGaaPd7gG6oTSACGIkdhrYfAj2QaHiYiIMe0pAjoLiKFXtiRJHZ8
xTgOcdgTfulQpl8BNus2zqFZTgDlj97bSGi5lvRq8Nqu9tcbEDVTEIQc6TAg988L
9RxiY+pEbA/dHOHM39Qy9KK9ETM7B1YEv2X+8KAu9tErgjDfrczuMQlzMe7ovxui
j8rMYohepLBIh+NUbYcFYTmujm5zGrE2j8SHP1tl2GAO5ZVuBU8k09n+e3vPchWH
TTDFc4nQp9CHgXtz364K8cJZuwEjk/lQDASxWRG8Hi/+mBklW+c/3GOJxdT790wJ
Wb3GkcEOXvmymTVWB8UI4JU3yrOqeTtIHa+1fyzyeXceFzCgtFjBHlfHPWIeE/qL
k8bi/0JCly0uA5gUY5ldJAnOnORYtqkzmOYyFKCiJQhJch2XO4iNm4fK10QV6tKU
xDGc15CYufd0tQR5stcIO8z+AwrZ+L3FcjxIcJ3elnK4Ll4BP2nLVbQQShrogvy0
Bq5b5Uu01xoB5hfegLUFdJvJezETs4FahO8Ypk8/k3wsykOs6UD/RCvRRp7q44IN
QjfSQbqL+/UhQo2fP2Qg6bBd7QrGuVoJ2Gg0h9Rhx8lmEBmC/ZY9L65VXtt3m65T
oycAoDcrkuGRELsYq+7qij5LOe+in9Q6Q9G46eS12jeteT2SwdiOiqnbBmDJsfKk
B/4Z9L4W1+7xFnbnvTQzTXmf2ooQ8z5UnuBCCGMWzaFJJDZi4B2qokcGxFRl197D
BD6kIjLKfGfacDnWKgPWrPKj/arbbfiiB4gygmG3AjjcBlCyEb4866WHcuC2+Gv5
GCjStoQnVQw4ERnMFOyN8Vvxc6i+JHytwgcJsM4xhn1Mf1y/gyiySpKhbFepKjSR
lcno6BYGyGRUePgkJ5OOUVHy4Buc4apLEsieY01+NO5hf+5Gi5KoP/Ol87qMWvge
iJ8t0r0DVfzObgq0C5jF4vheaFakiMkfRdvvhoc9WNUp046cOLczKDP3Y8I5kt4b
unSRzu+KFmcv8F+xxT5zeN3ybuHpD3hca9TCoTGvkqYGBQLZ7spsmJ4iJ3lrRHiL
ZsJANEcjacVPiu4I5RoDuz8P8nuSgZqiuZaMzG2rD5QBjNcYI4xO+8p2erOquniq
cKyievCNHObUS6vU2R2tPPJG0LC5DJ6KVLVyuAZLhpSVvTkg1FWaDmToea6JBO5Z
HVjnwMs/OnJDeDCPJMg1u0AwImHU9wjYbbpkb0GOIXhFJcPE7QNlPUHObVnIE6YJ
+/3OTrG9UEbv6Pt4uEPsm/IAwQa775GTKr6Zum3e0xI1SNnSj4GLWzo/w7awej3s
oDl1FmeiUpQi9fxhEGbfT1UA82LMWr4UgEP1D7eyGiAR1x4Ru2ejBHb9AThMvgW2
Tvfkxv3vWNkNmOPxgGBiUSQKAMAUvQxE8oXyx/3J47eSPC3K3SKDRryUHdcQOpco
Y0Cwe3/ZYLjhSiuFCprh/g/dl86Mt9auQgwG0aEmj5dRHBASLKFHJnfZ7qh+iZRv
XZkal2HMgdTt9fCqMr6Qqyuyu4rMI63DfU+d4PVksURl+KJ4cZ49wfFlp1mL4v0h
hyfQTNWXvI2EfIYeiItEG3/2yy5dDSyz6A17q0v9bgSJik4XBA/wXhswyMsN2fua
BVbyYjQzOrnrf79I4unurXk4D39tUIaw9Xak12VicUavERu1YaMieuJm6UGZtfcq
KS/PUFwfZbGxBcLQMYtRY9xaGkszujXyzGZtNUQ4alzmfgB+ToGANDX1Ciz3YBNC
55wbaITu4TAiRrLDds4jlo3WNrROjmEWGxCWrLLafjzmKZ50Y///slOfVUhxab6b
LoAkGCQdgqXVGWah2RTxVHIbkE8GvMUn5QYBASWNJLjH6pVpHcLksUZoi09yLmuy
aUCAoVwi8J6ZYpQEss7KpvjjCWYnC0WftaT33Baz5FJ6+PfRHCwFFtYm282PQKIH
3AbupfNPO1njfGF261UVEeY1OxSwa8b1l/qPnURqBSjbaNqKowI1y7/8CAcFHvQN
AbQG3XwvsPGJkD6spStQIy9FCQS8WeHI3yPhPfUh8DnqyxQO6IGMRltq1Lz5si+C
Czod5YcJoyVWrAyy39qRzWjsanZKBo8rowUC2ZYZYjQvQxbSNjljbLAI6jxNvwGH
0FKgehRxmffXtC7sP5X2g/WHZI+aONx4eNhJwDPDNXweSwLAgqfbyQJpXg5bVBhp
60fl6O/Ngp7zx9HNuwDiolO9rAbYDySvAAC8+YC8z5JR5c8w0fX+APwRgYrJnLaP
dIa6N4eUaMSG7SKIzNRtvDGsdQ+breeSFupZpFwnEVMZ/g3DXGQrGCQIDSVWs6fD
RKjGtV8RSfDpkBcnpMb+pKBN4Nh+sb3QG3NYFSDBSPyIMiimWhQRLbk/OBfCFd5t
pqDVcYva3r8erzcRc6FAyGYsfZtbS8eYu5GnOJ/irwMFlqrfwmV7/UxMcCn6jpyg
ayAoQnlNWB9osUHQq24YKpVYEuFb/OqeBXyoJbVjEnwI77d+t/SZPm+PNHUHau8o
2M5OjczhuCoCge6uuGEuKh6ZsFUrngVUS7uLoKLRVOfESunYz8txnOL6qSiKL/Gn
/tmV19OBynQfyu6KdnqSLMslAeuWdp5TJt0+T4cV9fRkeI/LlcMgiHBnKrlkCj0n
hhg7kweuPXoCnhnGqkv5kJ6jlg5mTvWZgVNk5IfSLRzyUjzEhO4pQR1mDKSPjziw
RL0+3HR4XsKGaKK9D8v+U2KfVftYbqRiZfPsUhmz88YxOWh8CtfFa711X/uEjHjz
CBpn9fmhsniElrZVYzg0OAkw92o2KqQwZTHVM4kycfNnx9vWmH+VBO/UkH1xjooT
zmt4bYs27T3QCNY56JmjSqg0plQY7i8vYjl2geTA6FNoSag8n0oNmSrMSouwMfqa
QCnrX+gHkBLPvfOq4OH5bM7SRXK3V+6AJTiFgmRaanpyzP8u/yYK7D7u/ePXNeaA
fDVhX7uKs1bK4CXl2NxEwZoivFmUWxr7FfvqlfwPZAVH2kghOz/4vxsiDb5boSKP
QGs64X2kqu5mnNIoz/JJnpopaGTl+MI0wnAxp+eCpQTPUhDg2b0o9zlsaO0cYPly
GB5Cnb21UHMygrqAOOlNCcA/A2EhxycZ58QG+8RbIFRbxEpGN1333iPzOJKj4v43
Tuz6k9IdtHJx0qP+A7/ghhzBpd7UnjZ5/FebbwapkXDObNsZLa+1ypKq6NJKQv5u
MslQNmhQGfBnrDFGG8T4yEBz4W/UA/2192LYLb/OC6sCS+9ktKeIWJz8j4H4a/Iy
jjPh4r+OokvMyCB6I8dmoRINgHWPKb/+VvvHn64Ur0ookUe5EdDDphRqe8VzRQum
gtvG2uPFfHO4CG/2x27FyqQQCQ/lt5Q4ArtOdvi0vUQ90ewbvFDOX10JM6dMztXX
WaDPkR5PPZn+a4PtScmQWP1+xGRipwxrI25+7VxIfhgtE8TRdk8tw+yMjvvGHywW
3ZnaMUmml2P08BTjXzzqZVSSTr9X7XMfXqrByXzYip83LFOn//zf1l7bORCn0e4B
GLNgA8yduJ8CCRyQDfYQuPY7eFnqvLakdUr4I5bWhTAQ+p0hRWhpj+Pk06BEIvLZ
tf1+9nIxoKzCkRLgBak6TpeQVv467XXIdr5ghz2sKyH4Gdq4mhJ+w5qmnmvfXePH
RG+Q+TfKgyh6IM0YgS0VdzTe2lEh84TajUb/OfCRnvX4Co7I5di14oJdCCU6eyP2
nPQm6iOJWCXkW/uvnZ51O8TAWsyaXYZsJOAaS81p8kWbt0tH/HLSXny/WDVHMO3Q
XyTLq5e2n1iEHPk4v6kqHvsZSvEhsI2vb4wrjPxKgF5oqstwrMN3e3HBCC957/0z
Zrq9xOxiGC+TDObDwCumWFYIbUx5lPjUZjKpE3cA2F8y22J0jzTDVy+unyD95nZF
Q/+MjkboeOvq82gnIzodJAbMlERpQp9xFrXzN5oBlQUv3CV4Vkq5P2kcPZ1zmZvw
NcHbCk0lC4JDzMCEKE0KoUk9Xb4AO4MF6d9jNhnFnk7wpEKHEMHa/f5mjUYVTqxW
xuiG1m1LQaHnP62ndumhwXnzU5bEDqk4reoNasTZC/e1SYbc1ugHQYygz1EG1u5O
JgnHyIdbNNlMk/TvfHSjKJv6XVFHUVFqb7fXS8YaPqrErft9q9b/TZIlg4oArJLP
rTO1KZ5gT66uhTJOAOI+HtnRiySgTQtcvGUhlj8crTTuV2kNTJnpbCFa5rMVFBd4
ERkPvaKSt4yDBCxIetOYJUjBpUb6XWFtAcV31jxGQXLD9W+jt0930v669UEe86x4
6t2uMza1tOuFrUFDa1H8ZrKAtkeya1lSxUHfx4hPoBmjbvZMfpYVKvmtos7dgVKv
pOcPjBaiS4NjZCo9Vvcf8PDYI+Hf6rtipYKOfFEAVShKfGiZrva86958jDFXwFvK
RVh72Xvhs75B27ZPe0AL3CDAvtjM4jaunbBi6fbCkJXlGR7nAIe6koicBxEBzhTC
ZemnYt6FccCAeof0bKxxBCid58oQ+aL9ldkJbtlSQzaN3LoKuuOfF88rye7A3TqF
XagpEABX+iZnvsXR1KvN3hd6XfRL73lnclrr4hAOfbZndPaW3Sz1l8Nb4JZVje6m
3FACPCKBwdqPY5GoAvLGmHLfQRZS07O9eh8e9sGnX6n7cpX54bMUdLVDDe7QOjFY
lLwtl3lo4+KUXEcqDfN5pfQkH84HGY/HMN9NGSRpAOKR3kOr364x2wU5pLnVAbXt
BsfmJ27WfBeHZx0rd4M0CA1MPwMqH1OxWPXkV+9uF9i7JO2oU4tttqaWwP+MTmL/
mza8W7LqihmFPdICOOhOJzrpsA/YUJ40yqHRmK5O2MhwpTDyV3FgER6Lcb6y0FNf
hMYgwwdSJj68oz1QmpUsKaQGobBhL6ZjCjoqZQyZ6aLhF6Yz8zcssMnApowbfJpG
OskxVtC7m8Z9vmS342N02oVN1dWfm/EBBIwo1WKIZbp6fgBg9+5DYZ+wyrtj2Jw9
JFKAtJdZgKyxzj0MZc+BNxq52FQCmUOxCrDKURiE/MnZ7FKJIQwCN4Hb88kWOD6L
UdyIgiCd5SuYWrp1M0VtreBrhi6cIgvKXziyj4yBOsU15Cvx++UV5UZZ9gn9y7Ai
ON3rDJnC0J4H6O5QNh0+ihkydYqjUFG26cbbKNISL43hQ60gu/QvmGAmw76t+k0X
LDLrbmgqCU0EBWLnGh1SiO94BpCMRKDSmqdqPbc1wM1b5R5l8RCxCHt2VLRNjC51
2vyM5ELPf2p7vUUPdVzVSPDjQ/wuJZYs6w2fgp4Lw0LyVxew2JU2/+4sWYqLdpIg
kcQW+rnEGaeksOz0wC4plpvHBWfGb8fY8aTZJlXyMNL78nPsE06tMuN8Rj7Q0fgs
gdDbycTH3J2Yk40by5xJ+j7QLsCadfxE+0M5KDknwnm30WJxaDxItdlzV+F01u8C
U/z0mfL4MwjPMDLAVpPXdJGKCfanbNSwIDE97hqlaMC4tzsoJaaG3akmgJm2NgSI
LmI/GvKQ7zj8pCVffCpODvpApflqtXWo5ne3WMICB7cBu9fK9JvicOMVD0hcsqW8
WgXeu+4nL6pOjArMFjBU6rv07TXMDJd33S0Bc2U5OgBbDAqojVRvABnnu/cLfD+k
kNS0IuGn6dmzbSGNQftrUnU0D8FiLAfjFsF4w2VGYWlNck3CWVehtC4p/dCeMadJ
sB8vaLfIL0bE7IwfQCzo+2JfnFH+1vk2oq78BVTPSykisASrhtcjcGvHXG4xUl5w
BJJW0XonHJVyQRNBzjAFrrS4K9Q3Uu0TTxGzyaYwOAkBWO03YDVzod14xJ6bEhvy
olh4+KcZI8njl7IHOu/e0xjfD/t757iGZXDYIwCZZzTg3JDIEpoDyOc1m4whubda
kfpktGBkcLfaN0gVQ06+jBqOqv37h4n7JtKL6ns7O2ctoIgU6ZppU+fq5hrQCDyU
mlpUvzNLvR0bZUjwdCu/s7LAmThQIDySHcdSSL9sMY/UM43Nymu+NLbXtgJ+RyYA
ZjF1qOaqoa7MV1OABHNujjkQKz2Tv3rM8hAZR+IDa9+DRJzQVrvYKuzq7NH+zWWZ
GSDEqbVgHEXUaxawTBLeVhdFoW8XH0Q1uO91nVAk75mBsdH0Xs10xsz5801q8OE8
+b2te3AhOyI/sMVTe1qT2yVe3KuDXWRKkFO0kol4fEIunzRW7hvJEDiWbVF+A6zJ
qt3ub2QqS/7JCqTHtOGddTcUuKvAK08IqbXyT1ImqNjO8PoWigXFy2m5qk3nJcmz
bVG39KDuJL6JpobuwVbcoWIFM3jHhHOS2XtThgwaKEYxSNwHm7IgjUsfzHVHSwQz
963vj0JT7aTcqEOfSRc9cqAiX+Zpv+SGoyOMZAgbeu13ExpFOAPT8azTPe/th8hQ
RcoXBsQ1co+NE5WVIZO25fwG6cc8/WXBHp6YMieASZUlXt29m+PCZ1VD8+ZRUlz8
kJUnxk/8rkD80db0Q+O/oWmRDB2Me9Igvpi0v459ZooBVR7iuooquAGxziywqf/M
6ag+n3JhPl30hX44wDVOqpHrbOW7uVSc7j06lPKiT7V0igIRV0RZ5jU/VplnSWqM
XV6YXMUPMAfPiPCaWoacTV94iCv3wNpptJaz0JBSEv4=

`pragma protect end_protected
