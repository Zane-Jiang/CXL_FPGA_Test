// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
fCiAQ86X92Rl6r0e9dLFqHGsp4NDQYNkaznS1MC94IItmZiPmKO78s5nL+/nceAY
yEZZTKb3buNMV/6hbpid6MgIQ9Dr+5l+/QTaH5CL+mptz9vAeEkeLvMrr+k4uos9
RQBdeVlsvGbhMBtx0UIT6yDyAGOeuathUXHfmNpMS0yZiK88DFxacg==
//pragma protect end_key_block
//pragma protect digest_block
gDxQxlKk9CUAv+20tAdbqNO0lpk=
//pragma protect end_digest_block
//pragma protect data_block
PT9fMIlT5bB1ZvM4sso3DFsod94pJLnilZH0HFH1eskWNsogqYXLA7NrH42pKgjQ
IZA/6DIskn+4qFQiJCZ+S9tU51fvo8R6Xk4X/+hCjVBmWkS3ucZbd8/IwBDKq//Q
+8ZzR8Y091w7a1YU1kD7fk4/dinXntsC72bHG47ubh6b21YHAUcivrTmkQllCpPZ
G6h0naBW/Dm2FGBmZ+4YSj0BWEXTRiFuuXg6izA0DngfiRHAHSFxus/ehXhGNfpK
/dr2+sIQ+3DwfnNUD0Q23VKjUmRvkYnJtVO4Rr1f79ZUuNHQVw57XI26k3JTSVbA
nPizQuFfrmVQDb5IVAbnsQ4dYQmDwswCacIFcW5EAX7Pe9Bi6n2IxopWRJKZ3fZx
4TGtfEVpK/r6lLHWgz8+eyyK/87R69gF2rwJcTHM+ZnqpIHSlwyM0Yv8d88mQCUT
Wr8BdT21vFA2ZEWD4eNXxSPoPGu7SPJ4ZaZ16ScuM5CfGCaQ78Hu0zEjBeoGTz06
mdOi3QrYXj0NxBZP3bOpzr2nUH36LC1uR8vxmPrXbVHOd9NfqbMJlmyYmlTcrALg
my0ZRJR/gBrjfHz2rjhCn4PCXJzYYqQtUnxyHEzRVWuU35UTG49PqAjHjiBltYbt
vAhLbBwyYbue+g1AnNhJ/ZTL/2DTN1yM8GY3dUeYkQD4qLTUjbPxLKUo3guZbp8T
L222EgSqMnZfufeVYxDpJoKKFef86l294PQJcPAF4k7q5sIuALrrIlHZf2bjVooy
VSjHteLX+qf24+Kmfqy0tJv1/4MWrUyhPPvwT4cLRBd9+6tIB3tp9w9GuJAngPwl
jpL4hH+n/IGDAyXYAURNn+wbZsWKA1esVoG4Bm+zzctzdlAMK2+eNm+5mch2AVX4
dHXQxCPZCaqEvsDnTaZP0YBX5R/A8vS+Ev19DGIy5yXwQdUmMAhTB/2ac4URFQ3M
3FmHbAvel0YRvC50ECL8UxAr3XqznrQPu+uV8NhVIulApESBglUADRswgVrvHAjm
BiG5AQBeUC1QNW1vlaihV9xBeSz/0iDrDPwX9ENmtVxDJuoUn+ZcXUoVcq3nAsbb
TcB0MqdR8PUiUmWN9Oa1gKsFTj9vqjwfVb8cJ69rjXy985TsuK8/sBMH5qCVuFvg
HwWZLwL41xyAbQOWy7G0GdmKInvBHye/K+zHozAEvaNuSO2ZuB1OfY5VpALM3cCl
eESAntW5wK1A+8dcuaw4/5dTUrfzMtBVuY+EvK14+3oQyLxWHrVKPoBWuotN7o6w
VG4xWC1rWW1gYc3Fel7YIVexch0ZiFA8NU0DxYLX46AiGEVE7jBGIYxQcfwkKs8l
lRugwp2vpjS2yvRC5I+HDoKOcIG+o3dlYdGwRlkfa2kimwSPOPNhkoEvfvgEhmdi
UkSgubqjDvIGAX+OcDYnGc931Vz9oq4hML46G8OEjx/LzlcnPmgdtEpYWYB/BBuS
Lb0cMnbolVfalbxoA6OwmGBoxPO2Fd6cz+WsmX0ExTZ+lQeXpVujMVG4Ghf3aaMI
t5HP3820bdWiUnybpPYIWpy7HvGCNzsvfc3bZi5yERxjSc1WI6ORbw2svuKhbXT9
irGtN36JXnottlndqTVXEc2DfswCWyzyExu6V8lqfnDNdAfkXv7mRIQeUQBx/lDr
7dR0I3XQrOYBUr+RucuhSEAUmz5WRO1+ZKpa2+rntziRrwiywqaAAH1zTFvGUPfl
dyHArDUd64R4u14+JFXfbUQjcT+1JaO7FPmIaS4oXVEvbEOwhevlMtCgeLusBKWQ
U5j2SL4Z8sm3yL+/TquG/439J5YommwDH59NrFBuWDdaj8hw3yPijp5tYmnai8Z9
o0YUypSHdWVAfYjPSYVf5x9c3oSKozczZ31TcA/ruZXmZvw3C8mdJginJZpgqrbz
5fQhEDPcRjAopn9s+CgYWY8RdGdPXdUZcecDAQuTzMbcTSJ0prTfh5PCwvAVyjBY
beYG1PiQ6543ZWngj6AV7yZFuDqllAinhS9YXLuzDVgIjR8cYwYB/wBxdlM2KcVz
6bXxpQxmSkiKTDmw8PdekrhLnoakGT1l+6yyh5eoH3GKQ2cuMvySzU09LIY48LoQ
GOPxn266/tlWPtVMM9RAcWUHhYemLZmxADuXchwrrqvRtiZwkI772HqkPFcvBS9x
lqi3aiekY/gLTThN2HBZ00G7k5EmT3sWLWCb3dQ7uvIOaOjpjmMASI0dEAnWlyQ2
49zuNi07e77ZS6JbwaVh5ZjGawmb+CvDxPaOxgDSd1b5Bb5zFtxmUafe4p2dFTWh
79dHKJMgQsx01fTVrqyN8SdJm7zwaX8YBBBV7628BJ9D4FCwjf+Qw1ShWx2J4Ihm
ZCyo5q7gJATgeNrzvOJ6jshjOkvnnec77gIAo2oX9OtzxLYcAVsXI2MLGPbp6JDL
oUDZwkh9tymR2o852TcPbVrKPQ2q6luyoGnttjYjoNB7BrMhgSJaxcGAHQrh/RMj
1Y34K48/7wNZAGwWaPLBqxef1as2sKaK8l8AO7LNa/AlBjMi7Asqdpq6czGOgBu8
6Z2/5/5bVN5MMMK/6X3I0qk6hlXZ7I2tGIOxARcmemnTTvFypTPtJpzumcjob6es
3T3kUD7kExfGjPd6C+zJNSQvKeBoDzCqPKYCTto4e39gdgG7OJMLVv307Sa6AyRf
Eg0JzrM+JF30SFU2+UTqcSHlSvHudK3gvdTYQGABZS1LFg6Xp1uoePpG9F9NPJ8G
R+RLczl4vGgH7b59e/VgteNsComOQ/C+Gq8oTSv2Iroz/GIjmDUqYF/3k15aI85t
lsqOysJHFE3kYPmp8Zrw0qy3LoQLgT42ch+kQS0e4xWN/MsYekaQxf6UIf2durL7
YYgSJxayGwzi+5thXlRRAKq+b09yGscQ2pIFMrMiinL7FVRA/EbVZxzECc9j8m4x
APtBvuL9MischJckSl1J75TGsC7DAi7nQtB5jAK7Td8MYaPEFmlMdcJLA3sE2G9r
flgykzq5Bk1wHWdgPZbja1h7gngrfstEAME1Sqxocgr4D1Vacj9fRMNJNW1baDhi
ZFStBOBa053sVI67/Z71/eYbl6tTIomeN1Io/2nt+DOuYFsUklgAIdMj2PcVwHFE
EfvgyBUYccaPeVqvBjaqaOJTLkKMBODkvqSk78UsXK5pwU7sq2rZe80g08fd3ikM
GDK6w8pBqyZGxGBuHwsM3pF37l5g2cZn+sxhrQJUEYxb0Y5ABBiKRbf5P/hu3wBU
amJIOEDXJqiQji+DN5+lzvRH5+Vu+VnfpGLT6VpyfHdLtGfS7otnB6UuJglgztCY
ET5r8L+iX72Ay1M17wmEaQV3dW1RhpAOBYAwSP3i4xhzbOiSz0GVhuMq05eBPU21
YsUfmaszOPN8Yl2/ntvSoEdEwAo1yG0WqqCjLH9KqXuHgY8ZRBRiEpVr/E2OvF8g
LMW33OXDdGiQEgezvCi3TcpeXYTx7bvSZVP0t4dD3u0a2FiwqtptjkKRy8ef3I5V
1BBN4lrwKJfV1N3yIebN0TRBG/bzf9t87zjuq+HACjLJAACK6gd2M1TvI3zUxphs
q1QdHs1+z0LrP9mJ8rh5ipsVG2fzP1pDkkeK+AI9na5qPUgRkhL6R4ZHR45XuRwF
lKgFGjZ3GaQODazsnWwkL6aQewM3Nk9pmwOqNK2dYhQhbHfYcj37h9NPY2TT8fec
2OG+kepqHudW9KUeNZ6re0A7uXscJifKVp3CbgfCR4gW4GrLDJeda6Qbj+N/mdQg
c06OhP1AKe38ydJ3PXKS56Zrc0cIMffTZvMNAJmVnIFq12Krz4H+36wvUSSL8JAo
GrrPoF5S+/oVErr0NqxbWlZRVxNfaf84GtcQEUw2YG1aetIOdaqVXc19bku8J8zi
BhaenUF9PEjpXUrfT8hW3sz9forEdczEtq4UwotjEOqkoqa9FBjAVsupaTI7LmlW
Ar2fq1Wg6pSFbFoDVTCcRFloXifQ+VqNUq5OiSsrX9tgocJ9PEc0OdbyZo/oLnTJ
LE5Bq50UOlCOLDnuZNS+tfpBjCEfxT/lzJc4h7Sy4OVc2hlWPEskpgX5LrX5rp7s
BECu0utTEAzI04HZRnexbgq9G2oTxUu5kEFNO+SFOg5T0DEMoja6W1bhQqcyu1EW
oLdYG3b55/qM+vw3e/rMKsB26Ld5KeYKVvLSsfB3F478WM+2cWpKL6m3xIzvF6uC
B8bNsDnYMjjwEWN8X1SgUsDSn+HXi0e+WGchEBfrS3B2W4OdpkFPN7gCGSuOY/Xl
ri5X7Zz93x6Rmg8vMOkIMKueK7YVzMizq4IsR8s8x8t36Tg2hEc0qH19B6UXPL8Q
0MfB15fS4S4wmbRAFLU4zUMbl/88UGTVZItfqTeKPmRadumc9WGYcXocbVPcthLd
5pcf/fKxQxUXRkwVRK5zxoPdljFVN8Rc/5xFxx6dinq33JfzcOe/Y07eJ5znGESF
+ex8cDgGi7kBSp+rOCJY5nvxK+MqsW/0ax7zSTccF/ra1PVBXpCxSQmykJGFdB/o
t2QvcrXw7qHnV49YDMQe7W/MwnjqqUd8FiDEekyGuxvVC9Ia9JAIHf72DLSrlqGA
DqVapg84zlafYWEDL+ZcZ01EaiuZJcQEItWqsyCtO23V0DGaAN09AX6iwYDw24lb
GjObFh5LACU8QKKxMyTdiI6fTtlOkEF2O1mnJF7LB2dajewL0bHLNESB3I1iuADg
+C/eRHEozk68Gu5mqIREH0pGeo+gJz5nblnA4Nf9E3eTrJYCWk0l8Cqup0VZJyCY
TB2KRrZWe1rfMjLkqNk7mwEbd/Ml/ZibcaoNKbGJSTrHYddRjl81XHBvXxcgFAGr
Eq811rYPO0XuwJTwZ5LMo+v7oOvqEQhkVqQDvmWD2CMBoyiffDrLJqddrI+6AbzO
Oz6y1T0LTpvBmN1EQW4sNlK57aIYKGgKtjH9Uakgyt3HAPReCF446JgI0ujAzha/
oL5yMdnMogS4ZFy07vsxAQS7hTxL/wOhXeBSmbbtR5xfiRFQLAUiwfByu5syOqtq
BUXZ2K9LEreuGAKsiScWwzESAe+ZN9GbV05crwzzI5smVo8BDmHuB3SwjNkW+20Q
haiXbm73/Sz6jfC2dxt4xMbEx5qIRcH3uUL4qJ7EBxENNjvAVdqHjcYpZS6UCNDX
14r6s1HjL0OViJlA4FSxRzupltiKtmNeAxqjZ0tbcjSlhAe+2vPS5v+KdkkaWP+0
eSTZ//wwqzcqbypH7ysr4ym0qafz3OIEQsg0oPLjoFAgx6uW2tawOeR9rkk4q5Ix
z/+7HjPag/zXQ8FKBXgIYFJEgwc1byw4tXrGKSKAzDJpOMKjnnWGvnI2X/pA1VFb
+kK+iCd87WFiPkj79aleLWmq8Xkyp9XuCQ9IPPxy6+7qlRv3jlc2V3w6E06VPRNY
bKNAkqeE+6yZHaFuZ2UbFoFK9lvOll+M+hF0BXEd1xTVzrMgZrcn6mbxjURvn/Fe
LcQMpbgxKV5P0T6JQvji7+DE94Yj5NVbEJmOTOTc/zVpULyhphLv2j1uaHn78dZq
7m3s3iNyc2ZzYVPUc8HzxTcd5emmRzhK73ajj58yKTq7Dk6pQ316lATL5snuiQn8
C0K4C+IFQbwEZLb9IMHwDj9+BxZDvTFDGsUyItiVgsqvp/W4qSNpgzmpg05YkO9g
PyzdMYa6xacnrwpYymtBBx3Agb2BCOZY9ficU10oMOlbl+VSoI/uRyv9DcjeYNHu
eMpNnclksXXYLXfls3rBD35F1z3V9V/+jFvlgCFrOTZoWSY20VspJl6W3UGVX6YH
4TiY4Mv9acyo9OiQVk9U1AJfWNC0pjnVo1vUBEy+QAoQYQpztvtzK4vfESmgU5EW
J8sbcp0KdGs7qQbVHMt6j8D51Mx8qNMuoOIYqEmUpwfU1bd5Ysd2Fm+3NX5n7Pj6
luoyc8cZQypEHfoP2kBsRrkqbu7/lPJwimiSS/1Lr6c8+/F+rQlWcd7P1yNJ+zf6
b2vSx87k/ha1Mgf8iz7HSnHqxkZ5SFGCidqvZkpj7OZeXawviGrbKfrKvNk3Orvz
Em8BhFqEM1fJfzP9dP/AiSNa2s15iIXImMNRmWTwKkNN6V1sHk1Utiwi+69hDp7m
+ZL0eIXqWYzl+ZedfIYeTC+Pq3METg9VfPCxc1xhKO01o9N+XI8Fr5NL7TA57oSt
aUd3M4sCx8sGgEZ34Lx6fIaN8t2SUNGEbG6Tu0zRaWMCwryB5N0mckQl3rkc2rwC
9bIHvt1B6basXaQ7bUBEt1SpphPd0d4ZtccFK9p/OtqTW82giLkm66zmodz6VRxf
Ol+PFBgF6V9WUGdU8KN1PKzPYnyFbDPsBGXde0nh+LXY8IVu3Sc2tluISX4MBTpe
ZyQLin5/gz2biOXJ0MvrHjyHY/IlI6B7TCrS0XZ+BGJUwaSOBnyYhi7Yyrt6zICS
oeT+kT5Egs2WH1Spuu3IkRu4YtXFiwZlJTAXuaZdJ+p/k3DqSLIp6HBK4ifcnKrG
CUM8G2BwYkE3CIZK4V0q6aIi1+GnU6cCrQQvGREuoDZ7dxi5+Ca2yWGxQDbeTcvi
jC/uzkGHVZdFNMD2DJ9eF5NKt4PBvRIj/KBfYD2jvfD9WBKYBlOaoZH1jvwZqvMC
6F+Fx7PE8Qw+HURQo5pGi2cSZD9ytJZ2t54reJcQgSX13KujCOAgKYSiHAClKOeX
jQrGDzqRO6ioFcHflEI4adZD7RfCeQ67Dff0KDXsoegXDYOqkerg94bB8nisdwNR
N/7wfam6tKW4FX4ZRlAI/ovO7nWu1bWuyIIx7LG/hivCKMiu5pKimnOaKo+Hz2lG
LmpIEetcwggyu3oGfCRTa/wjF8cWktOdKDh8Sg5YjvhFv8xjUC024ZJboAGnGQr2
ZfTqO4KVbVNPqezTLjWRO9H7YTDe5RatNI698QYay9B6v4vKGlvacC/p25XCfjYS
iHsH8gMj4cK9qeKmDaeBA6KL8mTY7mkoBy79LmA1db2MbbPtFRIRY/rDm/jYDLkd
xgUbSR+0tdUvAB23C9SLd1ubib0RVHKdYVdH/smOJVmTjI3nGWsk9UAhv56waJd4
IeEoZeEW4TXzC+zpIltK8HxJEF6/2fnkJzPMmtwcDG6Db4xd6QhMXxZFuU/y5DOh
dvqao9uthYySKbonS8XvLpZNC3SjjArY7ZVPv3EBP8IYO/2oE3LVvO2UtrleV163
A22mGj6DjJ1anr1pYcqQhUEzZOBx5I1xItr3hxaexAuTzdgV//eGWnOTxty7ZQVX
ARp6nHEV4tu5k2YQbf76IdLsWTXBWCxC1dIGnA4OJBh6hHBagO5RwUuS4ueYgsjw
id323IEFzFephBXOlMtQODlm9H3c9t43EUHbhCJyk3UMkd9OClINndtvhYZdp3XB
DYzl8eqs0FjnKogJMPZjM920GILKMohbLpE0aMIZp/H21pDG70t3sKBJTdEgvCqZ
+xP+BWcNSS8JqtIgszOmwb7xsrJ6igdw+uWuz5Z/SCK+9Z7EuZWvjwfHZV6f5wTm
0RcAlrayraE5fIagQNK2dJ+5lzi3cTex2RD3hc4FNgej3CFH75IZJeOF1rsgwDpl
XFDWbB3FMYLTiY3fjMWZVxxQsxsybbfL0ri8eUeZfQJwqLS2M5UdO8vm/772GGyT
CHPYLjIxUy3UpJj5e6WyrN+jt1DhResAK7g231XML4s/pjgOJeOldi9yKiKcCZbj
Ppd8Wvn4frRiZ+0Q7Hbo71eERqcoyOoMZTPlbS1SSevzuBzjeCyEy8LGar4q2L2H
FS5pjCbMJWThBBSbSpZTTy0efwDbcFrgRGml5zNPpZvXy47jSs8hjj4exRBsEYkt
wvFoZaOMDG7g1ch/u+k4aN5Av72tDUEL6Oye6XoxqhTRHD/ffNl8tCAgQMVemjmL
73GS7dmCvuhj0n4UJxBSEwXbAVDieQBpLpenDALUnIesunzYm3bjfB7TG0yYFY6y
cLwolgANqs3AmbDz4Hq+IpGETR73E8f82YqMYT27g5f56xWDB2rDlOEAMajAkfpe
tMXj6q6PQiI3RTkmytFWZaMzf0/3MCDIXrSKY37Fvr0mntVG5To+hxUZzNqR5wXz
IfyPVjqjWttILheA2vOuatJfMjpQHX7Fr4jZ4TQpen2SLv1O0k0RQLjhNjSn24Py
+er3Dc5MUJHYvuKV4d5WWV5z8AWNAGlsTddQ5pVSRxvBpLoJWcpGjxBielW0cijJ
XsEFh+9ubC28SdpnXPXRMZJ/F2knjMQ3XwbLaIv/WH9MrtbM5goeOOBc4WI8dAxa
Zh9NY6TSlD8jtQlMoSVfVmgqQPJa/uMcw6XcmkvDNo+FWSVHkDZg+4o8zXrV1zrg
lYHV8719LxxRIbNA5KWcW7vQJGIbUFPIWpnVmdq4xD90fuLJIRt9YiqD/Zvked0g
Dl+Gz/i/1BiEjyLzaGjucuchLNvXiy6aWKhvOHTK+20BKTzbgTCm+Xv9RDWRfO/5
gKpWbY6o2dd+eOsQTlQnsOtJSTMLEVuiO+2Wxv6HUclfRHqSzys+/o2Kjutjmn/j
OP3GnP9xQhKOQnXOidFvUDpROZC5z7/wviRVtwfeRhgQlDijqZVC63vSYWiLtlnU
RasdCca3baKc13GsPR7hez4m5photGKhtJeO3VnysGRcxJxpSJfmBlvguFhulwl8
JNQsGA1veNyu8DWXt/m4jzj+sM9+5+ldb8pu/WWqctrwg74VVXC6hNydeeu3VgtJ
k2o8I1ATPg7+5+yx5/jlzUKGk+LvhYyHMQVrPrBJF5O7rd2aMkd4C1sxd1TTIQkN
xO4Xsm+hnpLhwB4ByGSQYwt8RfY2Xkolp76oIsHg0HyHEEHEYK6S9FQOuFx16LLS
atJ5eXQwyG6un/1lX5ptfwQ1SxHh0QlQsEyNj8fctNhdDqyXbYVz2F+jHm+xrgZN
ErPQrmkCfdbsCKCl0EaNHL7MCOoyv6KuL2Q3o9AvsK9lAVkxUy4+vPloFjDfFo08
k1Qr0hECF5xJLZaRPerHcECcntBRH/v/U1LCD0SPbESxs3Q2mXWYjm/vq6arNtMs
En9DHbHTVl6rmYjC8vsgVuscrbDSkMzDoHefnr5QMMG/LSsHmf6JJV6kN3ilbKXh
61So/XWS2QykO9XGQjxbbpSmAb8+c9F4S4TxDBXobcUOLwvRz4hURGpaZrBGIJPn
pLTl0DBqWb8hQY12S94S8UBDOe8EzTJYzHD1tTq+MSCBdiikOmVYXWCBWPiMtN6O
x+1T4YmTC8ljGCMJFOtusHIXKl0wTQdPew+h4TOaPpqkekDGqoqOUFIWduV4N8S9
OBLXmPDwcyp/rJs33gkrHDGIckAtmHDZv8r461Rklpqoy0cPFYPN+Ex4G8feQjhB
YOGo2TP4gKqwrEY2SVVcC0nkLe0VDL5260jXQmtWaoXxlApZiqe+T6HjHFiizrBC
byFdBwPbTl8//qoiTqt3rlgDA7e/LQtNZl7JxrmtO44bxkD1JpKmwnjil3l6BKD/
Lg5A7zNoMAlMQPAqilhhaCfbii1aB3XJU+S37ecTbO4tmLWS7lQC/6S0i9Xl3eGJ
4ntAfYdEWll2QIPsEv+NUW0IhPgu9k6LCJHBSczqPVogGdqUVbQB6V5QhR4B4csl
Bf3ny2cuYItGbWaFSdSbJ6gJfzW0y3mKWtl9X/oNWwSi/DtJgZsMoI1SxKhGmqaf
2fK6d66ssn3z8RsB0CAe9IIWa2z/eosBBIiE/8m82h2p8iZnHGhlsA/nvLiab13R
6QYWz0cp0V4h20m03HvPGm8p6frQaNVHISwWbygcYyGyVM80XnFqsP2D7MjSpvbr
mXgRdmIZ9ZrSdHxfY6Xjl5PQXhwTzQ1gcj/JRNemi82N+bATlV3HfJemhpZLe8/S
T5yNQ7vNM7JMN5v8dZFm5cRHVeKPfL5HP3BD5oobFT6uKX4yUE1thjPK4ZCkJNeJ
bH6G0Xtmvuk7L0lRI2ogIOLflgxD+kggPR51q8Y/naf9TSY1/7CmSDCuiygrgqWO
glTo/XMdNzJfWc2M+b2VRGyhiKAsU0zb5F1J/8o4jTvTtN0+o+3cJAtCkU29OZEu
bn36KFlpZbAKvcta/KT3FSS8Z3J/aJL/7DqIyXIypFVhRL0VUJu27xbLNNpHM16L
5JrBT65x0sF6U6qDvbwlVAOW7lCc0Nt0bYdRStQzjRsIdhUJn87DI1AYlVWPQUvN
Y+pYV3vdG63gQAOhXchUsEbR/T+xKuFQpzipXWWI3ceFpLg40JHgL1kspjzDG5M9
2awOesaCtHL0v8OyYnXOumkxh1diHTTQDXGgrUadH2tPUlekpbxq/0JNYa3G7Raq
5B5sHLPo2otjEKK28ypBQo3OCLJkUmwKUupOC3jmZpG407jzKJJsVgK6FxtFjZuG
oswyMyyCS7L8dFtDa9YfW3R5a3lL/4G4SSMkusDCea8Xy5GeIKYksKOHnoGE48+v
3kU8yOwRLkaDLHjdlpSiUTMti8hGHnV6KGCx6D/8aPwigEO4V7eZFZuw6h4F6XCQ
4BTAy05bRaWr2aaHEh3j+BarYPzY8IO/nraNyO1xmTEWRvKWWiNNrwkkRlovjREI
HB+2bIqLcOSgfHiyCN3/o4RHcYTMPSHzpWPqLYxHsfMKxwE2wwXROinpcZ55pgfv
Lq1KL+pS+9AYiJXCIlFcikCVDD3bxBwwJC5q674CkQgD8leBYBRSmd5++I7jO7Oj
CfHO5aV7m6gqaTG9pA1dclFHNwYcb6U5R1bUZZDeSR17r5CnEdtGvd3GdGJQ9VkT
t0GuzQuABq/I1D6lE/A/TIl+uQsl1CkG05kPDFyKBY77iQVVGqmqAbVaGVQ0CkFg
6UvvxKLOFQo6SiFnPT/srVXvTIqTqfp3SeJ1/YRvyfN91d9SR/35e3kliR77O7x2
No5wYSv89G9LDs6mTu5Wc30b5sFVKEtWGa6dIjcbb50qJy75byX5Z/R/B5GB2/gn
iKmeJoNfKSNYopIUj5lDzmsz4Xn6AnHEJ3u1LMZ5ffn8B6qe7/bNp7NF8b7XBNd2
wnS6DnazbyRPjygnthjFDvKAdIm8BXlPe8SgLN7piGh+XdCobvgf30r1pQ9uOwW6
V+NYlCtfRwZSIXuY86RyOieReXbUAUOTo7uTXYBmqzl+5YVn62NmN9TzKrAbqcQo
kQQVVsNqPTQt1zSIAatAjNyoXFH/PDVt8+1n3fAlZ6duAxkP66sRycBoOdEeZzhL
i6MFwN1TzCaJfXUOjyyLXDYVvVNeIV3cegz4dg9+9lVKSrAYLMk1IF82fhjBi8Jv
bvYuXpgketwQv2HOeMffD/cwrN+dHt+2XftEIzq7DP/Sx7N+BFzeIAVRMdOJPKzR
Zyh23fomkCSQ8d93t31Rmol9UJbIZRj/v1NkZwAR5t6sRIHtkTNLJY1mFQ8M8pLT
cbNGQb9kP4Pa3SN2tWQMDlzGkKpsG2dfTivboVRvoMw3uk4K098C2LDA4NXemEjC
07sJNh5GSTuNE6MaiF1tx5inEXUB4MUpXJEncL06XGYglGlwLay8M1BnahllrCEA
VvOs7ple9unCBIPigDIp69WCfsl1L7y6hWGMfV2N9ZqpFpiFVqWx+CT+CKyzbPHg
zN3AA6GRFRz7goxVYTibM7zttxTR54bek4sLqbilEEcEyUpsK5w9clszCC1j5Z9G
3k47AM47/9/8gRaaan1zHz58nZhcvdUYF0wY8vF+oTCD8+BP7NBpcavmkcxzBKiJ
IMNdqnDOmB6gWu+QDhGGTd/95KdaFQ7qxt8LM1I0sM3APW/dHkp1sDW2P4nm8d1H
znbOylS1Tb5p4ZOIR3fSS5PNZjvnwVBwHZL8ZBtsvESCYL47jmkpAPsxSjWJcWmS
lIRnW/rVgZpmAfSHsT3m0PLMVbZbSHZiaQxdePk9CxrFRt6I8qZLUaC/aDTHgaQb
vvH7M2j4P9LOCdc1H2528K3uJ7RLHRdg5z1EJ2ZWdbvNkrcIA2LQy2j6odM9Ar1U
1P5K9BJo/QChdbpsLQj9hv8NO8XmDvES4PaA6Z4ysfYAlb+0k/GwAIh8kDpO9DMq
o9ywJZu7u1r+kRGtLpDja66vQT63vwX0Wl1nh8EIIO06yBXzjyLLx/iRgbYHVL1A
UeFhbGBC1Jw0yfFVCGBvmHH4iVBK6zrEaCsWM3Gfip1s2mXYWaaAhcHtvvNeSr6J
X1o1H+UJ600mh6xh5vRq1NYZYc/5IDnXrgp0A6yp3nUY/lviXHzrxrdbrQhtOAic
lwEmXGcgpXi+2TX75mm26AyaScTf2vO2q2EF5++GPsdp1d6H3xaQglLOvZGgRffC
4mNYCgP5zhN8vhSiUhtmx2Keu0IXMn4sLvaf3HXPNa7i2erin4zfIVhmC779W83K
rZVrgY4AjVuFzL/u/iN3sWnrnpM6yNp1wdZX9B5sdH6pI+WbPySpEX4yubJjXQRI
ZnlVbHAHboSDl22ATqxkqXaerfMU3dQAv1USrZm/5sEy0vZ8UVzbmEI54K4mqAJC
1FmcWR2FBeaGlXlOFJpu4XN43cbTQU0X5gppJSvGq1UW1rCUMhfLrYkaOqONEvJ9
6wTzoQOxU1lArqaq83dEf+R4GP3cTXxlHyBif4x+Nq2pHH2hgJOeN2nwbuL9tWEi
iO3hyIE3YiCiIVPBcYy5X8YYCZoxVA+CBLMoRriSxC+AqvlrxgUkll+b3//Soagn
yFVuQXyuIxILLa7u40KfYS4LV5uJWUw5j9igZc5VKllsH+tAbtJFf+K/t2UUljbi
nalFSb44C05jAPE92JgTO7nWGySWUoPP2vwfvvPf7uPlgiMaPmv1aolsoHtii9wB
rAG7PWJiVzIOM8wyKLYy0GMt6dqnj8woAFGveMmb4UblBaLCGYUrlG9InLPcT/BY
xHgOiUWE+yYBvbJKXFtPGdb14jwVRmeKTnxgPBxH3MColubl3QbH+ZZETMqr/eAj
A6KIykLcR9eUlxkDb1ll2It62cpB8DhUpbDf2P/qnT/K8xwjigYvwmbkF/PZzpzo
8f0WVGG2NMEE7xowclYBMoYPK3zgHrrO5et5zBPcqx2JnTJtUNdCk7lBaMiT+JYl
TmIqJNHA2Cah0lt/Ui06IAMjz81tBEpRBZNlfIkYhZGC0mP8J9s0Tclp75VnDaSr
c/B9XxfoDAQQ7B3+iScdjy7pVjylW9xpsSEFUVYsNaS9W9u6aJyHPEINPWtvPeVj
gbI3hYXUGzyScFLVoCOwsRDHlU3rTBoqB+6wPfGHrdvzv/hc946B4lT4QiCeWXwY
QrBaOJGkp1/mMEM+YBW8p27+lbZFOJTNz4PK1/d/tXAO1DLkMWVOPj08EfjYRl2M
ayP8itzsTOCEeHu5QP8a4L57GFGUOCVFnRViRLVWysvCg1ssdF5Cyr+eXEGnzhMi
cACyiMHD+jq/Nx0I0agIa69iiNZLNYir2uOsT8MjhxEkStZjOSwZ4bpTQHidK7VN
/00ISOmKif2B9vffkiKIQWN72pWXcMH1D0vT0te+ic1GQHqFV/NKvZ3TRmsAIf4c
JwcU5DbSHQoxC5vSPRW7VTmmp6xIMrn/48SBeEo/pHeVduFpLE/CzaBVwANaWBs7
vXlhy2yhwPgzh7GSPq4lVYrKHvAPzTyjjUbbTLS+W/nu4WGchQXFlsCSJ3uWyK4V
AE0qbHeI9ILb/qSm0xX7Yo2gEFHzJyhkrSzIL9Ztfes1qG3gJ/Xf6HJ0uYHqoywm
2vsvR2FMNzhnN7IQF33mgT/fO+qMEtxpRPZH+e/420JhtFM7Y46MLOaP30w2f9FK
MUI+HKfSTlgjGbfkK0DfVDUPRrt3LrS/EKm+o4saaSqWT0mevIFJABuL+Jmuscf4
KHWynAK04zXo2Dvy0D2lD8H8thLymWvxn2Q0WWYcae4zV970fMj2YhBLSGbq+Wt8
IN3WvbI9Ae/atPFm44mUDh2O5hGs2JycXSG8X292kviKn2XaYDZYaiYYgML4i1xq
6/xKJtWUrqbWpHKf7baniwHNeNlva8x71vNWcjCjJCELsJOeNRboMNv93gCFl21K
pcmcCyQxaju/6wpeHpDEnfI8pu/HU9BRJILHFYE69QpC7tg50kPaLmZqTJ0aidvI
wv7osy3BYhpoidPa37QDqDhtXrSpko19luiS99EK/UUl4KHvg5FNP5Hxjdufi2GX
+0IlOKdzgdMk9igqrIqpuJAeedjsUJoXrwIa4RzvkP95TL/QEKCjxlEtPfpAydmF
MheBh3xeAtvnr5d3M24CLjdz3WjdYBKFSWYhlIA0+0Y99J/OUhiMz8Uhlv9T0Rkn
a6+nzo/qaCEIX3jMg8eNB6xWmSVKz4f2wsgSeRxSy+CsCogxvqa98sIhNmZs1dw3
gskOwOSrj/sbK2EontTjHbw/sRemzlzkzdaNvc958JSEYez2+zP5RcrjddFjZPzM
7t6ezWqV7KEl7LBbAF/GDfJVJSxRPw9gTnHtns7eYFA=
//pragma protect end_data_block
//pragma protect digest_block
DUiFOrVar56bBJKn4UuFDL8yCII=
//pragma protect end_digest_block
//pragma protect end_protected
