// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
dwg0LW8A9rPcLsmtbqMjv6io99BzhmUL4DK+WTjwjO9RVcscTj5t1+rX3je59OP0
1FKz4oE4ZDpiG5JTC1eqGtMoHYVoC7kYSlVIr5bot9guoHClWDPEemjgxGzNmngz
GUh/uxtLxRQLkHLKFk9R6Bq1DRtb2j4P2m1LLfNz8tk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 57664 )
`pragma protect data_block
4z8LFDNU+zarNRMaKBVchWevF1gn9q45P9KlItrttMjWfDIsBLRjst680S2qRdDr
DDLU/B84gFA1sI5SfVFHuywTiCWeEc/+KsT+WhBPYBj9ZXrsr1rzFd+r9407iHOp
oSMx1QCUBzzzi4M+ywvjHfpljWqfjRAk9sx2oeeyzcN+89e/VvEVSq4Lb8JaqMde
YK27ODwBJJHR5V5mKilRD8twxjspIKCawL74w4SO1HeQcSlSNf3eqp2WSWXdtdg3
JU0990p9xGr3nLZ92hPbVW+WpuwiW3TvAgjGDXN+4SWDmqAzmmN2C+Qslgky3sSJ
l98zUqvOdN3GifiCXs94XK8iYfBsHc++1Fxy2f1SStuSyCfYUDBw7HOZcqO0VKN2
yCAFOc2hoxNRqv/6gIbHnhHArVBurzErQSzpNeYCgOgHB+24e4+Q1aChd3jFIBmS
9cWLEzpah7pkyUftths7CNuLE9QUJvtCyvZXqM1AMw2BoKhmwo1itEzXjq9AF3/w
5WZmPgOetxJbftY8g6xdxpqimohYbpHfmKnTAigc0QaBi/UH1Beh0gU0DoiJTKXD
sYuB/Za8ARZBOY4LRlFKRv2hjBmQd6S5KQd/TM+zeB0s/YXhzYScEe27TomiANu7
sko1tkjuxUrtBaJsckcVsb3Vo7K0TWgAvsKAz+uIAw4njDhYmVHpuXl9RJIagLog
f6RysszZpKBIdyJUiJH94gyMjwfAo96dupcQGWUuLipXlSUPgdHxRltq4InKn7vM
UNYD8DNf9bQMShte2MV8tycF17HxX4Nn1t0fVFh5Qae5OPWxFYGKtQeGT0NGEiE6
tkMUntmCXqeqz4UqnHAZy6XolBLo5IPr2bfDtrKmO7y1oUof0bdQ+TC5CoQ4alez
oRA5sSOXOy4lT7fKD4VCqzfL2Xc5K22546TRartKCZhtys7MVpb2P5NBLu66TRYK
Bq9VVoKRvzQgtE77rAzPGXpKaJkR0+CG6fUKqwJoqYJMkUBmdTip5yIjOJHyUd75
98epe4GFY1UyVG5s3cPsumrblFio82dM7iMO7lzKkWiAznVWPNN9tLEcQqwcQF/D
XQ+3zgn58wgMuvlmgZRoXzCHDub8TxZOG+zCWXmva+oEINnKXy+9Kv4TASShPhwu
YJGif3y7mj/G3OQzzQ1gtwh0TTP5Kx3q1+L887damIXw12oK7FWgWjzz4hrTUcGf
PJlgrbH3+mQ5GO7stzSEcO/7v7PcnIM/REQ6tzZVYs7eBBY3n3YWP61nKjt/qJza
GVIzgRyTBTqR/6d0IcVTvEOC4h0n3C3u33MgU2w1mLkG+i+snnVBh52/O0AN/LWW
llpPkK8CtKhtvxo21aYMnCK7AjmMw/gu958gZRdFDtfANqGrgxv5L3HgENZqWfCn
YvTQtqQMjLUN6ishzqVyfMO/FP7+p6AQ+v3vjT1fKzpje7ndxtj9vfUz4nAji/SC
qiJE53YiMod84eJSyqGiQMiJ4K51/WUlEoPZLwgdr+AUrh61eOvQ+bw3KMqPCjwX
sieJ2084hzYN+oop4JUV5DvT5j/k54QGItObx1dZ9Kdq1dIx/ZMFIiSAe51x9qV8
qgM55EbP9Thrhj+/l9zRDnTWGwpScxiGdvNvVudvjL1kIpb78IVriSLqKPSlbqL/
jgalz+XePT8HMm+bVBiZrNhELv7tqZoKsD8bwhXRWOwVWVSJhwAez8KY06/RfxSh
O3CnguQNPi//NU0w4hYPuCff7KK3Wwhu80sqZe7tXGDeu3RENhKJO+kWc4cvbT/r
IdLEaiHE8gChK4IrfvXAIS0XK5YHfMIv6rxX4OwZz6E/vYNDt/k134eMuriGnLvc
+beIy8KVemMNrXa3+6t6lj7aCLp127rN+83ONOLoNDo8v45lqSteHx4IrNm+TcTY
CXjUmiiUUtHzhUE1pwnj3K62cxphMrx33eSajmKUzbJJEDBwSErRw9AkIpz2yHC2
zR0pbEIBfV/G7+WNcj3K9H4F/alWUhT1ObAwQ5z1iU3KCQeDdtgdLfqwXCAIvYjp
XpONC+v9nb4Hh4ffzxTOs5piv8o8pKH/nuv4Twe352LZXjlWl3zr+isDD4jeMY3m
J2Y95C9inun70u8YzaW44BjBC/eihv3OxE6t7tkozTySN6yokP0grZH4Kd5h6yuT
8klM9TNvlj84vvOIqc2xIkvjOPWq3GLHhUPJ130WJLipWoXTHMp0z1IcHOdvq5WK
4ABgvRcTNmYWZhF/PIl9WwcGjeO22YQEfxAFOnyY8g9k4zlD6mD1PKOLMDosGmdv
NKyUx8+4uKbH2oLkIJPqv1hOryHGChiygFVf8MogFW9I+YM6BzayK3fA483JZYx2
DZZtXHAO5xfw+UdqdLBvPd3ZEDXgs4zT3LbMfckHYqwTxJbwSJRnqPn+g+bi36xg
5s4jMQBFiyLTUTR7dGUuozOBErGor26ZZllhhLhG2IB9FUSC6wbGdWLJkOV+ht8K
Kwv7/DwD/hMkZuDty4VnLpXJWWXlzh2ZjUXF8k6Ppz53S1KUoISY/hmUuIViy5eS
/leyK144D22HEiLlKKwwbTzowz4vBDuz1UG+zS3F/tSRnW6ClrrMmWga42kpWLSH
1iYkyofqWbK+QC6xzAppFJA6JSl3+TgLRkNmFhp8zZQIwsPElw8n3IDT7b+g9P+R
Cm6c0Ib/Gzv2M+4bA1Svd8PrkZH96FPGU/Pt9tv5zRjgtDR6bkmojYpFRnlNlw/T
Suuqq9xUuN7rFQ6KETqCgKpFbmqZ8EU8Pk1ZCg3cOUHtImb6Osp88Btt5g78TCp/
rOTekvpx6U0LbXteThM9cPbVcASwureRcCQYuKf05OzMkY+NwSq+nBQCxalRCPEA
+gnetP0kwAjZOgBFbQM+G2jjVcPqSgPOT/s6W2HC/Lc/EF5te/UO974lnkYWR7wG
hnSRDbfkqhNfNUKT4Wbnc7BntSVBQhLd2rIoxSIgS7PK7ASqW3ELIwOjwgQ5q9yj
ZWct9u1T7XbEBrTg/5Hc20OOnG8gOOh2HXpxycjs8GUb3A8OBp5F+jxH1SloXS/M
xYM7Ei+ZHuI/OW6yxqHT6dQIma3/1rRk8aeKSfyi8ttGg2dIiATKGfPThoGZ1IOi
F1It+avhfqNyVaVK+6BvVVUWI5GkJ/QfavkJicdYb4QaRW6kbxTxAEZWi2IExH/N
dIgsVmq30VTEku0QwDV6aOmS8egicq65oTGdTi5AXWyqXQ7Lb001OMHTbh2X4cR2
EHyUWXwiZUwy24fBxq6mc/0hVvCkguYJZ79ojaLgaRXm3hPP/GeCP+CD+WInnqgS
4rA/JOg9RfiQQeb/tcmROIlvHWP1PIvsqLsBaPWnWJgT7GniOfhj/eKigZdwx4W7
kd5Fu57ew4uml6PDXNJcQZB9QyR8pQ3wF5VKbZ3iusHxi+nv2rN86R+LFyQ6W6+I
S4+fMTe510KbkwS4BxKWuPhoGjDANl7ak2yMd73xnk6sQ5XxBcbXzDNmIRBvkvNR
mZxkJ9P+s8fIiA8fGyxh3lAbF0B523yBCHhgVRV7dudJR6Uu16nz/lr5miavr97v
2v9/kaTVeYXpeOPReERmDUPk49bEl/T2dQHNHzDRCzZ92nYfXcXI57jVaw4JycgB
pypkzs0WytbOkRHXIreCpSY5J3/Z8FmH9tQ0i/WllaOx+UlwQlEpUu1Glmx+7Tar
vXWHU42AmOnfIXlk/Y0OCRIhaGDLuJlSQirk2uQh6wiku//aEBbLciHxf1i0zZqm
1jjhL0GLIa90xBYjqXVR2UwEi4R8XOmAhFhJ4QeHyTF3MiNb19xOgiH0uSjem+L4
O05IDWgbppxVqdmOtIG2Yb5eVgCm3KfWu4mDoYcN04HU867ggCPpO7FA0v42FLf5
TxFIQCqvi1O8UXclRiPAMI8YYSmJL+SIhHHAInSgPqGc7BLNrxWvFsWH+UnTrW+X
MkQEaY+KreytjjPQrq39M8t9xGHpTqLxU1LS5HRTuKEftFq2J1sSQqt8K1nyOpTz
Sj0I+I0VTaQzYcO7xB2jiGLGRAI+kbFkfeeXJmRKHQjhColUTYeO32PkayjJPl/3
XhDJeGvv6ncyt98RgswUmdJgCKgZs0mlZIGDs3375J5CKsNVvcbqAIJYP3NRMa2O
BgjVEzOeFOCypmWQ6Wz8bL/r8AW0zDNM4EzM5QSuwVgHyzEqJhM+AM55cc327gBd
j8nMmi8IvAwD3APyEKsKCuyTtIOS0h+nYjkYVVPrKaAFAE8ldYDbKnjkF6mm0FVK
ENZN+2ZN9YDIhzINnCg6ash1fB/OTWMj+m2h6Dcu3+NsrpYRRu+aPTF61ioErQUD
gNILC4mXkmPdywV45kJ8RgB3p0KEV3PsfTkIh37L+AIRMGNTb6T0wUMfgqeFufo+
H4hCy5wyyHrabNVHflO0h6ZCXlp9Iq6sf2XeNVNq8PcdzYBhXN/yOw3JlRvVBJyL
3vm/0Q936Fij5Gw5wGzph80J/d6Sp3OXBuBOA83mnBoQ5WHf/ylxwjXARtzapOuP
xRF6+HTeOrJ9CZc9XztvwSEmc7ytzh19yyG9y486EF2MljUIojkiEM47zwZyjBoC
PM1TjanzLhtUYYMP5mJvtCXsS+qI0GHR6BpSJ7PQVTCJctAHVRweJ81icD8DaU6+
r9svez6L+hyfsAgMWElW5BSpqMQD4/mEYlAo23SYC6+ArlInMxibCImAVX46EiD6
o8IalxY5FYrMdmhbNyih6pnQnBYYAQdqNvbSwxbZrSlMA2D2mrarX4fXCWQt9428
JFHtNPVad1uuQ25Q+9KuBdFeCWY0pkY+0RViXv7fCgpph1hD5MnZDQ1loNQz2QFV
tws7IyFbtogUGYAGGripbyjR4qOQ47lJZWYhFM5+Z/wuOT+8byE7yJR6fD7yx+t6
BxtzdTINPp/mc3O3A0IoayFgSvnZ6vrODAGBje4ZCqBqUaQYSo/7yDFzJ7LYHCaE
EP/lA4sX35qwq+NH4edTp3HTSovsUv5OCRknnAHdDcAnCWYsykYxqBFIsw4bpwYS
vQXL7HX/2acXXQk0dPd0lZ2I+gyTgmYuS6KmTyGfeAD3hZV5MUTt2N4EWO6khw7e
izIY36u5Pz3WahBgri93A5AJ7MJmkZ3aJMEHpCS+RIVln/AqYq5KNQEsd1xT2Njx
rhnhXZ+EOaESboyJgH33zsLQifEqCBmtm4DHzVW86yHGX0IE59k1YZi7kz+/FKew
qs5/tTmzzUyebhi8r6sN+rIXiNeUMEyUHDHOfJFvqK6jhdA264HacFYUqg7dFQUb
OXyUG9q09DQ4LVuQs5oj/Or44CLJ2ZKN/AATjpcoVKVyUa9C1Mewc2FbXoncm+bi
m07xjVQ1efNFpaeu89Yj0QOToIVvB4ctDlHEpqX82v1XTCJwmsnkoxciKVXVBX8T
8vTZUdUjO4saf/gjyHGQLS/5S3vM3Ftca7WkHiBase6yWke25iNorPUSsPmLFj8h
xCoUHVEinlBmzwzgMCqfnX3jenBhZrs+VP7u9a8zbni0cDdDGf2P5z3AoXWNJ8f3
3tF/TzkQSsJtRtHmoeRaHpw7CBrFHUMGWiq9NB8rrd1FPYKFMR4gPW6JFD4D8YSi
OIP8YPuFSlIghKOS72tj4EoI57zNhl5OYavOPOvNDuQlIW45304tb1ZizpGOJkzB
tbUiMGipblokJG3iqa7McDK1rs0acD8UCd5suHSnXT/TgXvyx69kE0d5VSd6bIu1
rVrzNpKnQ/KEkuzIGlnHOBj9iNB8rhHyO0TSKTa1Xk3Gz6MZREOvLa6gEzDDjPev
Ec11bjsXeeO+D+5qWltd08W1QN/fmmZwR2qHvoNY6Zzj0Uz8p1iWIEGrxNhw1YPY
80GqMai7/vUGIUPEgmesewugf4kezF27YPaZpC8nQugLx5A1a9X3TGbned/iInae
TEIuCFcZRFEQZSZa6nJoPk2xTc62HK8lSJ4qtTOdObFR5Eod5haMj9vONgeWB3D9
6ANTqs66iJtnyoAZwyp/mkYhd+sLN2j6Oy5MdnSACnEb0tRN5aeRzYk9cV2O7V2x
o1TXTfqdRADLyz7w+Stp8O0hbc7buMGMoL3DCxo/NheG3fIyR20X1gUanfj51mBx
DjiGGkeAb2U8zcVqR7fVnyxS9o8frLlh/IWnCGt7S4Xm3RusjB76mFiMbpO6J18N
ixAl59vjh8JXQOYuZdumtAmjShbK97t1IODP1Zk8OZx6mfwky7X+Tc4aluZgzRtn
IPhMGPBeYp6hDOpXFElG6gZWWlpKgHxQyyzn9vhUZJpTClU88FbOxT/9TfiqBB8D
KzTH3FaAptWIEf4raxLbQB/iRj+vaVa9opLnN82r7RIuYPB1DRerh9V7v8R0vIIH
Boalo79ojg+teAg+G58d0d6hyXSwQhutFc113zBxexSgSjUWUVTuvpsfEiVq7qEq
RwUcCdQ4ILK0Am/x4biMT4nC1otaNI322CADRm8feCAu9aXxqAsX8FNRFxkobaZ/
fBJdSUqoBV1XlPUBcEipHq80lZKJIWZOpmEdzveCCzVhux4ufYePCBLao394GYq3
1E1DfVXPO/tkTESNtyNYPIn9Wo/2dK1I3Y6eH9CGCLue/06MIXslmEnrZf9W80PX
8/Fs7Ek5WGBG/QXjSWL/6bjs4YcOKKbCbNrJ1eSCI/589ybADToHFtP5IyyvIpFb
U9JJf5sICEl3tM34IgGGNtW4CkqRQLVC9Wo/N4AS0SLarGigfIQvQJbDK9dX6VWo
Rurddnv4AKPe4m6kFcGDmikiTXGE/Z8r9Mfnc1zs1AyovrBI8M+ZUQ0OyHR7t6jN
SZx8T+OjpfAIFo2t4qJevMITLtNTtm6BLSr+fggOCo/wbldFCHN18HAqZXqNq6hS
HBjuc55IRMXBHVNJNugCCAE3LdK6DtH3do2fNi63C+RjIECmcknQCqa0zdI6K6GF
7szGKOWfGhrWVeXCYJVaF6TApTjXvrn4wV5ytxWUKK9p0JWHcLGBvGnKcANMF3U2
1rDu2ET+f0cEf7Ubbdc+dYvT3UMJyrf/3TGs8K+KIcpLlMzc95f9TisqSmA0L9X/
6X7pRzQuCx/kpwFhDnQ+fO8R45NJFuj0pNXyHoSfVFARF0IXUBuGUKXCR97k4FLv
EPhkCKfBaYZ2rOi78/hHtaHhyRBziTohjLT25k941bCVfGoiRXgJD5RiN079GRTM
vdlNDVseF73K/nB2YEnowxd+wi08dqu0qcw2w5dH1R8O0jOeCpkSqj7/idTir8wA
2wkz1/+tLZ8olyfL2Xd0OvE2/ZEi0nMIM8Qmtgy5EIDA3LO0JjNiw9QbcZjS3TCm
EJOD59mNMUfbuCkeNrQyb22R9y4CNeVLRABZR8XSlmmQgse0RQ7kKdweopDjheFt
z/+v3ogxQYN+NNZvhNuMH4//47xs3w2TEkY6Oh3Y3yK8ik+ZPSBUEddaJ4pzrQ1B
fVyXBPHlu1V9x/uLDwu3OOodEdesTLebYM6BcLrROissmP5aY/UasdhonYr9wPlZ
FmGChnqgCdSyyHbBOejY0qcuQQ2/18qlxjLMSiRs5T/yCRRNOD+fqIL7gPwVn4cu
0o856GIM5jWH8KfXt+MXyy4sLpGim2NU0xK86l/u9et8DhNjcqOaiGt49adCNC82
lwbIk7L35KYW9Ehm0JB0QnvC/nIlxvEOl58ik8u9EHt5WT2MAKIlRe8FHhcT4DOO
ICev568FcI3JOKdQg1IXngH2X3ckPKLtNtpGn7oxCZhmHdHChDptr/XJ+o/sai3M
+yHD7CkNxR7e6LsQMLz5nnZDQdEOL9qxXfrsWCmfs0hf/4ZsDsiPySbzGiq1pso8
q6P0PyA5cMb2yHzlXOxmmo3olKfPHWOUbMxq7l4gxF0XeMIBFiuiH+dTJ/FWBUjQ
+JumSWkkFttGnfaSOMgrvxMcMVCNoGz8i00QQH1BtHtuV1I10HkdeVXcCo0bhpJu
ClS9gmyva636djMcelagplKEeowJjhw6FiiVAk2JUj/rtHpf1Q5DEWpP1dl1OyzS
kvpBsGNQxjAbHiZ5y+/DwxGIL8m+OzGBZ5uiXQeYVAwaGUKzAO59BBvaICwE/UNF
VshKlElrD20Rk49UEbU7zpVkyPghFXT6yRuO922jiyzxg6XY0lJmUGz6K7UrbR3q
R2JuIhaWW4L1fN++Io4RTWRfJy9sCXoDIfOvXAJ5xnmemBjbveFr44LGnz4VeGNa
lNqNyO9i7NiBRvHYXDaWgJB5Z1d7DCbIFyex6T2/SN95YaSTD4DPIukbevbQUt+x
buk2QsP1VrkpYau+f5n1RRvwr6tzZ+cRvWBcAbAIJ9SNhTiQr7KcJaogoT3SX0V+
3/uH2f0pSYldk0kQLfuifntSRm5va7Cpd1o5IAO4Vl0LETa1UKdNJQoo2w1XM/Ac
ArTHYHLwBQ4HRShHKvROp7f72UoVEfj3WyGaXxJLRxi3keKXOdEXUiUl0E+QzhaA
ys1ZIyNTE081HGNYV3BjCHjbNQcQS47mThMGuBYbhmOeKXQsJ13XKKivtNwk3bJC
EgSC++uc66VTHw3KqBnMHGpINrvgAxTSRumwc8mb8qfa7mRz2ObCrreB289my3lS
T5nnxdqsYxUNq08OwNbd6whOcCuUCkffd0I+zK5jCJ2C/IShJl8K6fENVG7UZEX7
cvTZXcLcLDfoOGNf4CGLXZMjvyAwCqS3OUoPArzr/RmGN/CXXFGkH6oyVbN6I3CE
tWx0/XimHfh3hzeSltiKvURJTlErwE70AQx+G97Kn3Bilrcs2Xepq4QeXZTBDcWr
JCuCJdmd6tmbkuaZXTn5/XJT8P5dpVMWDJMtGMiy68q8XBIDjOsmNRh4w9hAEAQK
1Dreq5CUJsWATFzgSB7xIj4vEZZxfppTtmqZJPRXVwPtHfMPfUfSxEZuox6h7EPG
n0bTiam0bLZ8ERZ5ASRjAY6hlJz/OSSoPlWmpPQtRdVUu23/rfSdBHb2ZGes+sjH
BL+cI/Zjn9s0baMOao3CwrDvanRzf1hOeE8GhQaSzdsUu6GsX74SS/FhhQGz4MiF
LaNXeuwW77ko6qW3Y04YPNCJbqLaVLGYFHdD8T/3VGWVFFUZsmgRBVvAj8pR/y4A
+BArQtsRxK1csXdRLIUC6TSLBCPFhreDW66K46IulPANCylfaJ8PJZT5FlZ3Rqly
qipyESpiBH3WVT6xd60STeP1oEnw0M5002pR25Mei15wtJ3ZW0cMbq8piuh40H96
gEgq4RfblOipmMZO+84onSJpLgtz4eJytaIBSDOVC0em+D5+8W6DngJUS+GUTY6v
kO/nMzSht0rruI3JgtI8O+tbBXHOTbH70E7jUmUKta/Kz/Q24wjiVYP2RpZtbb91
vBmqgP5/sVbq6wwts41bGLRXibsp2xRTZ4dB4f9C2iWoWrPZrTV3BFetu5HEPmbo
R4mEMffziq1Cdvrtdcw9YK50fN1zLvi/EdIgEwIeZ4sBlAQlRbltB0IL9aVnB4gu
sLeWZUNpzuwtQclA61AfQlzUoqEVqUdMwN+Ct2G40KQRUDa/pMEN1PzMdJp6sJFJ
MmJDMxjvRew7MjoAOv/ngZjHJNT9s36QP4uWpJZLx/qhtJuPQab9xZf1sTNXIJZ2
PSui0ouM8hjnRF0pcMDsUoRpK3lwLv1sECHWj0+6ogv9UxneuqSJxWrrVOjzZBgT
poak99ij+bVRBVYOM5C4CA5lFfj19mEFLm+eJeZPZepk8SY7+c9wXo7W+dDSVmxl
PNYzW6ZaZ/PtUrPP4sFJla0rbcXfcBA1p0ZH2CM0Bjl3GxJKzcPVr0TBZDu9IzOS
mlymzyP1Qgg5YyErIXnoRGkeHbUEkCp6gIdatmAuumXfD3OCJ5mFsyV61o5dSSyg
/9u+bSApZMusohVJCzJjZSTBHZYirRVYdlLFK567AGpr1nOyrrzcHEtcMw+oDO9u
sfzMVbjYZyROYWKKOoxBj7oXv0CbmN6LyUZiS4DFvTLIuiugBUjHWF+17Oqu1GHZ
UR3s4samcG/Z9DbZIy2Wp2N97rfkKD5+QFGw1B7oqpWiD3hhzghcGpN7uFnZqIAZ
C1nEyZQ9GiUV50P5F6YuGn8DdGWx3oTz+Lc5btZOIvhlGqLdckS07wgmGRgpVa+/
uo9xoFRmE+GLoS1V92lpei23pqrmb7gQtN66do2pC9QGo59hqTpftkowv/9+DCMH
s8gkj3Xl+M+1G1VOr+FjBOEnM0dbSi+A0bYuEZKGWdE8/Z37PrNPHeDfJCwsAtZ/
Tke4shkUq0vpEY6AU4Q7u64YeUAlsZvLY+lymyf4hXLJ7ykD/WfzO1G5UJMvjP3Y
Oc2ZZjuhhhDh55m+R86d1Q0Lo/gTJo0mLiSOSolDq6tEAoVFvR1zEYLLmce/WviE
M/tMtU0LhXX9TYdNh1vTQmsgY3JRc8KbSOx6Qz2wJMu5lYVgt6+jJBegjbHQxT1o
cPRu83vR5RfFqLp02GNhTdcJMDLcHrbpav1SnRH5igjK+l5KHe559PDe6FqK6NKI
8oo1MHFRtPpDU5xsLBSXQcZMSaqKw0JlJNFpdwa3ZQApjMydPh/nToA/J+atOgwc
sjkzjU6MVeJ3B0EEULvI+dAT/UKg9y30LJLQPHjpNE8XFJLao0jCgr8lqjvP/ldB
c6ayhN1PXPHDzixo5x8QWTkx0ApyCGfpr3TiPeHKKupciZa+mCv32o8iwVW28AT3
Ndn9a2ZCsewc6JbTspco3aMNgivqed5Tk5IZtMOLnSfb0sGx9aM4HEQKgGBnd+A5
+R0FkWbHJOF/woeY9aHeZjpdC3FMXlgy/ejf/Kd1sGm1tzrnjOGETeXupNwARToW
2CExHBWsez53EjhXk1pA3b44VgB/oorPk6skI2YbBXq48lfF/TKQzXbuoQYyF1ZY
V0TTZCEUczfSnBWNh/HtTSWhqQnKdeX5D+WQ+q3apymEpgFiqqyIEpoTarJA1n4V
ItvBs3No5h6cD3/X/J3yfmpo9NVJTs2sR00CaFPNcWatBIp/x4eJUF9JA53lFT/F
LUfly82g6Q9q9pPyY2t+J5ts77vBNsV+gw2W1NNWGPnYMn+LfgUWQS6lK0P/OC1e
6AVsOigvRTY2el9Sw4O9l826xRqJHDwguZPXuxJuVCWhl+VSxnSxnLzR588370Ya
hUWR1ITfpSKM3MuUBX/bGP09UIkZnBClf5SzfBLquNyqFMCkxJmzfZnXxTUuYDvG
2q7U7Qx5c72jHDnm1fPfzHm/9kLbanhph3m+iIjE6y97VejucbulYG59fqVGG+UG
GibThYO4ybWEMjXT71Ovv7k2A/wI169dnel6LzibVkX7fhjnlgXWT2jVHwCzkDm+
dHYvmq9czbC60h6aXwNirCPMTnCIuKWOz76JACoDZLv/XTKFX64VYNiFB8Y9aKwy
wetF3Ni0+xOi1inltJJcgR/IielClETD1vRhLGq8Udx2Qec4/L1cARwbRAoDshzI
OezXUe7+i55+wyuqIPBD37GW5n7vKgUBf+3CVcIEmAPZLZwzBrcru8lvJW59QVQb
Vr6xBevv9Z3K276Hmrm7102XAcq2cOhrzLB7nXrFGFkRX90P7nOWl+wfTdrw0Bwp
AyiLhA4DIa6WLRj+vL90Wnwrho+Yrd0S8NSddFM4VLk8CdwqGMYEJ9NOS0CLSuTb
ljJcKUGNt1B4kjyvnhntG4M3VyAG8b3QZcouqv2wH+neLyidl22lsgC2agILhbtA
lw5TNDoPPN7M1y4+oMKC28j23I8A+2WEga7jagwoyzBrtJ4WKRMpDxegwmakenHp
JUjhKhG+BsOz+4pWVo2ia/wVnloSwbmHE3B0wX/LIaDWXBma3ubuH5Oh+Y5coGJF
ubiiymZchdw/LKJg57RZX0TaHUNdBRlLXPpsZjKVhlceW02dB3hM+mqqfLZdU1c0
xxMTxA3EEIPtft647xViMMYY9uMSGd4jI/ehymmjdI0yxLrP7EtA+Nd9rv5QZFEf
y+tC4QMS7hJn/DU3wtFiAF577A6sFdvHNAPT5ByktF5F1bwzxsV4e+o3Pjzsufrh
5fgbal4lyGF3GbtTpdR8GZ4P17RZYoeOm4/YDc6c68SdWz5heuNaUlpWXkpoRkBb
e0AGbT0THkqyqQLpvNosb9KtKNU0i2q4h210uCf18h1Y6wDOfMPQivRzlKLIH7Ua
TkkGBt5fO/ojMN1E3BpgkLeBO4uyfcTEPs5UBgrXUM6poBLBADPXuwXrlxzCl019
OlHBAxhwn/qZVpBzzARXfsRCKeU4mY+KmO6hRuDdvndOwzhDEeQ5qa7a9Fo5mnbn
oupKZ6TdCocU94P/h4DeN1XeEZyfDJdMmoQXosEktbdogGy0dtaDesjdGvIAJFYI
D/OvdWf7sDrkBnu/j9pWxtk4tXi3d9CAHIuvrtIaS2dYsnc24a3OQBIkUBDh4/Ez
Md1coobm60NNWMbiSMD8og3gav8Q3+Mi1pKs3hR5VbTzfNaumz/7TUNIp7ro5d4A
h+IBht7r6sd8I/0E7GtRmaujUSCSLLeX1svTGqsc3NtfO4Qd6D18zYNCcbra8aGm
KCpMKSxnNrbSvfKAJwVTqFaMR0TME4G7QWTs+XBXW34Syqxtd06ePU1t2WHW9sx4
Ks5Xg/PbWOSZulX/Bmh7gGsxeODq71GffEOJuGgx6ADBHn7IJMjYVy2p06jkeTZz
Ngl2XfBElOWZuIQ39UhkIs0BoYF3iCGyMeUp+jak4rXKNkejSWIpfzEvsJt62YD8
mI6S9yLXlZ4SE2Ay4wyzxge8s3rjgPWuuETLFJr0HxRfSJE9olJQY/zvk84bn5QM
ucBeeG/kP8l/JLWRqMnl3KM5J+/cGhCD8vTsi8bca/mxMVU3V/ejRZfaZ13RujMv
gs2RqUDs/MNGZCTCBqL8hi3b7OwXkSqlGOlhrwZmtKQb3CC/I7TEmtxsCKYmEarj
8qco26RN4avddcjdCzYyowbKMMDmIxttkKi/NHJw1TgFcUoWxMEhtJ4QaR6UnCA/
+EuoO/X9+IGqwC7EQORyyS7HDN2lHLqt47LHysUypiPGTXCzXtRwQ+hvMG+bFXkl
DkWhgrOch8HegvoMETFwb7vIIGofmYvaUqaJtsN7Bky5NfPCnHSwUEnr7yDSPemo
YOL1X0qv8eHTe9bXlHNbmv4wppJUaSYocdG84n1RO0YOVmc0FbVSumRWfOvoOsBA
LtwjBATFOslNtU7hzoI0LyzN412FJrCDsj/dI++ZAdB7+SquL2skJ28geYFwWkT5
uaKT8QFf01FRaYL4i9eINo4p4S+F97A39hnMWnZNatj6RGFx4avyUvTisZ8uwplv
b4Ju0TcQchM0bZk5HmJtuqzSDbyLBDqjYVG+lTSPknYy3Y5lTA9v+KHuNOA6SAk7
J9lDR8QSJDa6nDQp5TKcDYgS1B1r3XCt9OnvLP7Cn6PkTFFioLT4uAeAReYYEgdH
zkz7NYkBF6UFWYtJhMpowYuSq7hhfBIpjfL4QjkOh+rnL3SLu7sNCJuVM361Za/D
65lqBHIShIbvEvocW2fo/DYcvLYGrE1csRU/GpbF6jJack4R5okPG6jJnKGpD9Ms
KQ6iwkSLGYbs0vScLRk35HvErdB2M4QDiTrmzVS9BCAtFr3wjGjTImIKmxqp0B5l
/e4nBLJ8DcGU6o2qAcTQZ0n3UHGGlIvpwID+ucwKRf8d7l/lL1/9q54Hu3ygopJV
gyZ3Frb9Oce96ey/DuH5szhwDM1JQ/Eyp380nYO6iAUMIidtnbyHNPFAlOcpA484
r9KSE74Y0xZGMcb6PqEBANcMVnQnUj1y0On9/Ru1rLPRm/n40zaZ/AfTrK8XLP3w
YCiuGKPpXYfL8o8WAyM+HCgQ764leie7frWtx78heX2+Ho5ZDBp2pyWZfDK/XY/5
2HWSI2TjTss1+G/wCp76s1oA9fEeIypZvsuRBj8rD1DIKUS5cgmlgZLrPZBxYmNn
re9IqZOG0L+dfktb78WKBp58F0wBl279v5eXptL0e3z+nzKg8dGTM0DWnyUlDWiI
KGdlZOvXzZKLs2T9sBl1iR9gi7KCphVwMXXfRr4wskSQ/jvq/sf8RpupySOKXakU
a2dtnvF0SyocVZkcO3KHfey42K+fLc1S3QTaBMEyj/3q2eLBQL5LiblBlvQqJcFL
4vDaFDbK5nbigmuqTIlCxHbkhhaTc/lEwoP/bGmnOpmvxmS7zFl00KIAEsYmU3uZ
WVa5mXWBy2fYnrE5Nb2KjOtFCHpHLlyOyF1cg0Lv4+8hpW9C/osMknnU335q7UAZ
mdMqKqftsjvihIwD02oZvwkzHxNXr0sy4Fg99GeB2pDmPhvq+ouFF/ubSP+yPwSz
zKgV3V8HqKfS5NlLWOVvA+Sh/iVZZ/z05Fd5+CbHHcydNn5lsIHuRPkNqIyd7LoY
89g+OynjE2MDf2zTZNAjH2DWSS8qRLq4Ikr8NV/JAQ1xmCfCG+8XYx2TmE3zKLj9
YSdEsVRPA9fvh9q2pVusc3EAxRG/7GcvVhgQLIM+LnmSzcp/454vf+5B4H8EtHFU
jBMVJkpJ2W44nVvqNpLuWMyWE0dmQwGragYlb1/Rtly2pLnZ6ZYE5BaDBNUAhVz3
lKc49xByOWQQCPxmTX7maqXBZZwP9/v9g29hb7wq9R/DjdqejERcLjGOeIkRwR5Y
V1hnjr8Q6yWm4wDLeBYtHcgQWo+pCShJ6QsMbtJhMy+XLiwHEAvqL0DMehUjHb1v
ZVWai5TdYUerQoC74faIR1XqBgWxWHvC+kklOk57mGa/cimC3+DEADrQCAL2wDUI
Md1D4uHJnvlnGScPPVmbdrPSHuk6Tm8PveLYPxSQP0urX0iEzY+OVbXrVlSwxfBG
zsF1orwB/CsX6btDptgpDz0a5J+0dL+Dhw7MsOeXCF2DMyVka4tV5bHLr2RwNiTI
5nUM0Di3kj1qqAEKf1ArLloE8WRPujc9qjZKd4jUxBv2KadF4TF65lREkK/kxkte
c8hC7Mh/XlxZoLoRh+fP17FaVFAL4LM7RI5wQoK0hLd/DnNV6q7tXrWb9nLS4dDx
biKVOQ4UZ2JM9qcg0x4gLoVn5rQkVuyrM5J+LkpxbT+ga1UAd+wSPERA+FX3/VOZ
qGiCN8TrXfucHLjn37/2Iw8WloJPOicnXPHo5zPiuG+OKHhX8UCULg8L6ecgiPF5
9BNxIN/WluJ9tWFU+/B+qvYY0jX6+4+OaaLk/uCihP585IR1dTjguqmfwvYxh5nv
du05qqa9yrR7Cef+7392IsZQfzZPhHW3yC0skCfYXTze1j6KBBO5Y6BGQvCp5I5o
U2M7YC6wmkcj0QbycI7veaYZS7itjMHqKfZYNz7FXPd4W1OVS71MuUkt03s1rJuA
t/OIXiwiS/pR6DrKcbJWIQRlLF8FcBdias9CdeshizJ+M1RRHHSQUgFysv5yJCcZ
h+z9aieT0bY4TrqP3VOLLSBM+g46QPbDQnv3HYM7zsYA/eeKqQXVKjI4ngaxTje2
IMuQccIUbPn7VE60P81Rw6P8rN2VJpXLuFkiP56awnVyzZ6x3FqM48DS3ysd7XJu
604ag118P88ncCAL6FASFnM4V83jN9/O/liUacevsX1RLpTsQpqG30+4C/qOanr3
P77nq3E/Yxr/cEUOAFxUiyvrsRzmBIlLE/89jJnVUIro4lu0+n1dypmWBVCdw+We
YuYHZxzsJ0jUnp6acabr5sjky+KIjAMKgHLu2NeHkjUpdweY2dhlW8yAcClWdCcV
gGswchCHSPDj5C01OQDGyrRS4d3a7d4tsp1BqA+SqUOYVnw5zvfi/DXC2zSWjukz
Qxy1gfdGIWH/3pLGT+oPcLXbCfVEPNFNrmn7gYypQttZUFcdJZUOT6OpI5DDXxPx
htwV5cQ8QDJBcOkCiN/c0X1x2mgJuwrBSue7B5aL9EFfdhlWAqDUp/nFRRH0ixrp
8XdqerGvFwItz1txJLMVGnoufPOlDfbJ5sWH78y3qcKqxnxAb6p+NhJjJT0UqDOY
odqzcS/ZM+9s5DLIhXeEZkkjNf4BLScGsCIriJPbZlyP6H3n14OeXZ9iZp001VKp
EEXAw6tmtr+vLxgmCoodNQxZgl1xAGdRVhHfGJbPpSalZnBnT1+1relxB7AvMiZU
IraQUYV9xmgT01Sqga4UPvgWvPuMcvZH8rOolKZYH7ECMXpPI8zPG51Z4bO74HvQ
gvHCKL/1ZW3v8oh9T1cdV/Hyutos3AOttRiTsXKPWekbpxhiqXJIQSyaDsuPjhkl
isbictZCTdPWST9OQIFZRUOcgoaP+khr+6QpDRG659rISUxUSC4u7HgFOx214OUX
So7YJJteBu09UOXHM39cNcpiwLvM33dLBPWT2CqG2yVzF4VwRXf0mCuEgnkQ3TCX
jgNWn7Hos+8g0EjoiT0tlwKAQpFflKofzy6fOk72VJXGr/tFxnz23fU3CNWzu8EJ
3glvj0EVe4YjB5dM2MY8B1utL/V8XoJifjkPuXeQ8n+LJuBblwrchv2sEtV39f38
hXwtdbHkv2pKsv585hoJpiZ2uhqB4ARhqKVuJCSVww5bz8/lL5o0d+Yki1/3e5n6
bSVjN0lp4cyj9cyJ6iVG+odXqPgpZiMsodpfDiKVoEHFxtFV8tMjuO6r/z7gk9ie
Hh3ZGiXBY8QA0hYip3b9dGfvA7yskQCz+uSTZ42okPVzICWniGoww61u5mV/CtKV
LZU6Vj2xfPpd0nP1dv7hRbXVTMsi+eb9MgXTABGY0AlJH52aOFDSdSluYrwx9wuI
4EYF81mZMRwMd9S2FaLQtvIOD4eMSTe60vrfGsj5VsvuruPRJx52T6lTVUDRPJzH
40AtNzrETbakwgsdn7dFD2Nx6ZdW0XPfYIGk6Mw3YBhGMorbkspQsTXVsylNUwjh
Cx80D9Vn6KS59lpfwnxFgDLhSszGWFRYLJ/D1M+/h272y/W7y4CjX407UGb4r1dG
pfIkEExDsBf5MjfH5lsR/BH2959bV3fLqHAWUP8W5KTYUvhtVbGbf+qB0h33qlA9
I8P9gboOfn5Fva65R01MnlwxeEZdUAq0wUzbjEjFBe9e0kMrKyCFJLR4C1qyujoN
lKSSS3gpupPpVTemMS+Iunufn5hf0mZHM6niAYNvdmnfgWKpLeLSDUaV5clZd8+h
5//en72ROtP86mQqC4iEt4T9vJV92I3NKNVw1jZDd0cFCwRY64q9tiZIIFV1AEMG
kn5ILurGRmZJil9pWkoWMDKPqBpnz9xVKh4z/2bJpEV5G+lmB7btf7txxKTGVTc0
A1QWVlVUm4T6SejfQjvm/uvsEdU+GTao0X0JKQwQQS3j0ygA/9VN4hvnmxy8p03r
VN9ZrmZWKIMd7n70qfCWJNOldcP23NC7bUR6oZ85Pn58VNybjU/iiywG7k8y8BND
kz7+5IsIKhELq+1Fqj+Nd79wDqzCnq9DN317uam0HN7ZXGWcoQ7SkBgauG30wi7c
/KzKKc8a8NPfV3ogXefoFXVEuOfe5lfQUCvyNObiffk+gZHqQTFHr/xyi3a7olcv
fgOC/Kmv9oDFJTcFHMmb8ZkZ6SXaR5fQWTyikvq9jCuBlKMJTgUbi7ZCUavkSAtQ
oS2UtCSYPenVElfBvf1cDSenjDH3TOa3PU3ySCOwCSHdongumiuuL9Pc9VS6R1mG
7RGSGoIGDhqM7VUEJkgPKmx5U/vsYJIoMvvXLY7Fbmf6a2uUsQPl9w78hEpuVayO
sxkOgmTnP/4yZbEHZr4c/TLJbvnTxghIZpUW7dETa43HcefnJou3ynyNzBEjzAeM
/rG2DqZk43l2srxwtijkPVmMZZVNZnIhzOfDZ0FpSKjzGDga2W7oMqQFqTmoLnSV
bWRit4rPyE9G6bwTsOr+fjegapFQPTPvOd428fLWWQUIJm4EIde8SrKfYFfT53bj
9/vf4KZHbzZLFYKDeVS9JCrARaRGiWIcxG7LDqG4kk5YjTMzlRGftrRPyEh9fuCh
3HthL6HrT4uHJK50kQimLqXXruIag+AJymFrKSdSy/CWY4CvyH/WWzKi5os2z/q8
NTvPND6z0ehjOnYaNjnR2NmffW8Ci07XV+si8+KX469qkrVTrZ2r+MlRepEZEMn5
hIscIE+0e6zCx8ieygi3Q+rF2jjA8vQNv2m2HOfCuLZRDeeH0SQCJVvyhIflOsGM
tnzUuJabzL7dpmNjsb3xcQfWkfEowvDi5JjTdWhVa8RfXtsUm5xiXBOpY0imkkTA
iaELVhlPL8My9g8ExOViR88y3xRBj7b2YuGzs6JkJ3iEgqR7kfrlt5BPKIpK7cA6
LyypHq+Wks8UPe6oyg6tG+FdwsIUmfPe9kFb67WaFvKg+OK9tZJVa/rtnQyq4fuu
dOkLwD703OuxsGuPvTMuB3AUUJr9I2Pq7W2/TvWvaemoHdjZVGuhA3frWJPBW5dR
Tj6WPVRX431CDpv7aokRoBp/dOa7IfnWOxUv56tvuqrnMU9EaVcCZRL0hP+XJH/D
nyKd8eHpl+NXbRrFs2iv/ZYcIu16kySgx+cJfDGOMuyQJiGr1jVNaUeqJUqyHttu
jT3iGZvXnfkCLOTwqqd+vY4XX4KNQx8XMaLbISBpH8KbJYnESH+GnbM6j+2RD03z
eTlz/wyZiYW7GctlWd5d9Srcc/r/QcHqGOAwfDaDKmE8Wx0u6RQ6nyM4DZmMFP71
mmvEnN2zepLlifZd9WqUbMWEO1upIDW+Iu5cQ3WmIJZ6lpyTJe/SftqieNqBesmT
hRaJ08+kgZMwJbU0Ij9zQfnCkZUdCKQqgTL5pAuNCtLamD2BCG0/L5VRxBmzU4T0
my/aNyBDmoa7PyK1DQih+YRdBddcs08DONSfNWqQYAIJeKxJeEpEWrPY85Dbi8+p
kLW9NOkDusBAWSQ7cslx6KGRbf9MrMgbNOkeycYDkG8lOxbxyDx/FTrTIZNK20n6
Ylxaz6ff+ITgjaJVdUkbWfdmBJeqHIEXHIqWrbRfrRLUGYgjtt2ognRfu8zt+737
0V574sTBuGGydp4ewWJCHlySwA2A51fnCfWMzFQRfWCaJ5UufArUr1xo5/i0hx++
bQ36moxJNq7APiOXp1n428b3O+zRItWJknYrwDDl4zKU1LIpYzGaELfqgSRbQLeK
rnaPfJ06Yd2k3QlMVG2bWbqcsdYCrKE1xsEb9kPszaz7i8LFOQRmj50kvcjz32/s
5ESZHFoePqoAMYDKoVBTZKq6OPHysP4VL14E6FWPEp65OswDoCd6iJ3tn7B/JTjt
HOrYD8QqwTbpLxQyMVsZNPn71WGVJdzdZc6lW2cZDjID3x6IZZ2JFOr6DwLTWyJe
3YHtHtDgzMHHVbRrx5ddl75rILPOvfpc/OWrc/p239y+GMh2QJSPawpE8czkcF+C
tmzYebT4EaDxKVi1sVj7efASKdOVfZmJSJlzJL8WLpHvCLS+/wHRME709dBuKwvX
npfk6I13HhN/hGOtYeZxz0wSl9VBKrwP9DmXmLJsOf1EHfL2LnNNb0uE5GgOoGSP
VuVybXavRtBuwcf1bWsuk+vBYNYFR7Q24Qvf+yyuHqd4J3qI9DDUgqb+cwaFEqoa
Zix2W/JAyIuN1evegbRL20p8YbnmzgHZBXlFLhW+EkYKzKGxITPjnW9JhZxAB6S4
RctIcrqZmBCYGrTNysn/ONzDkgMuY3sN4KlZgzKU3pUdDB32PPHloy3Vi3wbTOQN
/ZgKD5e3Tpk8WsRQIg4XK20u22ez89ZCdNTDL2cJ1Yje25XEsu4hXf/0T0okMZha
R1ke5e6lqhwl9Ql0swM8XCxaNRA+bhnPobHRLc/oK0q/iTe1qLjXnLJomLgZAGv7
QfEjP5RqszYRGu2clBsyhNNNeV+poyS0i0vVnOrxyyGCzRSfiEfzqHu7zz4dAEui
4s2tmmYul6JvfmjVL0hl4eQ9W7zRcFvx8UFYg2ONT/1yZuJ4WuZYru+mWOzTgs5+
hr4hGRVfT8aZtNgHsq1V5E8NC4OHUzsj+r95aCGbyzpy6BUhR/6U0vfhCKWnUdKg
LoflEUkXU/yRFa1iZGAyFz6wlFRAMeRnQh1xzcL2JQ801L5NmqmyVMmJoIRW2+dJ
QOfXjxWXbZX8egxi2YcI/VhO8ZrqEqDxUc9GqzKwUsmkbPdiTuSYQpMallnhWIVd
OE4Pj7BSYBZAiCD5cxTgaW28Fk88SmhHHiYwJ9ccGbY1JwQwcnAL8LPLuDR2cptU
T+DdhwgbOYlPB92yMULmXH2Oc9MqCRJUWYnh+pJEB7nmEaJUWmobQNQVSP0avsk9
AWEQkcdE2Ug88RvM5Cq1KHmh1JYeFtkqzj6AdTDzGcs+iE8wtYdE8etphxyUg+K8
TNmO7yZvDwbeCcJczr9ZTrZBxudK0/7Nv8tWoiYVA/5xetFF+IXHNcZIWHg4oXh9
Cry6+89hjC7HJ4SRZ//KJ6414Sx/0OguknOIl9x2iVcIOnpHH+PjUZhXDqxYkxh6
wdF6sej1x97yn3FZ9TOdalIYfQAmaKRmuj4IlKujaRdmbYQmk8vRt2xxAVM58CTc
Z1x9hGLPZboU3RZ8UCnadqxeuDWBfdYCrI/eP1Y7YfHd+dtIqndIlBV+LLJ/8obv
M9rtUuhkoklcziDLQ2SaDTztqihFAabX7pTlz8mC7Xa2enKnsMFG603HCloX0sn7
rSDNYkGDyaEtfFDbFcl6wuVJLTx7RfmTZmz/B8NgYeEQq9Up+C8xoIkwW/lKbA5/
7rXZdyUS8tmVM7+ndiPubZOif9ZRMgLeeCze+wXKUIyAB6b/P1rH4cEhsN521mrW
m84Md5L9Tl/20j3vhr1VANM7Cwsb9QAHXEkFnKOSWrBs6sOS4hp6hSitoBy6f2VS
+HPnk2x/YJHxvVq2rTQJ+qcNaUFhUBh5xWVtRC8VVIXtKHNfAl1qY8XRYr5PkJ/9
QxvMjpaZI3lecwAQQmw+F32ZB3AeHTWCC2qH0uJ8HlnYLWPLO5ydXPi2+wzqjLVz
kgp7/M+c1A8elDO9KAFAFvdTkbfhIpsAGbswGZzE2e+Qfczkb8SeUU7aq+OOnwKe
Pz7KOp/jsM8c9IiZ75HvgjXei8Rs2h5dGRxPept98lMYFmcLuNOMDoztuUaXe4Q2
9d7PC/vw/eT8DPJejluTq0nhzpEJEqRAAsfbG/fxUvqnb/W3U7baeMDsEbSuYG/3
fpBxZNL3ZAop557/z87XHL7QvQYt9ektCb+BFv4Bz+FFrSylhefsLEdnUm/ZJ4Iz
fLMvScHkwwD+5paZQyF+zwdiWS0Tm8jy7DW+7gxIyBlh4VRbufnHln3t3GOYIab/
qhAP5H+MGlAJkRzZBv3CygtSbgMVVjpkAM7mgKxh8Lhx0xZPI9Lm5Afo5u+zpEzd
hsXDlc9MUdDt7ewlAP95cGbrmuqyqcQhP/dD/c0Z8Xyqi3mZ/dZVTm5Sj58t/Md3
rypb6FhzTu6gmUkDM+A+ChDatmtp87wvi1Ksf6Lia9OdZqQnX5SwDtrjVinkglDm
zplsAQCUhZIuC86RVr+LnCXbmTSt4oe4WHqbB0tDw32FW2Zsac1bbw04R287tt8P
gHjU2ROhvN9aocRJVal4aUH9cXIYRNiQmU35KPTGsXY+33d2IhxlgbX1f1U2Z9t7
GoZIT5q+1couQ+bEEIsqI2X30dtzfAHia7L3LdcWw05dOYfBpb1X2MfPwLBfQW3g
RbzopeLcTRIV6mbW747fjB48h6NwKg2WLMU7WHEtHrUcBHHs0jBq9ZTX+8+FCR4E
sGrbR0FInZwHPJxUh+xwsiSfrUE2OJjIy/NqKBPaRkkr558ZsXP2k1u341OgiENU
EXQoN0sL6S9x7/e2BZk8Y7wZ7QTMQ9ygP9c0mz5WN4kDUMWtLtx86synXJh1WN0a
u1CgBFgOTqOsZY/fA1/SXgcdYni1jcn0snSJ8MN7kslJmzBtWFtcsFzMlxWqBIg6
MSxK+MSTpif06P8Nz03EeuIZGb8wlU6HeZXDjJAuQRVoeKokgLjRc7/lCLhW71nD
1xXpmUEkj0kxdRcwMnat2il83FQmeqSKrVfvuu6QYLZznvC2NjgnGnL+x38KTmsO
lbai0mBgcAcmQOhkUd70rLyK3DU6kClfOXyopdSUmI3D+Y6MDMUrISSLzzH+j4BN
HUQG4YMfXefFELBZQLnjVPOcHkTO1Qad7cj87kIrn0r7O1PSWhybOMeeM7++HH+O
zB/8KcFkStp9MmS+oVXlvzRck/lk0hboq3sDBPCKViBaZl3gKbnU9aNfL0VW69Mn
UT47gZ9aZKbHDRQDG8bNkGiF5+5gH6Yq3b5Ip4Bt0386Y/eXprotdPEniFSWQ+hk
H8D7rxpu+S5Se5IF36xvyGVPg7HpZYP0MeXaDnEhhzFqO6HnSOI8MVF/0/RKS80y
LDsCYdQel8ISkbubUCUbbQ9DFAfcUWgPJHPxr8YFpd3fdkqAYl0Eqz0op+08Q7T6
xyj5gbG903L+3dhZcQZSujFry43U+9Tyeh0PNyTmq5KxuXRU1igiSz+p0WzbrULD
OnpwXFTC8aAHd1tgGDUVKI+xftJSOkEqfc7FZa8KSGG6puT1WiBU42Fp68JhCmXy
Ieg/WZxhxWRSttiKZp6UFU0HG0CMGNBtqg11XgOboeVXa7HaRxvH1ykavrdbpcEZ
4T/zs85iD6wZ5MeOC7O7uXykxQFrxaQpPHr/ZQyVzrYGzva7KkX2sLWrgeqBl0Wo
/IlUsTUYCDqI5mlEdK0jrn/otUB7EiEepP5X2Rds2ltDBFq314Z2YxGlHI/nEgyV
P2V9nOxgWy9gvfBdieayJTL64XTLYCL7ucnogOEqKLGKKk9WR9qPlPS4M5je1h+S
3zeTmrIoZ0G4nqKNM8aXknuj0uEavLvKxcYLHPTyagR6CwNmV0u+ZYYi22ZSp4Nc
Y4zEye4nzmCi96McevSOVQZ0G3pgHSmsliSFOwhzHva3YZBhqqhPxROCKAzo7qZW
qvXXSmM20fsHUEaWao0ocSIlqKTsBXT8M1hM0A8/kbZcyxWwDNXeT5szJEHBcZVm
jx+2eoT7dPypsG6+D5Jf5uHtHfVO7reKizamdR6joRupW/XwglBUZzjFtSIREhSg
srcohplpyrD+HgR1mLb1f7C1yLJPQpx+JJvweESLqJI4b3yHHAmPC78SZbFmDan9
icITTYdl3cTQebzOVs9+WQ7Re+tH7SLOnNLnyFmcGi1qklvjwe9TZFlnQ/kvhe2I
QGFjuFzwM/kiPGM/pz4GaLFPPqohGcKpHOLj8DE5413eMj81R8vB4obTUZIcmvMH
EVgko+rQny80sgMOwS7OIwj/rPLBQvki5sBXJdLCFl2PmX7iMTRySJgb5x1eQsCe
oWqIkmtaGk4o/ft3XmPhc4hVFeMGwWAyW4MkUpctO2/gm3dISq8P2VWwkdjLXB31
sXiJ3Xx/ONE3ulLciKKQwtg4hBlsZw2Qx31epoyLBp7LEmDgPSFFwHNgVjXwvltX
zsKbBg2XEQ82fiRT70lqXHZafAHO44Y58IHVXo8UBTJ7o4+p4PER3pFUxBEu3YDn
ymzMjXf7bnaIM88P212gvjund0ZAswRRxdSK7BC/yZqQ1K8uMTjx4UdOoW8s7+xP
ukUkMildHCZj/qFKr46GH13PJfLv+FaAhWCX5aqLCgA5DbXycwgI8CISZnP6HMca
FXwV+KW2dSVmidEHzwHb0+0XHfMsVHrA0XtJZX1/jr1HKfkkfFpNJvVXhA26YG1R
icLVqkapZT0oflEpRVDj3J5EimkBY5mK75ZBQ9aVxTdGcaUwEAHzEHpRiw06YP1w
hLrOLM81na224+U+MKs9yhgVzgT+YaR5unBj0ALTKgccuu4NHruPOPfIUy9zbIn2
vvJh0Vj0BHukupy2a2g9ubPmwTKJCYhJJ2dV03chVxuo012BFrLkD9PpVWADNiGX
nlnRgHtJezi3UJEbJHYFLaLGTyyLnIWbGwPqQTBoPwWpAhPHqJWKu4Qes2gu9mmg
Ei9xP/myz4+JRLvPmMn4uWz9Zhl8ek4wye99QNFsoc3zWaqXsc/iaggXMcOLRO8q
eXp4/4HB/AB9jODv1k7qze6y6ECFszMjbVUZbUXxv/g9yv3c0t/yslXcEavHhPWJ
UzyDGEMhsLM3y4JWQ0xZ0uy3n5cPhvb0pDI0R3+lU6VzrxAYie9B1Luvz8uOZga6
wTjYgm4/iDCcEbkOypZO83WfOuFo3o9gieavxtP83P1q1hnhWt0ygaZHWBYJD5Ox
ayV4j3KS2Hx7tO15Fr2NuDtdUW+yCiaHz/y64M4d43zX+/DrXr/39Y2IgWlrtzKw
pI6b6AnW6WMyJEwNemiEDclu+fpluL34LRZ423EUN4pXTpYdAMk57qJ1dDcwvK82
Zsmm/iLReB5GSatj7CKd9+Cc9731TQjNF97ulkq893wtp4S/SmMzqBKy//3Z1HTL
xJU2MteD3AamgJy9pijSGomG74Nr+tHGRdnqoZoUQrRMlpFPEzR0czvwKVisCsT4
XMuXXxXoAIxMYBkYREVvsJcg8z2sYDigcqPc3rWL4ro8EZ+zCyMyL0mPDpOsPeRA
vzFsb5slZZIVVdXhWMCg69X1bOA/agZJGU4qEhAah4+HomIO+uyJ7UlvAxQN9+kl
jaN5YtYeeq5Mgz0CnxT2pVz0o476Q86nHqyJtnU+kEoQR9exGgaBqT/d3E5lCzXK
4jYN3Ip04M3uuKKmu7zBHWr66zb1dpq7pASkpPl40csY/52LWyCtGs5SrJIt8pNT
iaGqIZiN8yw+bqAa3NgmZUZGlQXXpihIF/cGuFIW/lgbrMJkJCrAGgwt4GnLnc3q
fUuSpSMjlWjDTTmXnTFsOXHlyzpw3+HWvezf38ZOkalvqxy3ZJ/ZArFnkX2P1hG5
gBPBcln5/N2ut5FQ2Otz11xw6DlZu8/ejWSfQVYHDvEGHG9biAVB/0J/B+j/Q/9Z
/XBYqklp63iqWkzMaEC32iM1kfcR3kHdcjtXKZH6c3+UaWFx8upZmtN4XCEBAYyT
Svho+uoCJkLiSdBBf6zghf+Voxo2dmK/Ot+NueVex+boQJ97czvQKJnuhLm3r6D0
v/pxGyX950qJxwIATktwjAF9S9nW+sAKTr/YoqQxShiTh10m43xi0moG6DqXT0jW
oyWzMFuDRjgG99TADmOBAV8t2nPG0+AqUnrrh7gFggideY0pgy1Zfss2ZebdZXKU
xO9TyyiYiBHAN/4Q1oMyerQFDNbwpNs5clEGzoDcuSyPI51ETa7gpu/VSgcr9ik/
gHWp6kx+snBsh16v8ncCsKZ6sGlwG2tLN++pwyXyMl50ohcoTwCpFkXl6XaSopue
KUyXYd7xoTyAVI7JQ3gn73FYZHYhLNyL4WxJl9lPdyQ24F3bdRONL+09zjqLS19w
QsEbUOGV66f8rkmtcrc8mIdZM68yzJ8mpc3P9MGXavaB+PHkEf6oCx5+D70dB1Z6
2kc8UMUDa5N5FHavHFU5djHGZY4jv5GMqugdSO9xhxnB2h741g5bEUotTk4b8a6x
qSF3r58Li+CW/+ZV4BYH1NfBWubKFZqWOrQrazRaT4Ne+LaH3dSjZaSzAN2U5x9e
s+eQYgJkoHRC0T420iGEY5aNGGjKwMOEYTIBdUs4E9p6xAsEOAEmeDiL8FZF5oea
/Ooc9xcopbACcgQTVewkKFo7kxj+oZMlQVcIpJRRAtu1UlZ1YPkkDNd/0ImzfFIU
LuWnvP7B5Cdz7HMWwh1g7l7F/UtRr4wyty67RguU1tRidPHA+/wNjUqZ6zbbDTJe
TQwGa0O3kXt8++YDh3OwMbUUX4vh9oCl1aurAtholXdhw/R7WStm76AcjSFudcNC
cQXwSQc95n37kPc18RySFVPaWVQ0vruAUlucC5dU4u83yIRbo8LhYZ2VAMflhhEN
jc04mqGC3np5ku4Ms+KGXy/p6yg0RxQ6beuGZCtr23mJ1qptJtCCvUbBlIzcH0FL
wEmS1ukVSzRq5Z+nWbFUGCSJuPsISwnZVmt0HABCD8sbSC3QwozjOoijHnt3R2FF
5NAh4xdDISoklHAk29WrQJ/U0L7ZvgP6sPr0XzNC+YKBFaLBKoFrdc30Auldp/Dp
5yXvCHwRZrMJsN4IJHJ8PsziGNdAJmXvTtaoP/+SoRmfivcI1FY/XEJ9jztqQy02
EuiGErREMNorkHxBL0qwMbbnoi7Kjf+ydK+TVACqG4uKilaFbz5b1Y05gRrrQKy8
fSYNjNTUbyI7keNq9rhI/akUzo05L27RNlk4g5/huGxPqxsv7GIgKBRbFAZhEwEi
vULbHT3hy5NSlR7JjX8KR248cig20MAoc0HH5mUn6vS/fzVLiIzYAfT94akaAhPW
coQNhfnqSZkJio1FNby4yeOtSsqWEOak4gRMLek610aQkfXuO5d0QOPeY6u9EjnM
zS8WPgOR9iTqeAztU/wGy7VCIw7EJjjCD64gB3U+1uz9yNOgu4syhkZTeYaZsRBU
CKMBTWa2Podo4qvR17xQbSxN/nDtFUBYmWLrZtM3ZQEVOBiJ0EAXEKjp1OxG8haE
WGUQ755iJtusSz3kx1lyVt3ADpkghTqsLqB/pPbej8yegwYwoLqMPHhhdqHz7jTY
VhukLarJ88JZxXtBtZj4Djfzuil8YkPRgDLH8K+3Lm/nUgBLMvkc5u9+ccHsRRpi
zg8OndgZ8k/Mc9nMej2uO2tBnYjWQMBtN/nKm4+AV/zjGc9wURIEpsCUEWgjQ6Mg
zee4N5qerkVJRuFMcUB1CG7ns/gwtN8wbjC9ojDkIHIQLJ5/LeGvy+QMckr+27Xq
MrGU6JwBIEDl5gB0GUPXI5CAquUCMD91JvpBJmCN8vyiEs4YkuA4VhdKX5YZmWyi
1ayea9rGUI3mB3tmUtqsGpHZDHiHWBXhkiDEQc4JBTnFYmYo9pU1PFHZzneb1yBo
f2JKJ6EVxVHRjwkmJMkvqDVlgfa9qrZG66WPgmF9Xl0XMB84j4QWyjINjKXWxu6a
StPqHKEyqjPk+zsTo4pU471QL732/NF1vZjkjELdJQ5VWX+ryvpKBCdjrof5N619
kUxk0dwPR6JzdezeGiL3E14Qyyt4WP0Ialf3KxAoyD9LwOh8f2QWkHFoyHjXGcFi
YIm8Oh/l/dttYGceyRKkcjRLyc2A7OVYKCnomhwolZUy9sJDZ1/4V0NZBcpBf1QO
duS7mbdsoW72fQKpbVESZHol65ZRVT8PIsiZj0tV8mAoG0l6gUA1Rx1LBYF/1xKX
uS4Bt4PFKLlNuW3D7pbVu9daz664o5AoyY3WFAqUw47BkYlpcUTesjpjcoSNxOOY
FMQ/WmZZVmmHJxP2+ZFY6I6NeBircv9Uiasg1mPqVIP7hdoz8VgQ1qW7vqny3JeF
vFe7h4veqTNFnKwf9kOgiltPkbk53ukJdGVRTW13Lhk1ZFtrY8F+qAl5rwLtpoA0
NbHUgHgKUzGWzvjtLccMOPmkSM7qG/IEPdKHDEuy6Mx1VHIto5aCyLe5a8mPr5i0
ArnQopnmP7aOWow20LRSPvU8rSt9D+OOJiyIUJE6Xlq7orfxmo2eRUTqijupD8RA
qKPS3R0dhLyN6fj0P8S71Xk/24wlRColCMWnOHQb4CmqKTNt2e0RwO5uAKB5X60y
qcBH+3RAkTHYZTZJGYjMnrqrQgq7Q1r1m7itdUx6OTcOhzN8QkJZj85ouir2sVuC
ADuq5Rf0a8DvAy+g9F5r+5wzrSWzA6oyxISJFWkeqxxgoQH/D9o3P+T0cEkON0ST
wty5gI5LyrOmsY16Z0TTkQw2GMfGGodTelFzLxbSLRyFpKHJZG1ZNzPB4ZKt7iX1
12x0eNO7ohYYsWNrLZquhSiJQKh8/RrfGoS2rCza7HrJYVzLfkMiuKSe2br54Kp8
qVQkbgrMcKvIh63bp+LTmkBI4HTHb35cGOf26bwYxk+tTzifPfaTeor3xMdDJbu+
81PvmaxnR8uI01i8W17f9Vl/EXwBUdIzxYwuZdD5w40ZS8DdKfBsxH8HGivHuqKn
ayFL74mzjPRFKWkJtm9LSSfowmSAywRt/A1vAw8mUlEfjg9jxJ4Kd6WIknw4V9z/
CjoQoprBOXtO5py2mGThdz+bUI7bg3vNOuunQmNoZSrnrbw0+ev3nJoEcYxmK0ep
I4NG/58UPHOCT/MoBjNZ0DFGIgqhkbmGw0+IrFnE78TIpL9j92aRI/rPUt3NVUTK
tziD35G5GknVViHfnvsQjX69WRoprga1aUvnsEJmR1e+8vcyKBCfNZYCtb+yrgIq
v5MZRKY0YgSrNrwtPCdylKwaUYUrTQ6CR2HvxvZemZA/EvKFOvdqntmIfO/31Xp+
xMLAcKA5KBHl+U7B0bLv4a7hJBYpLH8ZlDS3psNvJM9Cs4dJe12Xrq7LGyuiKZfB
0UTnlt2n9QQpq5gzlCBCbTPrUrpdXcURimNIaOzj9I5PRH580UymdzqMgu5ZPUmZ
ERgwsQbi2qaQ8i0h/btyYJ9xrPVqoPgnqpDkNRUKiu/L0KpbjslQ3rFgXUriAwrD
+JZQfpZANKqN4wGOPcQ3Vjc4Q83l3yryMN9cZ4yrSBmCfo90ronBDI8+zkl7sJXZ
pDT5HcY/hI3MVaXppLAuaisadVNf+3X4mwC4on94xCMC1icvQEtp5P7Jub8buQrg
j+9VDmph0e5iuVzeXQTdEpKD/UjxXtZsZASz+aIoJYH6nAP7wxZss3o0zzbrxLxo
B2AP604pmibTXFjNlF0n9yjjVZdInVvP+zMqUF2gcf2Cvh3p2ilQaK8rlZOq1/zw
e2GffoLu66boRjGoJ21e8LmushbadkXHshV8nqpuK5AGen9Pf9xq/WYYki0i8JiJ
7yCv/MdjATOlo+/3vRVp8TeD/PGOb1SeQUWDqreaUpKwhPrwwfLHU4Qwr+knMpq/
0GQLR43dxrOJg9LCmEEqVzEnG9esgGJEjQPWKmEnosymJW4P3bzzJg9Kcr6foGDZ
ymBy/gnuY6kvoAV7f154Fv2VG6VZdTr/lQDUn6UQdW1nt9QOGsGsS6c7L2+bxdYL
7wfz9N8zffDiCVNlQ7lNUuK4QHrSgt0CCP3ePSRYGW7xkbCueCHHrCv2+787IABw
xP/397VaxHPLgPPsk02ChPUMf+UyglkG9zZA1aG1kHe5TzyqO0DS1mF2egBCI1C8
zf/8NXUWeN8dRhajFJkNDSsvTc0WLgFayGgG5eLGneyH/Jm7BCfrBRKxCRZCokjs
SDfzNZfxy+IEjqYc6B36vF9eea+Yl+IjUImxq8WgVe8Su5k9oOGHSdxM7GmdyEvu
0ue00BA3XsXKvrSEj26zaUo2x2qdFqdMXNOOsXUmpN52ky4M8vQcB7ESRkzRh9dg
3DHX76SYJE0o9mwnXpEh3bzi5ikoyPOKRgs5dURUQyG81NvvtrN7p0U7/KwFP9Kp
F60MI//+HSKuHAom8f/QOnD808MvQSytRAq9YyHU2wdNlJhr/SdLd0n6/wLllTWk
/+jeQgMVblG8CwCK2Wkxy5UPxkC81MetIBc//0D+1p9wmrbviG34D9MLNmsj6GOB
GU3t6uzvknSPXVRitTMHOv01dsTf5JZNoin9Il/Y2tOttpI09inqcT50ljDolQYI
VdsIRas7aM8OcBybutZjHpXpAfMPVntwjR/BhXfL5bGmtLb9RjZTk3/Um/Tv57E1
vGEM8Y6CRkJvyEGTDWPYxFFJ1tx4nKmtZxt5Oc5XqwxH+uMr0k7cTZPbGxPrc3qV
QjbmDp9FK4/JthBmPtvvLsklpPxHK7abZU33TNKpZBR2JFXJAcGHQ0wgasY5Ge5N
Olc6yS+AKomBuWaLvwc6FqLXWcQvOk0Pn+Qk7vvFt7HFFq/CPXkFsOtajoGz/zxw
JVStSWHn9Mq+PfXMxVXKeFJ/4oqjk7o/jWEayhJ14jSpFzdFrydZeKBS1+hvzMyc
fc7jlqBIiEpSJEVlWq1MerGJhBcygNmt7IKfN1KA1iy/gpz8JXMwIvVo3NvLSTyS
Fj/YQ8O8tWcj7efsPkQfpmZb0rvOPX6nGqP5gONt4RK+X0j2ymwbjxy0d/QSZ8t/
EbyGYdRZYiHk7qtin92wEFQOwH+HU9sshPV/+Gc1fg/gHwy0DjsN+46DBLE5sa9d
AiD6sYb0ppUkINN+S3fLrncLAYMCc61Ab1lWs/sVAZ1lGnIupV+rLK93/Vx5lL6Q
wlLUTdpNkI8QH4G1GkyA2Rk5Ob/h1WgqrjvTCUjRcLsAU/Aj/GJ+7YC6KvXBbaAO
jEykcJCXEdQTqUypOht4eXM6dN0TzVJb8EPs4Y05wLmz0/Oh3/3lBOouRVvKQivJ
bXb0fAWd6hdgpGami54DMPA4H4ykFNbyjxml3zsp/Bt+HQD4yY1hEVGnw5dknYfo
PyUbiGx7L1IaLDMOCFzDOYISfk8SF0502BUzI+N0M+5UZGxCcTrMV/pwAWL34YKy
Ly9kuB+O9g+3xmhB7datVqO13dCuRmEI0Ltz2FIV98Psbb/9yelv8fsGDsg9ab+g
Q9JUEhNKHZbPl+TyFqczR7pnwxch8C7JkCMgUzDcghFHAA2akyZ/oQOJMMsNkx0h
vs1L8b9oP3QWwpDY6obcyh5mLnEdaRiik1yslMPIZlXro1KLHT8MVY5QorJLaXZc
/jEmVhiyp3uQdzGALlGRmek+PqR/s4r7TJTUsEqNzJumkwg5bTPzj8vBJF72UnEY
BMPyPqAZGyDAT4nge1wLRRycBxC1ycvMeibNVEWI3yUglLY+F0kQ8TX2yYZk7NNE
zPRdJGAHxJ4FWjr540pkY9vmcTaBEg5Ouy/4DsmGPg8h6xnHIY1E4kHRQiO5ol7q
ZzZLioNO2DX+W3UCT1CPPGPchOohvOxUhvT79jSAJbUsrPhYn3iDxPR1NPTXmg+a
d4F2AdmXCDYLr9AJ6r/Os1uQX/0KtmvChWlwKW5wAh72RnkbwfPPwA2TGRMCYLBW
tmSGtdkAnU+I+L9N9+UrZJ9LOMn0Mho7CNurgHf75ztHbLkg8Ct8JjDEw/jb5J6a
H6WCYZx0SSj3l/yU98pUGA48ZQJpMK20AVgyNQCFBfpxJPbpPO5onA7bLm11apYi
lkfpyAjttVBxR+Mk+Xj4qqAXy0GYwksODuyjjcjgPodAukNgJI2COLnGp1xJXDo8
2zW+z+SDmTtodl5soHxMnLIDoXDbLQ7rfTYb2qeshCfMcUTNVLCiLneCUJPP+3eW
LoGOBe14ep/mIxW/X9GPXEz9LfvvKz7okByCLT0fuyd4Df3PH/qMZ+a3Mu5JpAon
z5ECmPHh85YtcFncLk93vtQalL96+Y3U/yY+K5BsF27maWuPUXwl4/N1gLCVburw
nmUzM3ziBnabxMtFFxUaQAds0LRT4mqzme6mqT2dZNsGKnHAvREtR/a0KbOhukqz
UCZgF2w6vdv+jMEOAQcWkn2wIafioryf7RYnRsBalMiERmSfYJBX8h417F+G1o/5
AlPxfUEhXZTnttA99JiFxsVN2V0aUQCT6SLEuBbwD1lRvAaxts87dnAnM7i/aIq4
BMUeBscnM3R1fGJazwc0NQNCKfmN8znHUe7JS6HfsnUQVVWstYBucF3ghB9lp5rY
pkCJfZop7hOoxm9KPx9Tmge/RSI0nS0TJhcQJGzoNMY9gx4Zzac2Gg09y0Ex1mtb
S7XHaPA74Xyev+bX+0IVH43VRCFkbtigiyl7lpsGAyK+i3twG0qReoCwhg6xDAbn
cUJ1v2Ft08IXaTQ3vGnJ+XQ6nTYUU7QMiF73++FMnri7qn/+/jFHOFKVyOShOF0r
liZHuvXJJsmYNjwppJeKq9mdmBlYI4Iaz2SIggZwZdWmgTJwpuvFL0CCyWpqhp9N
/+e39BKTL37AUnw5CB4Lf4ddreVsPVUo/mEcl+RshYzFIEMoEoPUJZc3alPU1SWJ
n5HntdziPPn39tyrymiwiC2bIRQcWoOKezODMwMf/79BRGmTpf8YesRkCb52/Tmo
HG0sFPU+o5j3oiZu1YB+o0uMSF3XbLQOeGmZG+w8iQY4gHcGKvlDIJ7MGfY9GFgz
gtDrQrLbxfn5aXI++yFRh7/MzBNfKr0G07BCpzE03d0ylZWv3lRk48qawfYIIlh2
vrh68VnrUcPOZ9fbfGBRudKM+zb8IaDAiIIhab9Zjr/JpLb7/Sabr6MvrJ4DF37a
rvQKJ5GHau392T3Seu+Rb4F04D4FbPh14k91cSUH6vYq0v8BBFWUpoi8wg/Ar7fi
UMDjgX0/sJrTK5tbGO7tfP9okGSszXC02dSIkKWHMXlzMGQRVHbhgdL7ddmI+gU6
72Ms8oih5aRACSTJILc61L1vR53RHS5WkswpEwHDLZ4z7gWqLIv//dZieBhZEOZU
06nuXRUBs8psWgH5i18iYUqbgkSK9nePFemfdDS/lVgnL3K13NUuit+y+VPDFvad
WqllNQeZRiCZnpnHSolsCyZITBBakUEEu4QzO7r+v/gfL7PjI0TpT5jV18SuHFrw
3Lk3dyGeUeP+0+rIuE3R6d0HGsrIeLG7VC09xi3q4FTPhFxFYu47osYRuvvATcy8
DggtOYceX9v4PPb9qFWSaxDZKMYB08C/Tcbdjy1mqRofiI1a2+RXbv5KKdVlDrvm
sI1ISpJZxb7D3/6wH2xJF+Z5GqsbdlhigRgsiSjTFthz++l5aoZuxrbNOr5c5KVL
5RvHJ6ywusvzkEzTtx5x6EVgJNU/Nv9tOtckqsqXAcDjnBxis1LxeWwD4aKpKG/o
2mqYBGRUJHJxvaqosiTcRqpeCI+c7il8TBzSXdUWQWAa+3H/8qAuIR2EHrnxhpwY
STu6MT+AnlkAYxrjv593DK5uWk2/X/kT3PFKoHY6ijO8l4apFOC4qrVxD7aKWlkT
qdr62VrK4Dl/ETdMi3ywQ5hkoEJqntr4u+OoT6Pzf0q6xNH5ygD2rPKWcjrxMNhw
vWHpWZCmvlOJMD1hfcjzIm63C0fTJeRKNXZiUFP5Ft+3OWN0WhEBzZ0Z5QGsJ3UP
FKQo4BsZ94Otkq4Ib/WzcDvDxpAOPiU2PYm0ypbbbsqPKi3AYm02Edq4Plnotv59
ZJgVkf5z146PDoerH4IFj+Wm49UiYHYbLrziZPspLuFDRGZCHRzA6jzSwwIhnh+8
+r6lLntzZS+rU45PpqMO5MZfSoyKoM3iX0Zu4MMj7EjYk2G3oB2TJwpAH9sFy0Mr
bck904W6PSNT6UDBpJkar0YeYW2MCoSw2gr14aa/F7sKV8dx/XiMgF1yl+8r3K+t
9BGRnoo5B3VRfRFB2biMYnEg0Rg2EyqSmsOl8zHEPpQeoaqys5/5kdcSOFJQ55a+
sIAPMBnWF12pM7EQs2XM686Mish7VQfR5bPHjN6YtLwqY6eYoE5maDGECFdTGQrL
RGnM14AtOxoE0I98UEbbdOPwSQstnp46FDFbX8g0R5MkI7k1BoTLgxwS26Gt9I6t
W9KQ4fpJKKztpCuYsV6Tik2q/XqfH3S80888Dlg+c7fQEDepps2mf5vAmoA/HAZO
lb5RBVfQ5ZoI9HOsixQN+GxFol8FRe2976O3huIw7j+oFCxu7ODX4IldXdWPrIng
gRjBrXE/YQxE7JnoX4IH+r7qX2JApAHUu/beKpTcU5mjBPfS+XotovgXL2dzM7EJ
r0yTmoedyHuRq+XxhvDRCtx0YXQLJngqzEZ4IiFID8SWQcPEYmk2dJ4lrY+js92F
cwDkUUkEyZlW6LrhId0r87olEXb2DPjdCk9O7Vv9vik90lRfDxUYMekSbAkZlGfw
6bOjLOwSmwFsE6LqkhYgen3JJiCnEnUwJFG/3mCN0NTYOT9+pyfW6g02LzU48j2K
9+9UN2LlWDlygdw+umGXpiGLiTL/dbNE/NutmU8WKmJxZG4HIXFQBSBuYaQa5eH/
Mw4P41Bxffw4Dh5C/K8zyYKA4jlBZa5phjp7K7qZx/s+hKcsqRGj3H3i9OF/CWYN
SDRUA+zSp3v/xgl+9XXqollBnGs2P5AYPmU6YWHY4TRzrnI1MnxFqEd7106IUwE6
iozOdcXbXScOIjN2t3NVo1vANQqzYyZu4GPniIJAKBZQ4w2HaVwY990tCiddyQfR
7kMkq9N5uV0xjen3+v20K2X7pRph7JK65zNL7ZwoqOHk/Wp1YEojxfQjsVJvcum3
Y/GICq7OIgkTOs8siigmXX1UOQrHAOY8kat4bx4FjMTz+Y8H0/dO9sS2do+dkHgH
pawgxjhMc8dtw3RV6mRny1cQBhB2Qv2ygi6G4ro+jWt3AGgJ2ejKsVjYTm5yzRKi
MqKoD+YTkWGT8KP0MjHRInp8BXp2ZYKJgQGtgEAMub58F3azAsKnAg2D5XMysQlf
tG9lOKstQ7PwRJ/ntXO7jn1/KR6D7AXvhIGCxAuCFltzvudOwK6NZ/SmGluJ9yaT
wxMN5GBOzLLKGtlSHECXCMX20AtDcd3VSOlt39gULPgvjrd+Z0VezxNv+XB1n+jN
LXA6To55U6hTg2xXTDudR277klg9bXrPyEBZwi5Wc9hE+FVVnwhn+sFLI43va0+u
OtbfWLViIV01RU36QAXUhihyeaqDpbEVAzRLsZYWuEYrdFJPnoaDW+ivBFgg0+pF
yLiYUm6xsvAhYkv9SzoaOmRstRDRw5Fl7LVbv5dydpmJF9gYN8wExdw6nq5wji+2
tYxubcGOAiZwnYhpRSV48FYUvcTVkHqsJwZTZ+dPQG1PEepuy7+KSlclzV92lSvs
xpfCCPpzvF1NGdMsV695DoggQh3lKPgxASP5zv+mGD2lQDgVm+tj+nY22eMDFdRK
PTMHJagEvdsPiXYgTkcrnUrsgaeW5QgdmbHqbKg3fUX5/PfTO+NmWDkkAqu6RIpP
B05ol5bBV7xb++DZsiTpWdOTFS/+UbLC1dOGVzwmW9tPCyOY0kCqPg5HJ2k9okkv
r2SGfhNZzTTbp5ENmnG+xb92E0jrlk5DbrMO6sGUeAxnH1KhkQ+0h+CX5/DmvtBt
poOYuF/7JTVF7L260Cl5/Uyx6oxJ7nFsrycDSDihaUYurUhfdQ05YqW2taaua1JB
rLdhpj71csK7Ro//uDvaZR30a7zuo7K30EMPpirmKrNGPUZuv2Qn0jQ4nuEblMTQ
kRavetaaRmXBLwbJnkFdQpIJ+Qk+8vIiP7+gHVIMHjqgcP6Hb3xJ4jNqZFHU3s5b
pKeRyy7skzQoE+hECs1o+EE8g7Uf/sCAM8mWmuMJBLBrwIG3YnaNkoXF8f4GGL8G
gdAlCJwqR9MC82IlWXFRblFo9fzej7yeAab5rpRTLWgJd4Qb41xeQKxvJmEiATGs
dJTLggayCMvzgRpW09YBZVXhO5X/1mO4jpN6wpKSzH+hxwgL2nkDffjtGERRG9LR
PiUdYkiq+SgZ1w4HJK3UVLwPZpvxCNafQm+cYnG27kgTMFQ8SQ4+ubX3hD0r5Nox
PFNy6XJgRixPym9hKubC53s3FPA/HCTD486Gd7t8invtcq3g8wdoMnklLvdyDRo/
TgYp7O6P0yHfxrfOCDAp02HHe5mEy+Fm4L56MkKL09s2Es3BKPCiqgKWfcw7EeCV
1I1P3coGd55DHL6mJhUzsVHMZIGwK+uCYfrQa0xffSVpMnY2XjGr8gG5jGE8qAM6
vqb5ovv0iJN9e0ScWItBxB1SLABs3YtoZ1uajvBSBn8Ps3h22y9moGpaJKRLcr78
ISbaOFCM7OQnw9gZUqjNMS3zXl3ZtSaST572l1XYMe4DIUOQSLOafk09OSGK54r0
8RQJ7VijJQTJjv1JXks1d/nogzfgEv98f5ZkO9XvO2jviPH0kzM0SB9UF14N7tBe
bZwbdRt79Ku20pj+dYosibTX7JvAHDAKDSaiiK56Aqbql3vrB9U2e7N60KvwhzfJ
qHiUIRRI5QSQzmfmabkFNO5maQi52oPF83EWwb6VpNit9FovZB/bLwShVAsau+Q+
y5FTbH04SXgZIGwjkqtpqk7wLnnX5zzY4G1cuzX6S7kBl4lUaRBU+p5JSdDlT2M8
B2Fy4mz77vLBbnezlIL4xaexf5/zrzaiju3hyQJkFtm5yhFx4exvrKfidDRGXMi/
IkdX/jjCDznuHsA0CmRhADHrUiKBhIKoJzk6uu8R0qYoXvWZvoqsjFfyK5k2U2AZ
EeErBP+6syAzDNNrI8G7w7iD+PI26NyJSJzCJ2phsFYzDoAd60PiutlVaGCx7WGT
VGom35mmMCniru5Ui3zE9nXwTywSh2WVCd/VxWPK1oPFKiGvDFdq+2ov3Ofz7VPJ
mE6Q2tipAAmNIUXDForaYYJp8zATjfvUwyBGqxkKNW/nEaY1wuMBS+lMgmv/gok3
q6o44eiPgXSokkymcRhYOCT2wi4pJALUGwyeSC6GZjSdPJWkdhbGADOZxD8N7O21
8xO+Z/y24mklh9vlvVczzqfJ1oicvPqCE9f3DPoNEIb8s70eearX4oFCOx74jqcI
8NGzev3ikDlBKw67j7BksX2fcuOpFxfpApwZ9lMTu2poudfKZsMrBFJ1edntdhoy
pl3jaasIbbw7UDEdP8mWBr/IHOTHovvlQFuGjGK0+m0Cq1W5QlwlEq+SrRbZ3nPH
+I2UeYsOsVDtcwBL/SL1pSV7JspLIeHvmsLPg//SgLOmKok2J1CxfNxBEhH8Hpz9
bvZmNCRNwfOh+CMI/hb3/aMoQewD6/LldUlsmjGWZuO7lqoljl/7OoHQeWKWGQ93
j63BgTv7WLGiFGQrGyuN4UzH8ZaQeI6RXTZuAoziM761CMbmrj6UpVWk5IvmGl3p
bkHyeYilOkMc2DU1FTBtxGVKNnb92u5F9sMD/2EVD6ZfUGrGIR/pvf4/oNUCrUz1
32iTz8PUs2Zb+fWqHR+64wa37HvQ2QdgE8KmkKUvC+hxMzuJzXsP7cL08ALYHUb2
HalcLB5rCx6HNTl9cBgrDhbHPzRAjvaocuvEXXrJPVdPrH4sBb4TlOBVP8Uu9P/L
a9d5Y3otfYR3BoWLZJaVgk2JkINCDzFDPBlsQJUc+IfbZH88uEqvd145U3qnkhF8
LMBeofJYi79y4UipKSvdKdX2IlqLDuf+cB70CWNNgEAVyzpV1ZWT593WcvD/FGSL
vuOa7BAIeiUD/7JEiSXM6kn4KbVTJhnWAUXhJ70oysq9iZf4og0HGPDzCkdnRrOD
sHKHevKWucaQ5ElHTVkHRrl5UhCLb3qk7iqQRFWs6ubfncIuSRi39lFRUWwjJAq9
v2OcQg7cb1wMUF1U0qK8pceyp+RDvnoa+DrjsEzAf1HyxMHs9q3/i1hT4l2aGWl9
RtaRy1K0RH5dANbjYB9suz12CkEEASvPGs2kVpKwV1fZOhnm588sA6+8Qo6JPzA0
TH3ohXY742DGgr+854Tv4sPh16hQ3cetRdY1YLidPbzW1H2mQcWfbb72QAXZ+VQ4
kGOTeeOB4p0K35eErra6O03BXZVtJisarnO0dEMal9BKynlvBxc7JEKdfJv7L6c2
0oE9xcpAfqpKyw1UXgT71Q8B3EjesdZW8l/gOp+2ONm45E2m2KaZu9nrpP7a9FSc
UwMEr+QCMvm+IeMDR8zwZKaDMAYPM2Diw0l0cGgfIOmDE5Zf9YNST3mD3puwc5qZ
bpvnhMW/AP722ZOnz9u43UQLf0PMpCN2gNafnO7sPksvkvPGadxDjHokonSzJEyA
wu4fG6SQmIfzne3nJtCzbFy/FB8xGbhBLd5eKNWSlVdAGjOcOSuAL7y3DA0g5puq
QDpT6dVrpGxmdidc/OPRiAYdZ1Fhs5TcVJBMaGcYMJeZPtdy7GDCLk8JAmPRcLuW
Q94ejmkuEemnx5Q6TZc/FuXM2ko8gR7Y99MOuwgin/J2mhD9rvwEv811Gs2omXBo
ML3Il8qZvLRV3QK53OO1bb3QJHlJeEJqo8+tKRlJiQ1Bdj90uGsAj8wugIRpHIlC
lsUml9zGC/7qGZIAnL2JKUEaaHeTcJ/FVX3EN/8j13m2z+hi2q00ZXGzXAHNYCAK
bJI7EK6hhaPAbaBZa5WE49siW84B5wVvtSQPSvni0UeUkb1ODWjd4VgLPDZd2t5/
J4uMiuL9BHVh8U8RttzVbvBAAM3omnWeBg9JsLSNHSAcRWJ/tyeifKYT77lqi/OR
5YV6Bw+uJFeHLETz/cr0Qp+Reqifk7/5KHdtYe3IYsQb5nWsMIwVWRtWOiXCbn85
yaDolAES59obaB93FgbD+O6r1v49Fh6CvktdBHN65LmBnNhtO+kaOkg8Y/sDysbZ
5A8xbq41QHPIPHJKLMoHfc/EtJ2ekPZTPNrwdgL/e1naV7uOoOFnLMTxW5WIS4kD
0kGyGVTsJOYz/Mg0TlLKjWLlCUJW/VULN+rMfmOxgAHU2wYTprnSTPqSBDr7iGjn
v3FG3uR6hG2WS4CokphmsGtkw/wGzyKm61c9t7AWvomU1RxmCeVgaM4AN7z2uFoR
rFY7Q2JvJScUY8ce0HMTrmp8W/Js2DOprQvfZJJTPoZMY5wZ1D2+xi7Z+cwveHNj
BlYYYqr7LcOYrHVynyP6zEqn5SriKIb4B+lE9UjrCPScz0yRM9RvBM4ShG47slL2
HIBQncr8ogqibRw+66Zgj74POvyu0eiziYTP8/JIS3JubBQ46RLSck8loP0OOxBX
Q4oLt398jPjySkiRspZm03FoDEQawDWYJfyeRVWn6Y9JD6WpKBL0qhy1TKSHquWR
8dSTSiRe29UD1QPREsbfNoFD6xG6liO3XLmUNAmL0pGn66YrW1ZgKZ3uiiJiQNeX
+7byYMWPdaNG+sqTVtF8NwV7Ulo40h41P1fb//SjLpq0gXOsszugvayVxYPr+9gx
bq4PloPjuMwd46qD/WsH9LKMqErMc9McHnUg4b5sIrnmExkHJoZCEudFPtt9O5+8
pqhrlktH4rGbYxuu/pct+fiLBQILtwPRk/y6ZgtJjMeCTq6/+7khhsY4hUZ2UA5k
tkhtOiVC/eHThMSfwMIiJ5KH7lohkRJGAsJ9P72JaXy1cBfMXJm/CMAdZpGlKbXn
fzDX+gHafKN95EMuAOQUHxaS6Ig8W21swF8a1POwqR2h0PMaifDtdC36fxl1j4uB
4vnItrLILNyIA8qmLbhet7zckBBBHuhE1Xb2OzggbPfeOmlpoN0QmY+Vwf6Na1qM
tqCe+TvJ5RbkNFmZBRECTRN+h5hzyySR7ErYflYkUJ1r9Q08/6k8KrZMx1elod/w
nmMaZA1WhgKVowssiku54e+JaOJ+uIqQkFZbpaHO96Kwwigz8Wl0YGWMdqaFECHv
KYnrNrQxvmxh/OaRVldtpo/mrNoEIsTkoFgtHpBOmwUHJPG5ZG8rxXPRtLFMNFJl
1j2Xy9zebWqPDSNGJp7RxoyrEX2Nn5KAjOFuGflbCMA+OEeDP2GuZ9zgqdrODSQv
eFUTUJPqYwwuiqjXN0EYrxZlvzL0uh08V6ni18bSaJ4Fs7eYmduNTnhla/Kz69mb
exIsU2XjMRpYPF79ULLSpqP5QfmjEyXSwiJ1Q1ier2/sKiOMtVMZklBwLyT7riGG
4KPX8nlZMrfuk/nWZwsBSJoq4bp57uRODOA9nGCrOCX0lyNkTKvvrNvWP52V47fL
BFCNZvZb3ztY9gJuEykiGb39+Q+WzwHkddAPX31KsRYCny6/SdqKwLwZLKn3zR5o
Rofm3RQsJsZm7uFgUpSEWLkwMS6xgA7mRQyzcSERAtS5e1sxsB47As9kARMoKDYG
DJ38jZeoPJZDFhtRAU45pQ0mcz8vHX4BXlWIpQdaKaW0xD9nvlJ9K4OYjo3XArVW
8gi8dEIfziI45me8ZrziGx6gMqIftU0qt1pAWCEmcRglRNp5TstxYY+WWVn7KfQ/
oUx/s4ds/pey1oHPzBQ83TWnHvK7PPt6T3zUhIF+QqL9SogLvCCo9DVnjOC7tk1i
ZBEcz6b7P2t72u4+pR6T1EPY2uHhpn2hEfV8y51Rv3JiWt6qjGwNOckbkJm4+gWW
fiMihYXxKYc3doBtR0upLD2oWfS9uQtSgZ56ElsmUTVN7dwMM1pWfAhqaaIVDbrU
M1GbkZrlitFn/bgqumtqPmbnOOr5a72v4BucgHwbmjKnAWaFE/BL9Qo7r6Qm1LCm
PBPNTzVBWVG3LKg3Rn+bpu6cKOCr36ui1yCS14TBg8qbArpgZMTSaS/m18vByVX3
qg41ioJ1xY77WJgO47JW0dU5Gh4jMCC2umWRh8aavi2vP5oZyGe1MRjRgXxR/stl
/QfpgOJ1hbIxbfiT4qjvqsUwzffGzFw8Kf4vzfmpYztAm0+gkJXZlO6OjGC//ZmI
P7gygkDsLVb1mbKJ0AOJqGdFiYiUhP78kaZY7pkKUmwABG3mplew3vsXE9HAAqou
sFSJBkotVQCakA3ZfhzNAAgMDQJHqW0+HIB4C8LmRjJq6xzRw5sYMV+v9nzSRkIb
9NrDV8D2+/oJ/Q+XXru+PMM02d49YZ9VHsBnxHTE2C+Daa3Mnl3dvWFzpEZBJAxp
8+6N993R6XfE+fgP6KmDvLD8/1J3pAfwGydeJFjFJ31+ALagow1/unBGLFl2qBXY
ZbMiBtskXaZ2klk097lScxc+zoJCxBryBYoLwNvnIHwIPKagW/TOlTfT85VPxzAd
EDlw7sIdmoyXH6tbV+0FhzWuoaQ+DNuiOdyH9r7u01r0uQwP+z87xruyuA0G2o89
lDvi10cEfJmUh3248r0eHUQKE3qG3eG2uF9b4WiHFnnvreA/VIqobsEcsTmXdVUj
0dO/4ha6451LTxoUWwtDyzT1HsvYTEIJdGUoLvwI5jk1KVcjpdouuc5lN7wFJ0St
Dz1nT1SUxKBpcmHHAxhxfaY0u+G7/LLKE+JpQvCDzDEuSqJ/SqEwSnTfHsfTx9ST
BZ6hik/JFnqpAoWUKa8xAbR5twEUlXSemsYovr6gpLyHKc6dPMXir76ftug0mNp8
OjsmPJV5LoqrqxWICG1r57GkBy19v58E0NAoSnew2cCSIO61SDaajI/cnZA01V8A
ckvEYbAjEtcGBUsdEr+7IXpa5hRt8zCrXOwXeGFunD3Z5WmGFT40SNeBP6JfSlq6
YLXWMzsFIbGWWJcb9VwdtvKQ+HUZ2TPJxYpEm0ZYdSkEcx1Yt5SVfz03Ftx9yT+3
qSCHgVRNeALM/6Lu1kaMTDc4Ev8De68jd+OU1ZjqXo38XGThjdneggpu+GW4j8RI
W5pzD5YNrVx6CAz4IYvlBcm3+GjFwJ3c5jBcU11X1wrdrLtaOBkkmgTyRGk8cvaG
HRVBFAMnAMjTgycP2YTKNg19x0sx15KnYc2lpUN4hPKOHCQv+fYhmE4oRdG+30pM
ALw/snCGdshreqRLbOmVjtqsQfmj4npl2HSTEXeREVs8k7FiMiYQvaIAWPrA9k0i
XSQGO3ANyUR/XThXXGHgHbnov9QciGbnkyXE+unO5awyZQILfo2ourTCdzoTJPvz
xCQunz6YACVMoXlzoJdehR1RPsXXX7RsLFNWZvw27qHIdYjF5e2on5LzdCkR8/cP
JYytsw4b86HBElmI5IYD/a6A0QzrFhfhQ8gg8dGcwwTb9nP4NiKedmDnfH5QnMOR
46Xz2RqjTjcoS1lMlNqxgl1cjb7lssRHa2x/ovHHOVGWf1HWYNvyTv8n80dZd0f/
pYlj25NJ1lhXBwkVoGNDdAXk7m8yjjU3vTeT0Cdn7jRx8f4vH2dOa7RwN5SABrAl
3Buy4lMBZfr7K88L/T1NIjy6hdhGgw0CDgGJNP/Of8QXmD6BUTgu07Yu4MjjJFgT
DbCe3gmX87vF26rBgHnAWs3CTH992HS+HMNg53jj8kw5jEimA+I/n2+eq44mpBvE
tgHAglD7kDbeTzRQbVvC9zSQGoSt21YdVG9QLtW0QIsDQ+s/2pXQFKa/uZPOKt/I
qhkHEONC5bVuOIklYOjBGlwG1YamvNf41uGdfAggpM+4vnl4pBzCjRLxcVRTjybC
/rfuq8DXR2xM4nGwBoNTKjz9cGAQyKIghajKarZhFbWV8N91yI9vkhMObi6ttcq+
W3SEwxK6PvG18O6bJdL0orZS3vtjPySJ/d4YaQDf2LGQAMV02tFrSRRUMXUw3Vyw
rgEUGLCeJfnqq7CbHRsbuxnL/tArMwi5z2dIckUYi6sF5Z5mpm0YkAKiUZ1ldnik
zMZdo1Ehhrg0gSqgkgjNe49mtj5haVv5D0Be21zPGLfoyIDxbaWw+CJT+0M4DIFA
EMeZ7SO6QLGczJyiw8nuWC2+8l9xaJtEzs/B8LxzIuTy+grVTwCTjg+uchfMM+wR
eLG0Zr1Id33nSiMtg0neDCcRnmimEsdLKlm4s9PStJ9k2pAfkHMD7JIzfEz6wwCA
IZE69i+7wRUftK23WwTIDc0ktRpmmEKgoC6sD3JaJ+jYBpBzqQSnS4Kj2jgiV5Jj
D8E7ZhX4+RBFbpgWMfKj7FghkRqrFLVMIirBeEUlFYRvjTGJOU8qOuHnAg74Ucln
MQR1eajm/v6JhIAFzsdfor6iZvxRgl4d6JxgtJMgFqH6gmWMT2vbVyjlPoV4YdQe
HoL3WfDgPCPmQu2IjwS3VMGegg3U/djJEaoicNd5TofHHX7SK96mUFbtZ16ADjcR
0aBurzXol8Pc13arsfBHe29VYJvV3Tp1TRgmWnoUhtyXrQ7JNuqRV8k4TuwHBeSl
EvzAH1Paf2dNDm02QTqFpNja2qCsbse2XO6Igrd/9AqUQv+2llQ8ObAyxIJXcS+5
HuL3BVtwM/Z9syKVKCmCaqPHn+S8RprSp+OYSvVH6hiCvYVzNPCEDfUiAMmWE3GF
YPwgE/Eu+FM8eHqs8YjHPC1rSGiSEixdt0SfdTuPOvlmQiY+u8woa4SgszZZXkYf
4CzSEhNS1hAK5+eY3aWq31z3nm4pwguPs4dFYyXNB428A+PnZUG/+k1ZcI25md+f
Q58d2bGryn9Kg/p03ladCnICrM3wJmrprFLhvUhThBx/4JMQ53dVjhSi8uN7YsIB
5CtW9MlsJGPp3QeilSMjn6ZVlKHo4cctXcMZn0M1CxBGqDC/BTudlb/bXP3b2MS4
f+SMnfYIvsOO81FYdsoN0O8LWXCwMTbZjkuHA3/XFmpObwDM8UElVtXWrBofUJmI
4F4YxFO6omhgO5KSBofHL+X/kxtbiY5+1pDOrXPLCAkmTvL4SORX8gnJq7QvsRX1
QdVFIni2BniOtmGQGvJxI7+01k+ZGTgDvbSfeF0DbAVfQ5v5/QEdyb9iJ31En6Ol
k0W7OMaCe9rKi9lqkJHcjm0uzz7+Bz6dev+DfPpAEiEzT+gEyoR8oMtkgMOHtG/B
e2+P2reauP89VO0oaoRS1qink2oflfrERo4KId96qNbYDGQoOyZKQS0k0D/ug0pi
ZBrW9c4aDl7JCwfqqmSoEhW7QGG4TLBHkKcnTnRP5Uq+PMUAIRwqI22CeSjfOBlp
cx/i/qCJ4Lr1U15w1e5HwWl/3jt+B5J5JFhBEdIMNdUDYOnmu3+2GyfuZ1KJp0Nv
EoYBs2qu7paC2ItCKe2WflAxPXu7j4lGvcz6ZAmSRgh5JRDiMJKtPF1sGUjjizh8
tRr9CQngGywJso7hW6wfSR2hwiSKJIV7Sr+SGQTnkCBbTS5ZJDNkfS0fbo8fTakp
EhVQPAz/oDWmxKwus6vPr5cFhdFO/yVU9QR6UyFz7cUx4xJWfO8aLf5sfr40N+FW
Ag/L3F5oTbvIMlR7wux5LuRdno2LoQgivlpptI0eAwYp7m1IDnKGwq4/OjoYubZu
jWZbpmnfrib13nOU+eNTshc57uDvZ0j6WltXdBsTLKD6RF6eCI/0uCt/ULCgu20O
qOw2Sa9seKsKNugmdaIUaQyHlBReF1HOgNkMy+cdvydgHPAXe8nnxr8xuPcApmD7
U4yyEoMnS3kumxSwYCVxwKvmW2jM4p7TxCzyeLx86LmNPMMCPFm6qFUBj0Xo6EZP
DiM3NMnFphqZf6caA3V4RNR4PP+ToCnu0fwLq2wt6hqXXV81jxEkiM+jcdSx3PVp
oM5GanvErdgS0Estxn+wYJQNCzbDeXyaOJkG0ZOlYs6frESTDqVKAvKN44+8hBRq
UcW+YnsPoiY3ekJORnBWzV618jgE4CpRoIPsO8mOHxwa/2MgnXFYF0e1ygfe5obD
wUacWyNH8Iy4byNdh8OFK+1eUerhmxzekZ5ZrImJw+xFYLMnpxDMMCzEbAkiK1Nw
KGpM+qFt4tvTMY/hQoULdUpPo1Zcqfu/ggACJgjiqLzq/D4tDMFKIU/8QFUO8Emz
Pz79HeVMo13MtMAMrmXo4SWjdWhcVbSl45vDxiwudqNvuG6C+ki2bQ5xHbS8kJrp
ZY42A0cxjckRmKzZflPziyX7TwPzNF6hifWW0Gbx6jDkEeOjOpQglE0wN1ZySGOj
N93BlLjQjg0Kr1cdlQqBI/FDBT953T3XiRrtcbqueb3nJRnsfMRBP1aUZjuMJZUT
yuTI1NQEX+YRzFdCdRgChwfzW9cSuWEcbAUgdz+9wFJZU3hErJJMmmvRtw3g9VA0
Sxu6Vz8uLIEdf5oMcXTHYQsiRWhcFHqkWpEeq/uOOHV7ZTMuJbfhn72Q6WSOnYAA
LcZMPnCZAnHlS6Td+OJPIiuzO48YfmQBLIuB4Tow3wuehyfcEJHxDbEfrQZkQcVd
Upq7mdJSIbzSiRHeMfRF38FkSAB0YTjekqo9SOofSwvO0nkPm9YigitTsCWJEYRy
BYXi7y0jlcLz45n7KfsTIb4WTcV1YNgnUzkLNevgSMJILx5IvXKN0HvBWZUVw1RZ
uHeiWq/OZUjtoc3uWKhTLZ5Wt6jO59J7HLw5ThuFaAyor4cbIzeUjRv7Tbh7bG1r
BJe1rFnjNwG+4glJ/1QzMD9xX2oO8XQN2ofOfRIKq1htSk7mwwYTAg4wtnD66/hM
Sie1ny9RvJcEuNfM47SAJR/dckyQQAdWlpO0VNygHLXc7WNeydtNQIYSzArcVH6V
33jLXUXouFG375mqtcTOYwdo9Dqq19uxX2Z5yBwtb5uleka2vXunQDFN4P7T9aji
NCY8JXZGkS4ZyR6q1NGhDuIm0DCGP0agoTpC6R0h4aeKSsG2taGgTtkZKyXnucIq
fk/jrYmc/BmVM3WkOVWSDLvuM+0LecHLlkQWK8rMLfACEElC+6akIRgMX2YI2xPw
Vp33kBOhAXaOxLNGN4n/xvSjSnZBjhCvn/VOYOz+iN0536ibGeh89QY2Z8wtfXxw
RCuHUe60bPA1b3MTfZzMLhuTwdVaRgKM56no1wTKJTzajvoImcyLSjkAncT6ZUue
mGWVbsBP9tb2MFzXP+qANhUhnd2FNnZpKVEx0pSl59vmmQAX08E/hRBYvPeEN827
PLRhQpAG5UFnX+1WD8NfW+GGTHdmhkLGOoZqC+4cA0oFmjXoFdqL/ajPcissE/CW
I2TpKh/7KpqCF4yi/c09J1EBeyHRbDPMlGaWNHCBhiXojYO8qbsyiIYwoMk7gP5w
1hlC+cKEP+zjUKC5wvRfNH7X2AUoPWiH+Rxmqrna0rq+0LCQwTRJ76P0tBcV70Za
UvqSq096oiCjpP1guV2LN0SW0EgYcU+TI5QCntVY6TZZmOxnisp3zja+ziJchwt8
3sfj7SANAEc6h2W2WZ71Jg8WTsVqtet3YNLp8WLHMXhKYwqmQoE/l5kyBxAlMOaD
aewY2YUww5eYPv0qUWR9ZUsiOvTiqI5BS+0bKhlZK8kZPaG3TUwIc8cGZD9koK7b
8phMUuLGixpcCv+h3wbMvB4dS3xCVSYIhAZYzSBhkVwe8BA4PhSDyCzo1DhyiL99
xbkgVSBuqg9Nj9tvCun/F9W0JbArB9rKN2rZ00PL+FqKrWIfcKF8tRZm2owFWWDH
ELfGRtQvDi0mwkfnThxrdoNNg89LWg5XtQ95EO1wNMRCVrzqak2FvIlRgdGY0IsO
hBseHMSWS4DM/URqKPsn/PtRl/+qzJ6yy2OgPKv1NHyEVBrv1VEqF+YOxCaxyoYb
m8+IoeJyFoccIMtUg5/qZFhT5IX19BSAkMVNG28vlNAhr9Jr0JBm/ijThK9G1ykA
ujkelQ0/LD8ENB4rDBXPT3BQQeZNjYYG0kYbcM7nLfn0UAfylCGl8oY1btVeL1is
kdngYrwiDA+Oc7ziHOsUGfU3fScE9MZfKAB6Req43r7aOF88LRtEGlDpnMDIaZE1
zaAcvO1ftBSiUBZpx88gJm7vWrv0JvT+U1B046gGbE1B8jW/8j4FP6yUuvE4wzz9
8zWDxMvEXGyodvSFWV1qXk5xcL8YNAS3ErhvhU4M3Dcq0EGc43GWLyT4o0qlGA5Y
p0a77jg9wRWNGGXLm8BXeAvZ+GcHrxbyRdxGqoB2m18JTUxgl8EBAXIFHvQAjvgE
ijDf6rbxn/eKurn+caU72bpEivlxIlxiBxPBv2lOKky0MmsSJPdv11l0QIbdnl2M
T4UQNCYJfgSLxa3I+ZcdGQH2uFisn6IQRV7vJhVkHkZDZDK5PCfRbfqIQso3GzUQ
fqnda2TakBgQZo0nsKliqkElb1hG8eXWWuvO2BglEVGPm4YUiIfMQTnQ0MI8lgoH
zoXfE2qT6mRWVtluDRXraxho6TcMrAEGDtW8Ots9bjC9W6IGiCdKBhKOyjrm6TFq
UO90bVID3+egphYwnGi63kTR1Z2C/utX9RwTL07Z1ZSSV1H9xX1ej509t/o23YJu
sWmzMbny49KycKsIKG9Iuk4vNB7aj+UMTvzPx4od+O4fnDuw/0hrzWS3UV8djM+J
zv3J6KNJoLW+9JzELZ4+JMwQgy5WzukRfhtLW8Oc/cCzdllOSTdUuwJgtEgiGNxx
oxLefzjDOCxCo7MIxZvcAdafqMEN1quUW/yoFqFk4Q4RqZEre383zWw5wm6g+zsm
gS7cDmBS0Zx8jh+BUWIRd4iAEGhd1j+k3AX/xyZHphLzhZuJOSPS9gua9PC/7EE+
vHanAiOo32VN9RzwsAsvoodNoGadTX/j28M5yvzVzoD/W743UoaJNTyUsP85lC18
OalwMYt30SR3SFPe0TuOrSp/KM7HS1WpVHrtaA3PWASviTuyWgetaLkAHUWqhfqw
1MDIzKaZQ4114RiC23rB1zKm5FKIfT6AnK7fctTT78IYwzVWRlsRiz6fZ3Fa4ijU
FexoBijXXP6x6cDtNdvqfT3bFfGCAnH8ziqrzG0HLye5FUCdDRRdsIkcqNdCw8TU
WOfctwZrlAf32PJ180fAv/LTRGCT1ZHYCdIYt3oNhq/3+28AyBSokjR8inUFg7zB
6GSSdFGxWKbaBIvK/mIymvDgKDsrtNN9EXJ3L8GLPigM9aq/MSDBw0PcDfpxU0S0
cOQulEXur108wUVQQ5aDe0rDYsZeY9DK/7BLPlb9ILF5V49AtLrRWnL7vX3M2ijc
RII/JWSvWBM8pOKkHctmVk+67Py2jIIrZroCC71LX1WoMoxw5pft7Ako9s4nEBQq
884GyYJ/SDZwY1aZalJ7GvRZanebl0jvzOnYui/zh423t0H86qEp1YfHDtGAMYz8
YQqkpZAfyE9XTMZ7J1j7A2y4oTJLoSBqDcVHxqi0sRJSN3giBVjgTNMyBDSEdWR1
xkNDhynrNWk38YzsUiszjcYGNUlAJqm7qaWjmQst26sRsoTnyjr+5zlVqlpyMZMz
XSmhDgdEN6vBFQnuF5VXk3n5bqiUeRNs7c6eLhc3cafuM3JnkoB7jaJQKNgW1eDA
LOjJa6ItHe3s+xo2LbPdWLYaTTtnrLE/CFtf2q+NXEKLFZ6IBrYiM/4xmMmVvqMo
EMd8PCU8epQNDe1u9FnXxSktmrcUxAGLQyC3I22Orjbp5l1ZE/3yBS7TDuTM3SH6
arZNebInrYBU7cRIlLnn3vIOC5zhKEs2ixsYxi0Q/IHoQUaSOlh8Ej0YxtSsmqnY
AQUt4qH+lKZBnDrz8UeKiOc2w4DZe3tyF0Q6SVmNWXdxuz1HUc5fiWp3bnYZB3Yr
y1eFgVFguw+B2wQ8XBXBbLzQLCd9LWjDDcPOK4Qa0JGVxZWA/NiY59ONprG1mOlJ
RSqOXgagXUA+tgxFOhqRl4rLpWH0Ggz1vatBYJHDDJsH6yd/OavCnZoo2uL+rd4M
N49EP41cVJGxsUogY4b2kRTjsEyIXOUOW01gPSuxcZ4vSY2/XvWzfjEIy765jWv+
01tjs0r0Gu2UGRJ0f68b1OhWSVfaqclLFv/9dMXGuBeRRJBBxCSshMDxRHqmSJaV
ufgJojQW7RvGGjWzI2BfykChkJmD45hYKfTmkb+GJnracQHcBhL2W3CKflq1spEP
G4O+kqYv7tA69upHDq0HYRRK9pkF0n6NvgewtVFXJuqn3jCKkeEnx1i1HLzhbSH7
xIn148qS5smzO8IqWlhD5WZzb0eU0iXE6HLJXQTc7bDdpLh9c4DxEzguLdSppPVG
7ONF2afKTLw3aUC1bGChqF5IIkDe/7YDqohz+pu8LdunYVdb9WNXoTbUvrvfK5Az
dfFOetPRWylmbuUBWy463kOo0wOUq5DjLCIfUsh/Ky0WxYy1fysTRKJX140mlXHR
zXp6Im8CJJNw4ZsKS67Rua3hI6RAYjj+r1gdklE0RBZyxiF5tKLgZWfls0RvJggp
3wohyO710G2T3g7mOTxqoY/n/YLxSWRjKdeF1qg/izsBKf40SKzb5qFAw+Po6GsA
wz8aA5lLiAizmzPKPLAFWr8WWhl+xJoMo2sO4XQ9TxTlgAfcomEh40AqOKfXXH0b
JBtFyoVO5nXDZDJQGLmXaDT6qEPOO7FdpJj6DVmSqtBM7vToWlX1VglMVpAOVVMO
EVWzyORTlpqWa1XUnIl45k4DeJWFI4RoADh/l3X54EYtZMho7byv7jza9bxW70LQ
d1XH44C1pYxtSbk6ArodqGI2SK/sG/Qf7rSkboUzzyZ8Up7vdJIn07e8SSJU5EfK
FWvGKJZGy8JO/HTJcHQ/3V0DvRcay4ATgNL9tlSCFllrJkWhS7CWNS0Zl7UkwSjd
Ep04FaxvECf1lokDU94H+RbfM6PeNsi35hHDH4W8lQ8p0kmuIhaIhKVph7di6uNE
PuU4L99hY65BA9sDJAsHeDjzP2p8m/40SqHfk8qlhPhuqSjfNzFo5qa+s+cYK+HZ
x635BTCCJka1IGcfyDBimhDYqZzZ4BeXRP9k7BTmGuMRq0sws1A/APa58K7NZ4i7
z0mRhy6jlWucqsvLso8yTq7XLueY2CtS7bRxV5WWS39GeWAwQpzATNmv0VrlXbni
VC1uPWgzqGqJe6hk8hbWrS8PWrs8CsUzMReHXyzMRGozKOV7hI6T3YwI805cdZrd
K3e52MiPml1PnVQ3ph9D4kD16POdiMeU8tSsdqNkqThLUfj9jler7etpXlb6lLKB
sL0m0BzjKBXSSjG9ysJop36kPAGoDrbf7cDWcHZI7NjLeab7r38ztutwhOW/L0tm
WXpjGDybD42VdHWtabY9yCp5fzah4FJXZ0ip1I2g+dzD9h2Ttvc/e3mrUDPwMN6d
H0IRW+PHta51VZ8YTIkO+k1+Pyh01GFdnSNF26yeufPP9Al9syMRZ0lVWgJgDSje
tr1NIf3IOq+AFFUn+zfWZthED/m+oPQ68GHm0oBTqGcELXi2pPY8DXU+N73J4X5O
gvnKUzgf5bWQeoN0g4m7AiLfEhfei3SJHIFfGkFfgUDgfnqYSFkdZjBb/l9r5Y2A
557qloMRyl7iH946DAGXIsvDFGbIZ/6hICAux78Hh3HC9f9H0pr8qc4hmFfK4Ug6
vgrVpP1KZZGnj08RAf2cLLxMKiDjd9CfXB3FRPhy3lS7PJUTGoMYqDBm9DfNZtL5
0A7cBVqkVmo3NJQcQcZBW1Gdhzfpq0HOfFkxBSVuaADJuHp60qnII+nYiDJZzWcM
chERc+JRVXeZY4jtBmMXQM4n80u+lUhg18NO5l/YPzPos7AjlH6yMFQvm8MUBo4I
b1NjcPuR3ELypYIHfm1jipK1RGhTc9uZ9DWx/uic+ai1ft51yD/VFFbUEc/Tlnbj
hMiuF684z4iNY8ElE0hjWn7Pkir/X+DlbFani9APnN+nXsIP7SPLk5DW7uXrc6kV
HhrVB4ka7s4QaVrodr8DbJGJN104UO5VF32nKHwqwk76eTCNWgCAEafdFQgHRv+e
5PDG2pS6hLoFPqHERxW3PKGV1YWgwGp3Y1WJwiI0mTjFaL2PlRb+UfWyX3ADokt1
4rc16nC6lPy+TmeVvaBPgXA7XE4eSZPht0dOmaxyude7di+8fB/qVpl4m3+VHBLO
dNvLbIeoEExNyMpiHMQdzY+JNjB+mgaymi9mt6hKwsRwGjjf56u4tjVUcAqnMfPU
UhxczbrO0EFY+DdDXjI4VBayPWT/ePlgy00qYUALzCWyqvvT6rOQVO8Wr54d0EZS
JGrah/3IqnyVWtrVz8tOeK4rj3UIS7sFbuc8/oKKMhfIUIvM/k65k57Z1UeA7/4i
nS/z3emTVJGGq27drRS1yCkSmyeP0Al1qDJ/GnBrfM1n9KsXPDkCKIMUoMlux+Sm
XIczV0m69PyA9sF8KtMkf8lnJGU2RnKszryFWXUycc47z3yXr1ilG9+j/FMA0thi
4bUlrgZCAV46Fm4whLaygXy4T8j2AXiqrQXQXApIL5wIFB6nFG3ruD1rD9G6BQ67
iJHTKXaXuRQwpakzVo0jyF1rAw9+jy/8DyusWcBY19nD50LrEQSmEg8QRtkiWwZ3
110btfaLYLbV9BCU1I+2LtPUEbK4m6bHMAG4nZm7wqXZINJtWl+lKNVPA8N97V9R
0u10+hy409pu7c/nJOvyNwF/4sYfo/NiEDbLm7xRd54MznKLPds/qenVZMCKm5aG
iu8wtsV83VMZzG31AMaMJxKNRhGLEVjCLfJChlBWpZiP/F7sUTiTDGOPPyzwAxLf
mEVxWHM8iml5sWAMLTTSPGsu+fl7VHWQNoP6UuWWPZHFn3vit4Zdxz0FTwXxtNwB
qEH6D5i/bA6itioU1OdD5QjiFa2s57/jKxe/D1zhl2SIKgNd7LOR85A1jYgKCXTd
+LPIUPwc9qRdaNdYY6oQbpsf81M1SEU9Tmzs+Z0yvh/ddQY2YvYrrFRVdRfb/xAZ
luwEVW2RXDj1I3u0wWR47ftJIohpFN5z3gtlhTYL4DP23qFVZW/6ES/sKYFGtdZh
NgD1ID0UiWcl96at9r9K565CJZJebxR04ocPsNVgy3y5qZUnZ3ARsL1+Z+has40Y
kbztNyKQ2jXlhKgT9jmB9iWm4z212JBJ9ByZtzPnHCiReKKD2jIxWsrPZItPn7bc
zYKFkKF2djsZZZDbc5XEZx6209y6af3OGhZfOw9YH7HTnF0IqKbtVwK+3RachQL4
RMo5TpOsOkAa/yg0mXSp1c/fLSWtxtTmG60+PGaoIsKXHXW/gaHuKcT5GF52QW1q
B+jTHhaGxkB4OeG73bjWtZRR4u5Uv6Tfh0L1ZYfnG77wVHZtg5at2iBI9t1BidQY
OG78j7TKokNVHWTOkgXGHpeSNsF5rik1JAFN40qDV9reyRQxDk45eF5hAP5OwBj/
bqZYUSh2ME08Ao4Bs0TUcQYhwaPxW2FPE67/KDQfshDcXhrC0iZe6bxWD8yFopil
Krt5OgefBRDYfxx5XyDpMWkyNZ/efBzA4Iy3yxEFR2eGLElPHHKItd8ueFvQrLEO
4Edp1QTadCC+3YoK0pj21Vdbm2ibDm1yVfdfnhw17eQ6xMUrKrQ/6papbsUbKExv
F96jNhBUIN6DfvwOUxKxUW6jAOGzxxevfjk82+kRtRYX2lJu2hAArJ1KwGO8dkJG
RjiYmwfjw4qCrtg0Ogb9w+pFz98/r0fB4aqWq3n50hr+AS2HFytukwC1rbGgJnLm
url9KEWSywYGL4eNFFG7pIR5nfDF5tsXik3bKVxyU8aQQkcYz5AgeTQV/i4sV1dl
eIokfWFVSRfq7ek34H58zyDyLDvgaZXrY1h4fRaVwcVSaZGz0BQxW+fA6JI2jtDF
xPhepmPVOhX8kA/8u/hfRej4lv3ZF4sslNb833K6ehTeUemRrzQv8tjsenGZ8Sbv
Ig+mSsDYyyxxRnef5p01GNGe9xvYuCR/BFALvsnG4MhUl/n48KDvsQ9v6OiwoHIK
FRJvUenJvHScGVrGnWlBsMCZKrm3gh9lF0mHqSfIj0/3UOv/epyqPmQESI6NHKI1
OgtvLzhq9U176/M9sA0e/m521bnRYg8VNfK56zn82xR4b65Op/FroTf17TP15A5R
v+8Yxw6WDtOwmAlhqapLsrSKA6mm/78Bf1lwA71qutOjcv5Jt8qqtzqeiDHuncVn
3hpDxMhFS5iPH9UyhY33rQJrR1w48Phd1/IM3qxH7OVjAObLTsNmeTDLXR/+8JSC
q0tayIh3gQB3RCtJ4E5tzhsOwBvmadVfg47f0wcdKwqo95fkXBir2RZtL2dqdWo5
LvmonyZnkU5BLoKL/3JedPi4AyeR2PepG5F89zWrJeli/W/qXziPjrMRFMh8xxEW
pzUUyLU8DCi769PiG5dRZx4qtcRGgTb35Y3MbCRQxGAaMGHgX0bPLphm6oXY9/Ln
I27QIrSZkHICrBOnOkiAMXbq/GEeyuHi2P+Ewj5qSwZaCb8lzl9c/ZSNtBUBCEyu
1T56aOsw5D3816pOZflw/fVEKwtxLDUhtzUKcSOMXD2U708ESkT5X3Pt90aCrDuC
hk0WW00uz/eJQCfOkznMVJc/PlKrwHlPW0/tr5/BEobjgBsyjy90erpos9RVtS0e
BpDVn5BCiROZgUMSCeBx6RDOWZ9v48IwPgvMQKlG9j2gZgs3H80Az1TwnAkNPSiD
7NDApKiUEprOyQa5huZ+R7cyNW7Ba6eebJ3O2VPST+YdRdQLdCG1JPWk9wZ8+Hzq
m6G/8mtgGgmjhhO33w3po1kM9yfgK6REXtWZpTLOE1UADaoYh7U3JS79s0blUBQg
3oUV4Vo7UffZ2baZFRp5JnJ/TCmZwotNPUp5LhZmsUBpg23Am3kEQB/OO1Q+NJpV
65UPltZz1LHpyFNxEkMxFQgIX10boKu4YCoJQibhFhz1ofmlfFPmLHyw6awbd/Ga
lk0Xh/3iPKwLqcq5X/ydBXFNXFhbDLatWlxFR4JO/khOwX87BirYeLMKpNWd0szw
dPtHBlSqj15eWQaTIlaiC/2k6EaJApQ3muUBxuQw5+4nMca9jFa7eUU4eoLOvxo3
pLJ+YEs7lSACrn+/oejGzt0oANNYkz14Juw+7Q6Iat5/Yy45kuOp7ZQaKA3siywh
FiAobKJraxCrR99J5fH4JDdKC/KFwjMKFn0mZibbgV4PgYYG86pjxh1sxOVKHU6Y
Xo9rbme6uPy3B/8l3BDqWpRf3qC9cC/7/CUObopjcb/OnLD26lYBmNWW1LnHwV2j
9zcpVTyKdt9Ygu0SQjeett80do8sDmfgCSBGnYUOGX/ZWTLxIMu3zvBJLQBCq+B2
1fp8xMHbEQdcur7i9hO4OE9LKngv32HqEFqXyjVZr7DE7CyTajW9UhU3tzMI07A1
uTE7c9pig3t5NdTNdw+cuDBXWZmfSFXQhi2vGoi4xmCeVPFu5972HLCl0AE+JtMO
SLpPQnunxFFXPOJRhiTQ8jhr+YkoK7GOHFTVL+ZgEtKWH+9vomC9mzu9rXK6/fhg
X+VkinQcbVpHuLkc3dA0Wxi4xWBnloDfQLP6/IOez8uMAutSjxwrkj25SzkNvt1N
AyptAYOQZAG9iuf1XNNsdMXt/KleAyblsARuZ9ykqYUP7b/fowMRS81etrwzHIUq
/tDgVM8guP/NqoDWrNh7xcydl8kD/14Vn5I1zdIAzzJWxhA1StSCKSeAkfQF20lz
EhP1agx0mvSnzrtk4enx748D458o4Oc+lrVzKVgIhSQYMgLeXC/sFKtlXNrOG3Be
HgPmus2tbxMhlyW3cpac4gjPIrDLGLjOeLDuAEBLZN35pHY/ClCq1umF+DVpRRPi
8o5qUqWVeyWBqgQVkNp3+tSlHUFkOGNmG98rhgITUPzJMI+Mnl940yhikyYsU5ju
1skpm4DLBo1kdFsKUGMoI0oyIiSTqyV8azygYv3Lt7L/p0l2YNH1bhT+nca5QVzE
IlBFHYov9pjD3D0yH0G7JNmhDYik87DPTfxwkag6vK78uGHxbjCm1fXl18HGgt73
YKyhARfaMeOevCJ4LOSn6UH770CTOYUGQC/0QIH+TIw8ioSVCs56aJ4Jt1u3oCyQ
VnaFcd2+3P7matEJrB+S5S/7xTgG55hQF6zoNhmnTbdfuQ3WX5OeNUBs9Bun7IGw
/ENJu8PzVnDH/8oB/GOyHa0RjyKGEqofzbWtNta7EL5igDxKeAFLSkjrYkbc6p/Q
bC3i7DbJotOTpSDT6gLW2th6PKAJOOnkyzKJDjF/1OaHoPUVoD+RIhkyVwRswHQu
AIB4gEy0mZyi2bcs9qE2GKPaPSO+8hWeg7srFFcf8R7ExT7Zz1daMlQq0gSCVZN1
I6bGCEGDUhU+sYTWiMVVHfg0Yv/M9G6B4pi2ABzkGV5O81lHDk6SIYmpxJe6yXGz
trnApQijFV+SjyX+FJLDqAoXVVwkts5Mb4Oy9WTn8WB8Fpdjg5QcczOFAWk62vS1
ATirMqAXYsYJj038e0tuNC7p5cOkRGgKj9RdmjZ3em730QPF9ZYeCCj5xPj9eqif
Mlr0q4MTC+ATaWtyzWn13Mb2zOdkmdId2m7q0O4++IG1yWVEb9YU8QsUMhtN2ueJ
4DZJ8K/ZTdDkTi2tYTOWgxbSfor2ciG+lRAaGbWVeBb36bwrlroccS4ZTixx8mty
20AD4Q6MQYhy2zLfzeQ2h+ZPVDgIYHqjzMju3qFVESUknjT85OEL/jwiDnj0ix7O
cLXgCCVaEkpniY4A/gQfoz7WAL0d3bEOOSZTVrgk8GfMzfw5DfDUPSqT5K0k0pSp
1PFmyE5E8fnaHDfOEzAlsufpsHBlMOJrjK+65YWJSfwwSmNUAjB/i0X/0Suj5g4p
hADU1c2zUrtVyvH3PqN2QPhh/jL5ct8ZZ03I3MZMKlrYikEDw4p6oqrXq/T4FR1U
IvK73eAlqJ0LwgWE4sIBQlcEfIsiBFn2IITY08kBq+OOZuLX4ksygu+gZsIOp0Hp
VkGStUGZ0YeDonB/cdmRi/S+uEyuteP9HEfDW0HMH0rqLT/+U2xf2Js5NEb1V67v
xCuwv7Qq7cSfUkYhCYELfi07DvVapAEEnJvoUKmZOFylzywjqcobZly/jzNzt62u
LVg1LcQAJjfYJIkACtNorCNLBv1zhD1zAoVGD0qbuhiDpsJZWWleE1wDE45QDD0o
f3DyI0WziM7lZFupnd3VzVT9VCB0HQ02zmwWDjqwjBJgr/26r16Xay8wYSVYbImx
EhNas4IqMMD6dJfkeUopF96UMD62VUjKWh54hapWPHGSGaFrnU7nbD29J5TUmaB1
11tg/Yo0rLfH9nLYBLnWIdvjqYsi42U7KJ+AW58JG3VIQVzmUQkVjpjRYqmbAU7Z
njMIt4MHWbnKaWh1DH72RLwOQhxdYaJG6KnUBtf13s3rF6YcCm/FHGMVch1XgXJ1
ZZoyDIl33qSH2mYeL5XkUX0uwMR6RLsxz3hv6KLzJtSZken1vgAmPaEw3sfZ/usp
Gv0JjiiAvCSzYrEa5E1ill63QZQ7dMVWW8NO86sLIM5jtvTQttnPY+p7trAknfD2
JTgJu9+BEnD79HaYJZHC19dOcd+3YAF9eOYcNHzI+nRFb8SzXxqhFmMrkFRPOc15
0PtzyNDA6TKKCf4Vt04QbyyheefZcNuFx0NqgjY/xTfW0QBsAaglPw8xVX9NoxiN
rn+/+93GJCnBPFjydtx0d8sYweYwJHlmHmOKUiGWqMsGKh66JLwRnsgkdp/+pX/f
pqnVNT5YAVtULwEYU/C45HJUQbezd6J30rVXRZ6YTZeIO+9lP1A3kRQkuxvVHwSJ
EIqLfMjXgN3frxMOXAIiMNJWHdRtZP9nS2RVX9Ea39O15MHb/tVTIQwqqcgk4LW/
EBuAUJB82gMamLEoeTmX2ZKpirdPFT7u8B1WxwRkLvXi0p9oVmwXm4npkOvKOG8o
68RlTAxnSxw128zOKJ5NcBIrngG8NpgD19btkljDc+pmMr2rYTYOqo0Fxe2MTKov
/XGlf3iUGmw6Fthu/dVv/V5JwWUiQRqOQ1XmiRovXU29FUt0NGrifd6trK2qjm7l
c+NN5EjLeltOhsPzMFZq03JYAAHfPfJpAyg4uYjr71s9s4qsiYzZ6VTK9LdpPewF
Qy297Sath1smWccTO8nE54AOupFspLRSmTEnvmI4ztYz3EoE9mG8Pa/EcgAMbpVn
tmRsxY46RWPyvaCpv/f7DJUROWZ7ESAOSLnizHqhARMxJoDd3j0A6aZIZolOO7fP
B/j/msoxlTJBzteC4DPxrdOvKk2NZHK9KZmDs6lfpoOhZBq680SPdszAQSsv5k5Z
LIDJaqDXbihxbKY1xIfJHQGOI0pNrVgcq6EOqknBpCTUSM0Qp0pFbhsZ8Fxe8HW6
TdISyAo+1dV7RNOGYCfaczv952/8QZ6YoTcnqBvdg3aB3+JcodRu5wSvzevz5Fu+
MBObMgWuc+wvpa4QhPpBAX7pntKtj7547CutTx4xf1VNHdEDUhbfcbmm/iujNFvR
8WwSghbJYQ7M5q5yJa1ZIwWhz3/uFdVWHHHgdcSX7HO/zbcXKvr6Qs62GBEAjFkH
hYWQ+ajo6tir8FLprv+6mZUx0iqQVWzPWKvOFOI4gOnAXU5j9MPJ+vcD69taqtMA
R33nurtl7SpuSMB6sh/1mkZEbzTOOEhcqOUVGT+CL+oQVyCWNDYEyBP8ewyVVQnS
5Q5AK8Bnm5k9CThepRWFHQMpsIc0IRBScggWNZ4H5cwzdXlViSTTP8mAOWAxfga1
vhhkbQaOF5Bb29qQ8VM0wUMOnby5KJ1fqtwudyOH3WPA6stQ/cq8Mcuh+GQoXKNN
i8WhHBhx1Kap8LwpxCipTo2SxzPAhJoCSB/T5smQ71TxQf0vXQ7qx+nS1ERYigKT
2Q2ls1gb4NoTNxSkpNUupkIXvxQcayAt/mfOYSQ8L8+krAXECZKga8e44Cyol4eO
JPBXgPSbfuaj6Sd5rDJY0N6pTRPmYWqCuRgsoDjZNERVcpguFwQATgfTtHLPdQpv
+kvDfoonmlW4slIrrcgETC5cuxFFTVqAQfyq4eJhbRGBkIBoLG3EHy8V2lcs0Oye
XeQZV3LxICgJsifIxFClqWBjNTbWVLE9zNlgmoRzdkNhI3xorNOAK2nKJfdr8aLh
v+Dhx5gKZF7CF/0v9NA97gAh+5RHxe+2ezJSU5qZBc/om/jO1kQ6DtViJUvdtBXU
yX2xPnbT83iJ+Y6zuauNJKkulcSu3RmtyiSEezqt6nG9iZRVRsguVXzXQdJjFYY1
fAToOEsin7ZN3GTYMdTub1YDKKqOKrXqgQ3tsyu04ZiZ9IBRwsl4e4s6Yxe/F2xK
BrtPNiv+6ILLFzfuaih5/kxRqsJx3rFm+F3Ki5zLjIGWMN6gRMaUGBe/9aSJ6wbw
ut48nBZ48CM6ok6Unm6sKmAjrlx+svCkfHYSVhtBDNs9GtpthOy/3AKkpcY95uqp
9FM03swnzQamGMib5bG/sXwB+1bSyFa6EgizXiA9OMhLkS0Z54GEUC9KB17kzEPQ
3ssuKYIy0EEpSByIGAQc414oxcEuRbX0KqRNetjJIOUnzqIfRHL+1bjjYc7fmBVc
b9KD0tHXA+CRZa5Qb9MeC5z9MTJrJIYXZDqF5Zy8A2MI68mXGZ9CSK1PZvT+CCW8
8y7Arz/9tdQEEuYgElEcpR6txyd+qegnEpZRX3SCcT14K5uGT9TcyHLf8qrFPFlJ
V4FUf6bIfAKiXVOh0oyd+XyLlCdFAT/hTfK9tEOCVXSCHlzyOqOVbAwDS17+fhw0
dpOnONDt2Y9wMwuWvyDNwS+QGvfI/K1St9AXmaJ4KbYjcN/mppRJAT5l7d1j4nTD
1g7wNWYJ2M/81Zbg+4FpFwepwHekRm6vIK9HuFTyaEoDEmoBwKOjm2VitEktR+7j
Mz1E2+n27eTF+jeMjarkFK6KLzRo5VHMSjO3/n8O66GEMb86tFaMCoth+V6XbLEJ
pmSgYOPVFI/e8RqDoxdcXb4yWBNB3iacxJNFY6htwoAfOz44vDUAIFTqpAtfTXfW
o0MVNMe08mRBGTVkHAjElIOsLkumtaH0fm1Rk1iA+h5JAH3q9GVrPkHdey2fErdY
fIEpaY7rC3wbry6Fvyb78Q0g2jNWaPFNL+t8CpHS7tTVpioFy7HAUQqMCpNpU9P1
/B35pIuM50SNlCLarsivrkI7Y7Vjl5V/mDY319Kd6N9lB/uC8XXkfjmYFeI+wRGb
JSmo5DfKvWyH5VFoUBZzZNeHbndX30rB/2XjdREx9Yfku4Gmm/pRiWjQVpLSTpTL
AfeYccy0aBq8yB11jdhBOl7osjTSlB/qBMtV8Xop2SP6qFYbn7g86ZBcrR3R8zCD
q/orhSmXJZUcGz0vRpV1aKcbdgPafa2GRxxBCWSz0/Q91oN9M0+JaQelABebck+P
H8webIaP5tmz6gcedU88dshHDWxvEIAwiDioB+JZDkYd2xQrdu/6/joluxj192tT
P5iVhHr0/OsD+XNcN31dRDopGJYds642l1RkHrBrOqcf2YoXC1xmsi9t5huWws7M
cDCXoBHDcKsDapBm/ZODACT2RP45GQMtyBoswVfPguuUcPrQHKqebkgh9kEdvfpE
+otWM4cPAHwr1Fp8xC6DW4jxX7+j2bhe7u55DIn0v3NXMCU7o/0B3pNnLkQPsWJ1
WVpScvXdezDMCh1V5hDxO2CWCLtqECOwtYfnXfScSy/2udSuuIGTPaaNVKVak3SC
HNGXA4/VEM6UDkGXL0g7zx1lvZdRa9iLe6S1UBpHi/NzWOf46j2+689GlZrnvt6T
WK/xqMAER58Mnh2yEcon3prGpmuhMVL9TUzWDS47ZE77YBl//jnPs98LxFdjHzQK
N8SJp7NNM2fcrxociYfDj2VTTjkFZyNTVa0WUkIxiAO2rFg7pdAAVC6qbI2t8esX
bEFqQxpUAngc0zpu6QAtgcR9ONa9fAs/j9iRSIHVeiYIs135/zBTFdYiDWiSwW3r
VuwDxmYHpFcZylPrBxV5icGIzQ0lrmkpk4c7CXP1k2bv2XOCY//oBN4hmD/G5xFX
gH83yOW0F6/flDKfEeLQ11T8GQX0KGIJZkXS7aF6pKGF+b88VCiGlxcR8fXcH5lw
1YZFO5dYQhYwPgMTUDl6Y28YM2zsdu10tm6owbe+bJyO9HdoaiqA0+DmXRnpOTqa
F189rq4lMGoWtBwoSVSZUm/71XbIMNteYgAVPwR4aS5h3H3GLY8T9UHRHgo4hCsv
l6BxKe2bRy1fMKwt2wwaF593vW2UMuhwaOTB2c0wrYU33NyyOsO0IjVSkvFjjvuC
HqNchp++5J2CySbrYfmKu4tVkUrf0IsC6pWFr/a3wtgVq1HEnfGhQBW1/mTIvDf2
3ofnsvQ21cSTmWnNdJddwL3K88NugCe1iqhmt2rH8FlOe8xOLrjwG4YiucZ+Zu3p
YR0TWtXPg2pBz+B0WX+m95DFnJkAgqgehE2z52yLl5zO3eiHdCuzi5AwuUheHhKv
prEVVaPuHXYUWgr8VUwH/dMyysBN5778DxGtgrUnGqRH/avg/mm3vsjhB3jmt/uZ
7Ti8GvgoS5LTUQxRjr6HalCHzZzvjtMIQZAy2Oj+GdowCp7uSnRnYk58A41sQcKB
CfLMzcAolCSlvnZ3on8R3No4uXYA+NETy1xQZ2GDG/ZWRg1xwXvQ6f3yTZgDhj5u
I/d4pIq9vI1WatFBBjrsV9A0UKz63UlLI1DwrifINyRbmpkhsIAd+G5RvZC0Vktz
5lQIUExrjfOiQxvknSeHwFEwt5nO0436RjIQSzkgl1WLZXtScLvSkKxMpPl1zNQ2
Quxm2Mu46BG6YDfCII4LNw4Qfv1dE6+IhLslKSNKGcmZ/TcxH8aB8PZptmQvlHe+
qtfRVOi25bHyqxcijMlLLHc+BhjyIhYN7frFZKe/x5M2oy8hs/HDBgvSW0dx3yiD
wP/qHSmNSwysASThAO3q7cCOLKUHVdR8cWPXBjRPuVVeIwRh38R1StjlZrqUoqpS
Eg8ehaHleb/F+vx5pDvIs35xb0+ffdP1yjKZb+r8s0E5gj8SjeIYUG0oi1GTDIq8
xzMp8rYQl/FR4jflCFqvxiOmmm6ArPKmX2xfEF8Mhh+gaoUT/V5XnONAlg9vtscf
iD70mM+peEH3lnwcV/Qtk4qt/TIjM48+C/vZQi2DcsxRbvAPrr9GJ62D2a9FXyZ6
7DPV3PSr71GhGVwlK6oJRXcFARkfa365FJhpfoJT35I2dGEZLokkCKHB86nRCH+i
KD8PNoKcQhlWFIi/8RerJHkjRPGY7g4+7c5lCw9K+oeasnN86nHaSsxd4psT73xO
HDP4zjXF2HkxjzcGTSSo/35s7BCB3bGsz7F+l/IaNyPdLYdBI+V9lkpSkC52Cn2l
l42bSilUtzif5ILf/n7utm2r97HMtZrWoKItgvzwkzvNFasiDmF3WXIEkgW3lQKi
EBcNn8bY3BigwoODBE745oQr4XWp+3wozUSTCfYFuNhAAOVHD6I1/50wnOJM7fRu
L+mJftZh/vL1mCRgporBsh/DzYwdy/92LwUPcIkPTYCHPRZ2nGy15Y+6UpUNdh+Z
prxMNGqtN6+xIVyemp9rRjCWbC9lZTzwejTTK3m2pdqe9zhMX1X+ZW8WT2hJER/1
IStvSy4CpXMXXlZ0XWhmsFSHygHnjgt77wR2BIP7UXZAwoYfqrT93pEl7Lpn0fEw
tDqW/9RccqdkMT9HvxWj0qvDKPHT4nmFWDAUPGXXjomRZMdS4nGviUXxmmmch80t
22IzUMy8fE/4SGC14i1K4mXfBQwDzy5PKy6V5zlEMHaNRRAxkD/xOgOeSzCBZxHx
sPyScO1i2J5gE+5gmO0fsPqzU8vWxsp1ufwBfKs/YLEsej7qn7HPDbHgwCmFRCMY
JbKzNDMCByvnWOYPDsQzblustcZV57LxBiLWVyngk0H9r9Ey2zi4DALE8BuLDiwG
hahZCECP7P/P0KAIGfViRH88XgyAYIfL35OgAclehMh9Jy3EoExRE0YGAZHynq2C
k45JAeIT+RwVtzggafn2ek4PybUtg+AEwFrVPF2lKAEGhfaKvC19kAzRulaTh0yz
dRbD6medqoGdTlnTrPUW5rKXsOiFyV4ZgegBNcflWSoMaW52NeViE+mmHdfRdCfy
pdlArJ9GwJTRekYvebGGvGmkL7sHsOrj1eNfdTAOQNjAacQdL173WZiizjgWay7v
Y4nGmAZE4aQuzzhSbPVUKPtLWs5QUE+6/jmL7NxAIp4iURjLADhUmpwp21ibVISF
W3akDXmdEERiiVTZkJW8fBv5Be2nq4kVc2yuN5bKP9tJSAGM/qQkM0821Mx13aR5
01/AbnXCNVYjiPl/JToWya+CEevtpkkMHAlh6c5z4WA/lAnmto8AquJNwhTX4aZ1
WJGrPHTXEs7M3VzFRq3sy8IpJ7ugoiBIGpGfaJsrJfyjerPl1mwouWgCzbndGU1S
ZApx9QxHl+OtMVugsBLEq/unurRL2AKulIs6shPCr9YtbjxjfXqNmb2nDahNazD7
X+J1nqpz7RCq3Pl5bh8WoJlw81XHm0O8Y20lR+clr+q30UuUBk5hi7vAGbecYP8Y
yov9FbXiHbZUTrwEW+qc0dxsynUEtVinjvIXXzan3ogYVh3HU594AojQ0W/A3v6z
y/qL2lT6qbNgVC88GQj/wmGAo4EIt64V0j3i/P5qGdmOK3EBttDiVos0nQofXA1M
tAxJ40Uk1flN+1oQEhnH5I30aB+aEasdyn+IPrrmzyRNsuODnsUByJpiEgeC2BZS
hCLD2qqNSHvQsPd873Cwf7yClbQBwS1P4YdCbbvpMIMP+BDtgm3qXvHEXII+5htX
0vl6V3Tf8+FC0uy2KwxliGOTagIpUFie1Qb8rTTv4hGD5uMJZ/5OQCRwDkVKxV7M
5U4nogf83EGskBxvglD/fTaVZErCw3+qgmPIElKDOaXtGkjEHcFcmGH2vfiradxG
Ns22CXiJSHdNU1nC20EdBVtIWN3yduFviuRRMHJyzoMKhAqR0ygXcXgMinHEBNsk
6ir0kjtPMZMRRXdna+eMWyOjCD0upqSAZqnovr+Uw9kMbgTXOJ5N5j3U1DvNxH7H
CHF4768JtDa0ouiGXlCJPCv5xShm3JigsLO0BuAOVKdsErtT4PklnmwMLZOuWxyY
UETmWhVB6lFXTrhcA3owzEiqX81EjrPxPagyqMp1p5lPmmYRNuH1Jm1edr8lCd0k
oW7424dzNFk3bXmVA/DZeQJZhqMcT4eqMkbdU00AYYrciy1i3v7rqYaKXtLcKVd4
2V563l+1DT/qZtGhcOcKksFE/SR2+yOkNYTfSA4/8YCZTB0KOF4h+4bPK7k+f9ze
p/LB4ONWbwv/Snt4oE3gm252VX/3zpZwl4x1NXhkSpnI42gfbQzaEgTVBk3MxoqE
4+I7KKSWYyWjB9tOsQw3FlZXZy2Q/sWgIaGxKn3Y/XtwJhj7qEOPRpnaVks/4lpW
VuqB1GWZ5ffJ6dHgjtNQG1QXNKnuJwCXOVluDQhBDzpFhfh/Cop2aNYwzQ35tLiY
WpwnbMS0oGCFvae+UVqjgtOOJ4vUpW3F1KPAHkBz8dbLI/VT7j5sGiIwLQI98RLj
udkb/hjMywkdSfq4kRb4RqAxf3oB520hqYrGd1GvmANvGm8EGjntxfqK7oC3IanY
ryN8nQbN/GI4YJXjYvLKLDYhsdR4YFKRA0jfUNkvMQW6tRbXJwgI8HjUbfhberUO
DVicbUSAo1Tpp3Yzs86RiKpbZdqh2EioLfvLTj4P3BX4ObV6I/K1py+6BaJ5eKw5
CF2JhhVQ42uD1pEXk5MO+yFul164hbsT7BY5Iy8NRkzFYEoMq2z+nDIQA++m5Sgt
MCmVAi5XwmuoWonWOvsQlvmCzHc0mhIEKyppDzswFl30v9J4tkLpQAgybtOOM2gF
5KPcA8AIyDSSMfgUw/2RXCekwMI1eQ9G0IdU8sCoTa9YsfeY0OYMSovILTHDejYd
dN2oQHQZB+Da7qC4FTJ+0j8vRzHq4lLqnWVoNW6xOq29HMcZfyohWo899+yBbg/W
3gxDPvoOw1CK60O+ggLBZU6aYwwig33X8zjFkSl06RryRe0lVLlkz0NKmeTc83xG
YKUDMqMtTjD6So42pvHWbNKu2lTSVYLcHEWaPSUDkIAvSC33zl0/rFZYYi8jF7X4
+WXVb+ZOiL2WtJMMvvRdeL960drXINHvZBFyr2y1sVM4FcDlf17fpBNXvddx1l9f
fBsj1ERW4307o+GsNdrFa/gxP8Q66JiQSi6zv7A6aUR2hhgwjYJLXmDMYL17tVCw
AzcV9Zy77TbJg7kVmaTTLkv7+U8Xw8fv21fQiPln1E9OIVKnD/y/gbyFgfnYg3Pq
0XOaXYhQkUMcJ/Kk8pPFS2Wb4j8yTei2dflWYJEJJA0ZWtnHPq2T67io8kizCYRe
6T23u9QAdzEX2o54I3cc6Rd+fAXRcMeOYnHs2O9VJyi7tdpLA+B1ReVdoZiK7API
rNYYq2MRGJD1BkV5R8ePHXaVO+UNFuGiIdaBl/9qi1UC3856PBtnU1kByeaqNt6r
ndqCbwh+4j4sHG7I1QhLsUoB/fRoZcS7AkIb6Y6OqT/KT9LkI/0iY6mFPYf0I9i0
aOEFuCMwsWdKpTonFF0wDQ4Fv+Pjqlj0+ETNiM9M4AB5lQ5aZW3ed+lJhgBybUgJ
lmrpAUAXwq+Vn2pAd+y3KZEjurkbdpV8U3dn31c/lF+66cQW6f+kYEWgjSghw8+v
QEvw79uScdi3kOrVFTyL8ej/83fU3Cec232Ya9ytvOLcvKpna+9zJY6afb7cre3i
hnGeT017VXTKPDmEfCWM04G+Vs+eilRd37syxctYeM50OKVGNEOAcAHBniolL4+Y
z2/Vpk9qJLYQBKwwQ8dcZ4iTe0maRJXFBofWpGORrQhCHxbBAPYCfqx3xK7JWk8W
wSNwetj+C4jsbxeDaQTnslOW410Z32qzSfzlcymAWhYDic12ofpyj82rqoGdkbOX
gbovTJ9eVJzdi0qLGO4YuingS6Mvftj26yDtzps0sXv6C8mtUNjJ2qXCRatzf7qo
ggexuS2nxAnctMAobhAC8aX+NxQi4EXRkGxVKI07nt3Vfak3x+PiEB5Pv4ptUASc
mHvKn3sAmlNEQnrjB++BxN3Iss30WpFPkHowUIMAU6M3PplhM0qcFoQs9Nb/q4Na
Y+N6pOKKRKF2te8fVrlypSMsp2kYpV6dhPQp6awueejLxjeqmfrSdZjIlB1CmMBk
ZJtSsW/C+U1gPy1eBbxQbnDCxFQRNIfj7KynzCwcR/Bjjs1su7cG0R408UE2LdI1
uyqqkQlDtRQAWWm4XSA9E/Fv9nTNJ1AE1dBgT1wE+OSmMNSNRxgm7XuLTd0WN8cA
xGp4GZlGHRZdKfsQjbQaVH84k1JEZ5EGHHMdeoBqbBykl20XEk2cEQnEBI+bLLlB
qgYb3cXeNDZKncx/YNeTwTz42thS5Faq4brr2wWu1uqak9wN7Ip721HJTYTgrbqH
cj3kIlEANd86tX3VKo5ECVM5JZ50Z6UeWwXpn1BuMhNUdWiYJizp9u0POWvGDf2z
cg6DjGyvDEhStHJOWMWHFpD/fT0LifKAh8+O3c8mH30bHEtYU33KbvxwUzRpOzdC
/T0ftBNohk22ACF5xDOyL+RAoXuZ3ukqO0kgjO87bVkTbrjpB/L0Pha+C5jBngBi
CYLazYd1NdQSCKImbKlwvP3g0L6KH+7FQEi3ENFgGvu8oRbq9vHsV2JM4m5sAmbM
zolcqXkSz1wGxr77JNcCDrDo2zpDBn59fK3GFePx4SWWoLzwG8D5v7lveKozQuxZ
7Y0uhT44KHRk6lBOAlHfmrBUX97ut5D8hNGYMv2AiS2VG+cKcOPqNsTJ2toe8MTb
LedmtrFF2q6Sb9LVMNYmPWczUYn7YbZJzBMHmCoFUsBMRgoXquaoSPA+b1MeROq3
VDhcoNF51vjmkv/5XwPdnfjL4tsJ3tqeNyQp2ahYovE2/gozFdbttIwATeVsx1Y5
hsLYBWF1RXDQ9ZrS8zWylyUMjrRSSlEg9xgTBfz7+cLIugGR2BDVfEI9JREb4OYF
Jx2zKJzawyNkMVbyzJO5qV0Gay8N1lYREYC3l+s5ODBAumGRWWfOpaJ/60P+1U8A
Ca2LDUaiASPzuB3H7mD5BcM75+uGcCfXIDf2mm6lff+Jmc+LbMGcswxHZnwxtVDN
w5gNo7Z4ZcJwxAg+MRwzhZaYOaH1UnSXfqlxV3888JicjinCiEdGs+4uW+JAzSTn
+L12EZWQ0TL63FUDoGR4qxyg6FV78iI7seM+rf41nBk/aNISjdKDCwbiaRDIWc0y
dXtBmZSPIgxB55D5bEbJW5BkR1RWIxG3OlJ+dS7H5rU2zIIrYc7PUvHd2IKfDrYk
V47DfdDj2Jqd4NUtLLj5OKe7JlMZbXfSroWy2AFqZtuj/lWXb4Ydx6SZuXWB455G
iISmTbD62N0uScxP4ql6YEfYIfPC5FjUpYMK8KmwYK040CPblj3yR36sPLvBIdW0
FNnVt2YLJnxeSTL5fbO5v7QD/LZEed2Ox9iszFRRTnPxiMXN90yq4A2phE6kjd65
UugtnHckykykkuYd33kBcQTv+T8BxLMAJbIwM5JJ8q2kBsjSfK6L1G1+E7jfk9tu
H+mvDBPxOj/oYnjw1WepfZwDFONqxlLrAU2xLnxKdrPfYziMjlJGEP67MuZ+qEFX
2G2T/RWrrXqwB/i/UK9OX+WXLpaFqAb9rBTKbQTWA1uVSJpVWK1ENx3U/pF+W7Bz
PkWxdlER4KwrGBwKrelzmg7rXk1ViLzbLmxoiUaMg0pGo1dg0TZ/Qf2lmvpfqUjS
ZsgWuqtjatULGks1Mosc86z0s4hDKS7UkxrcgGjSOzjz+sl5M7UWnpK+lYDU3Ctr
NmxZ4CO7B+L9fEsYz9xFooXlL3eDGX9909ZL60Ma1dKZgfmmOeXstN9kk1MPIPsA
jQnDMZ4wg3k0liSnxWwna5MU6EGiTBejk9QS8zw7Gptt23qr5yoEYbuQ7Pcvu/fE
aBBDzlyOgxGVE99zzRXKJZzZrw+TDjsV8+/wUvBB+i0JsSRYYjCXAtYXSYteVcVf
V2x/4o2lV0viGwMji7SueyR6x0uxSS5cmtsRYdFdMhC9aZf/f1slvuiSaDmpsqxx
bc+TBt0h+mGeXG6BzmhGl9j2GzH9n8jPl2GcCPQKgV6xw9OEg0QVg+/mMo3alFD2
Js5AQQh0lsFeSBchD2ZIOJN1B1zScLV+EFF4WbnPMBAlBPBo1ri6E90XYH4Tn5tE
yPJqJie+/in+rftAklsVvleN4zubKJ3fHhfc5NwJzHntDr3CHWRwB9H4pfPOILS0
kbZT8UItvFvL5T96Voa58uzITDrClsyUMZ8BML7hZucKXzZCJ//sdUYg5h/kOqAb
JnbaBfWbAZk051vZ3cAs/7zBmwJRpIelgjKxVW7Yk29q4r0Gs19ZcPzvy+wcvYij
2kEwFCajP09xaTPj2IPxcXng8cyK3MppY0oJqjqZMcXH/ZQfjeLls93Umbxuxb9Q
wp5sQNv0SlaUPYu8w17IrKkAZtqTarUYUC9QRp9zxN4pwg6UVzQuInMn2F7zDnMC
UXv+m3C/RaQZKEq3o3KLK3vBrgaSok00EM05tUaSEOPq9+5MeSO43QlKjb7rjy4L
hGNH1s3VZr8yjo6tI6Dmmq9gpiDAnBZLIQVeOg1NBZfbfOlO6OBMuUmyVxcWv9lG
VVSuggphrQqEtlorHIaUzGPnmvQu8aS3QKKN2hDNurFvT2WdqrFD8fEU6iiRa4Ep
NU0VbAikbU6s3APx+8cI/OAzTB86FmxzbQtopbMDnZBj+Eqsa5wAg+73An4dwNNe
zpL4wsxKGp24vwZxvjcMbsXygQUJfIci9kv6tB5qMCUZLrOZ/j+7XxyG5BGjKP9/
We9T3i23F3N07HORZrqEKfBmUQxoOgRvPUB5hBUHIIPbG99Xrys6O0pyDPFgCf/g
kFKKjbrhBwJV9Mcnl03XPmYRIWXIOkvciB6c5qDq0V2QzvDN9nT7/ZU5kFLAPf2w
+0Kb9eLF5G9H6QtN5NdqyOWFltiTGy95d/n2i2XmfhNK9YUCwJPVv/o9JnfYjSeZ
M1pHS+CADAoyrmIIiFY6gkLlesnmk+Jgjt6l9miN11BElGRDF/JimxY4YT6eGOgq
h6NA/XB1CI1jGW1zIlK+F4OFWV8xSpC6OvJ4c6mlVY1kh3J3QBjibuQd4q4d0Klr
OPBg+pXoyvCLoldXdpuwl5PEYsPln/YIcfzM+xvck68OVCdgnR0rjuvD3sBrUNPs
VH8sbQGHjZw+ASIItccqaz5w7qu4XopIDxpRcato2RicPybJswooq7lkOuXSUb2+
YpLJYqsIMqr6zFrTkGUJk4whmlMYXqbgYRiloBHk/sF7i3gNmoKJ8a+eTB7IZ5sI
y5SvSxXGP7OhFZGgzBEYyRonHhJj1gp7aBlSH1Dx4vEyV3woW0Xn2ZYkjAuvV9qQ
3GFGBdMU0CdRYpJO0cjb/kfDvwdOByU4C7Yr6MrvBZUkA91twYXYyrTwZJ1EWMZF
gjIsIYaScsNs1hml0D/l5QU/zI8F4F+LQePBz6OTNMUFM/K4YbdmFZ+cnUxuAeXr
0KyAcdbHvm+Sd3incsc5TWxBNAuE0nO9E8043upDh/jSerL49InEtbHLenMw1V/7
gPgmxU78p3jfZl1we3w+ZuYNnoBww+GK3hnsasO/Unm7kHn7bxtrTo2hWY4Tg6aD
6KtFaVOL4l+qj8QIqzXDLs7e2rykBGRwFUZ+IUipMp+C1d3ds2lBEog5pnfRFH0f
ifckedSHlZr9a/ceC6zzgB94unH2x0nUUeSr1v+4NlK6gu19U7kwidmyXP6wJ1bm
xuzBsrKqhyzcTO0T4s4+H513YgBwQ/5OybJ8LdqWY0WbFewbzwut8od9ktGqt0mt
UoAALtphu3m/3Htm80eugJL83/euh7ffKLM0UUFtfEoFAU786g2M1eGbeCYOXD12
VrsVMmTIW3wuojf3ek9QPssZe7jqO8oMPQe6WsVfdKH/oZKNT08BZJtwq0d6puan
F9jbzfFbsDkHTekAX+Kbtw4GnrClLqsQ6ItG+aApHrNWK5cq24klYqaqIkCc5pIz
3SjT5nJyOCyIkoMWT+YkZXh1IwV1GhUJyL46wuuxNiyZN+9xJG6oR711sWmY2PL6
6Sn48I31iDz6iIbKRJDPFc2a5zobSnIr/v/nNn/9MAYysaNnCyTTSeOyZVzRFyT/
uAnFt3DxOodYg+atXEAEsxzEBwj/0li+TxmNnlXQWzNnilhByq69GXGmDv+0dUFW
qDPSHDW2jM3SslEM2Z255nkWPAMMjVPMdQmmnCPytPGTGE/n44glhCHuTqf6o1ZK
BvKsf5RQg1BUXQu4JiGxBo44BMneGzmb849kaj9kiKgkghxVdetK0yxXOsNrwbSC
60NmcMmpjt1BjLuQfVxCHxGutIi/rJOTUE/D0CspDRZ/FZdnYUgqELFrXk/RovEb
u21YlmRKcLTz0TQ3HauY6CO1rP119B312Vs+PW3yDcvqsgQ2Zct0+UiSqe47kAgw
27eMN7ZpV6ipXULcUDQG9HHIH7Ds9bBPkOHnBDBGeMUhnP4c6Q3wEsq9wjvh3HHr
hTwY16owpngsG5TF1Y9XeP93sqGVcekbANIpapzPivRKPMFTwTPduENUWsUA4INm
88AaAt/nEJmTTv4eyTjnRWSexNpehnEAYwfHphUNbCTc/hZNFoZ4W9WErrt4BXI9
oT+PBelOQi4a42ufiC4zeCFJYJiXX6uGn7UK//BZETPDzglPcmgBw7PTyHPiADuh
CKo3PajhTz9hxye9MuE5CSwpvnhUQRoJB2eQHgmgysw1OsVwxEc1o+yEHADYKzwn
+Ho5unn03O+nv0ZxKem7JYk2z0N/M6t0Z70US85cDYUADaElYd8eDY70xbHoIJkd
iLGP0ZPcK9bWbYuz9hQAPkFbF/+Su5C3Jc2RzdhyQlPMhO/cmJyZrPnR40/4Na6g
oy3VJYxoLwmejUBEOVeI8QsUuLN9ItRoeN+Qx9bZC0QugsWo5uMsNsbhQVrPOqH9
tV1KSAYKbnU2uV2fawpKPzwf8Jxg9c2PpgeIsYna/O+j3Mk00/q4eAJNMW2OoslF
FWix5Zuj03521V3I0oIc0YzQN+ustLmfQI4O0hORAQBRXq1eyrd95sgbakV8rv3q
aXaGpwSpd2zXh3DruVE1HSt65WRekskJHtlPuLzxB+zCTPVnvbIoyWBmKvRGYyBf
5PoAnC/16XK3c2I59HwnMsK5D5IJzrxQZ8cAssInTKGMEOiiEnYI+ioFY0W3y0sn
NNFCh4E5fSjdSnMevc69mMJuxY1jLtkHNDRgMOIUyk7w6qIy2BW/zfa+vjVxH3Lw
mGoLJlSwZoYPq9+7zDXwVFGYM3M8JyooERUfjEpTUnDVFbZ3vdnB3B7OafxhQuWl
g54oREj4hPTE3XyWT4rYeAL2qbEbao5PhyG5xftMqb+JISzBfB5vuUpu9RNQveU0
ymCfzxg/Sm7AetFKHMF5CgbxwOpM7dhhOyIOqeL5FcSl21jKrnO1gDTVSqediEW7
oeSXIpP+ruyykehRndqrvaL50qUeIoYAniee/nuq4Ir0Awiwoswi+/D/poC0uxC7
UALhrahgBBjfXlduSqsk7RrjR7r+9EwYklWLQuII431/c8DVyaRJm0dq9vux9jhV
k3QBphd2FcCxFhhY2UkazexiNPUY24ALzH4wXDHqo7deU7LCpMsvFT0YG07/KPIJ
3GUJI3dNTFOar9s7qSye86aTbLzlnvBzkQIXJ13NtuU8wgIoHRoPX8v4GgD4m6/1
D8jGdOci5B9v/FldVk8EcvyT28NXmZXzoc4cvE+ieuG2svCx7fEEjoa2JJIwP0BR
OLiBWiBhveipctxWek9IKeFAt1m86eA2Hfnx/pA1XEeebc6VTOIq0Is6M376c29w
Kuefv1hjRpC/c2ghpX59lhsBryYyw7D5zOq6n44kP+2fcdMMJgeSCy4jz7ka1fYR
2sG0e8IWbWAHJYnRW8eUUV/5uCFK/YXIraIlYAQwSIb+rvPt+88a8m42G/xP1yAN
dEenPSfMDprcdIAGUA+gk8/tXRmHb9HjW3A/N7bfKT7BIMwS/WyN2uZf73i27AX+
h/YLpJ0lWNyGMQtdf+bfiVit5sv2Gbpbr+zFVgiW82iXA8EQeOd81HAgvtkFCWye
twBCnST+JqsKl3RYLDAAsQcgLEiYWOYebR01Lh0J6PQiIM1HbdesQKIFInZk0wc+
2T9j3Cns4M+qFAJjKvdD9A8A8q8DkdDwnsC1dLB+fOKuXM1Oa9lnY+avBkN9vV+1
Zuq6g1GoWlFRSwC88GsMjtXa4KPSeGpBoJ4cMyx/XDwI6ko19csJBVLp9fl4gWxP
kWncGyT9b2JBXEIXVG7uGONotM6+ZhCT+uleD/HC7EZfR8NPIjpvkQI7NavQdM9k
stRkfOpntEuWt+FGBmwcDZ9aNssrlb3fiRGOpQbAgpTVOxjyVXHxz51cwjAhDdZm
523MCeS8UK8nh4s5ZHxzRibdEOrsYHSn6GWdd6QEMcLECSFi0+5UF60uNwvqs6Nl
N+T8qc3ynky7gnybKSsALXAf5w9Rh22q+RdYqdbj4z37TqmFUgDloOx+ftsXIVVO
tuw3sjzY81HKWOjlYedDtaYHNFXhh2asuFjoU6y3ubNam0GAF3gzn2gMk2/3ML78
1u9lmpTdy6hjm+r3Yq0fPEeT9grs6bQPDsTcyjw52+b8WE3hYbJ32kC6/N0n/PUP
6DV47ABUvKK1ggPuGEbrqvcieguhGfmCsEt5RftnTPlCmZnj9paYau0ervGMMSTp
kOfsggIPL5WjFL0CQ9Oi9qK41mawLxlTidZNZPMrNnFshCkGdWQuoEnwpCwAxu3f
XnFgoneVhgSuxFVjeCSPw4PLnBhiP95d0N57AKfOfMHQrw3eF3YPAqghSQ0YfQkD
N23jj7X91uI29kFNy1uKBVmPVevLJMSH5zDoydzfsbIOcRh2J04s6BXGsojO4LK1
8JjDtMpe4wW5XDzImfHRpLDLjHxur9PFzWHze8SuroyHxXNp6n93TDJtLk90CSIY
MU9e/h9Uf1CACruON+5Fy92MM7HrESyRAmCOL8ORNIFH8gRtU4fugsfmNJTt9+qc
h6gmU/lMvnhBoQkueJrNXZgBI8DNjGTNfqfQQpjpR+CDBhfclhKIgYbgASPy24Cr
T0Zj9mhlDYKPBsWw2pABP9/31zKOBrTWhJIwbCXjY1zwhJ9kDfa3/ysVGKS4Ws8z
h9kvcjvk20m7Az27eYil8TQVdeToXMRYqa1AT84VtIgoxWoeWd1+zjqykCNYM8tT
ijnTCIEBq63qDEXdKiwbnhf+UYEz5KCRCm1BbVt8dITXF9ZS2cGz6rd1IdwraoIZ
jNJq7M6xnTy78QbNTeoOGwSMMuXpOEpBPDMyQjXJFRqVZixJkjKsbV8X5SVFt1s9
NUaa4ql6gFynmoVZskw7kh51rJtSqTIeXVroSqQQpkA/oUkL6svbfuB7ggXYp8nD
WO0ZvWAIpazKr66+qApPqP4RI+wSDtRWFi7ShsFoKw7HxYD7kbKZpEqD3A3Bst4T
6uYxdi3zAn4itW5xDw/kzOoXscBbc46qgjNXcJ8z+I8S20ZY9f3vc3vQZo8WImr7
PC9BcqdmNhpB5xlPt0cBxFyL/WdBi6t3rsTTsZrWm1oESQ7v2jpqi3Yg3m/WzaDB
Let7FKqx82kCZn6w66bZVsVg3lY0O/n591OxZvPTmKPUSfm0+QjfePXi04ewSonl
wffpf/SjPahxg+6NylxJ2e+xVcU2nt1Gp+zvBgFfWxskrzdgDYr6ll8KYrKYb5qM
+DBpR9ODz+fDVKXUstn9WF2QKxMOGBSFP+qiKuriAq/ZRSOrkE0vF5JzzvZ+lSLV
1PPEB95hRJmaPjehQEx1bazUssyau7wYx2/VAwYzM7nzgaiO6Yb2oivdwnvyhGCM
G6O1UefoP2FJjPHK6oOTjS5i08+lkiIN2eUa4zRRvVGIKxN36yL+hxDpxBdtBCbV
Vczt3bTd0OBliKh+LPKCsj6GrXwCbv3eHRGLrh59USuvZ0K8+c0QfYmsC4IZWZ1g
HOjl6BOH30apYAQ/2EZ79xQKXqaziYQQF7RIhZftnyRDDoRCCRC/okJlrZi0o2RP
EI6tERVqzWsVc/s57TW5t36Dj9NWgNl63f/oIPK/0w1YNVa7bYDtr53M4f/FKtlp
yuN2uJUhDoAmy1wwsltJcffrcpOpq8j3Os4dNBckTbL0D9NLv1laHfLXlI7drB7s
KCctXbtrUVhSwjHrTuuy7HCcT+Jxe/O7+Xze8ur2t2WsWaeLFLz1X84ldoodALll
xrhs++6Qyu51naiL94dWzGzTs7r3K61v0cGIYZ3iSMCYAHmG/frQX2dpRuS/w8a7
Pq29HAZmnmD9v+c9Bx03ARK7Jeu1Xlxn3ydK31/81txuoNMCni1iWKCLdLljYO2c
6erQfs36E50QmQBP+0vFK4SBCBRG/eLfjOqRy/XyGCAfJXaqt83IPgFry0h+cA2M
JReVhi3nMv4PmsTEuJHT49knUC06AllYCQqbZahFmyGtZIEIb2HbW4twTqdgGDyj
eRqhbViBNbJRdWfysvbX5I7kYF2foBN9rMPMsCMBE1xUNc/Az8vpVyG28uOlst1K
wz7dwIQwwf051MwKDLHbWCTyc56Pj6F7qFuHXKpx+pKFfIqiRkoOK71ysWeeaaRv
U7FyQ/W+YHw9u+21FLjQzUMcFWL4wbBaJeCRTiDCYdeSVSYhfwXA3Jsj/7SMJUt6
L7klzO/MD70TiOlg6Gkb/gmDNHQ4WjWrdjqfUAq0x/24vLDf6OcU9gLgaZ5YdroD
1pWSY2S77ZK1NUp8VLjvjJfi1NDVO6odKNlMJn7pSrN+HHARwFF5G9KZoDDihhdw
iSAibDX9lYv+GBqxuBBvwgBRtPPS5qqHR6GNnMZxH8889g3uv4pewWjW48sTtoRX
gzJVFMniPt2N3wd9NhO4/phHpbL257xgW7C1m/uY0y4LonAVSvyTq4uxvZNDweWn
KcqekSEdhBZ51ez72Pwf/h2fsvseMVTfgJ4LKS/m/gJOZ4ZMxaXdI7wqx2sm71X2
peHFDanV04Cyu6usReLilhl+G2l+rpMsm66RGvmPd6bnNeVSwf6hK3qRrEzvUKT5
6wVecOasVLrL0cpi70PfXUaNaogLEXSv6gVIsKhUMK02CuVTynoXohZY5J1DMpJZ
0E5eY/34uL4LrLfJmWpL+Zy2uqalpw7H/eR+ypYD4lP3dbT80KYWuHrZ6S3EBYXZ
xdntfpZjGFsEQ1p2QJ4pQYB/o2otVWsDcEb7ibUL3rEdvK7+/bGAiGu+LhsKKIot
kZbSL/eJge5autBocxSOdLtmZfdAv21jIzuDDrKFOs+KtbEjPJV1UvxDxamnyAty
10iKkiT3XIQe7uvsGwXslhfJm45NdVGtJXfUmwwEWLkv7dc2pxq2z56JvLHnM3+C
GQrUXzeR1NLUuXoIzWLazGKPkwty86r2Km3BUPyNr7jH8GW4Kl82EINaY+ZGeRSy
oXssPNK1SLS+1J3Zgm6LiVNyk2UfFtZBVuRWz9PuVJvDpGRfHevdeWtIQjqXR4+5
u9+juWMqreiBMO8POdGERkJYWvYMVNDMA9fc/NowLSDnojwvRTsLNu+F391HmC0x
Q9LuJjD2wf92TzwDvbG9D28NGQGqQf7yWUXeQmjd7nT3NJtkZblVCitn7qoc/VNh
n06oF+pYm8/2p8WMD9wtQDuuhJxrWJgJN9/IGoc3DygeOYsrkKbPJkQNJx2tKsz2
Nn+aqfLK5mYTS19w73QxEObxn2GpDIMk3UtPW4lROBohhsWWK5V41+9ElyVzNRdr
9XRkLCgZTnAks6EznJf3sjdOGxUBEvuARBEmPNggaX2GJ/L/angtgDbg/o9B/3Nc
6y5Tz8U5EOzSLYF40cHFnSN3pmn4KpXAdJGBMCqynAreqnldRzBsrwOcacYhqr8F
BQunvlS5m+y/k3zvGl25ezOJdHhxdtxyluN0XL95FQfrk8T4l/2nylStNPLDtCRv
tMGMUmGHk3inBzet4tsGUOp7hloGSpdmDNrvMU9PLb3t4n+ZX8jqB5CApgNHZf0J
Cyuwrkii8xdrKPInZyf9ezVwnxBUQCEf/LaZd99WRu52He4H9TUGHRG/gqm1exL2
HoYCC22o0mv5XR7nmcoc1jZMaAtolIiDcUnrzUbIN4Cn7/39HeId1BPhU1V3nlIU
HqKNyQbDsjewsIHLYwHx6MyokUs8GTdBWqbV3D86hTI3XHvWeaS8ef1Llf/Vdjda
Blp29/C+AGUo1xoA7zhbDCPigcE6TyPThMdWk7RV4/Cn+6EBSVFzfAHEsSYAn6pc
cLI7ed/mfWBFWutLs/hpqq8Xy94+DODd1G4NXjnAtKlqZHWLIzsSYbA/r0sZe0by
ri+wtTpCTNkQaLJeuUG6VQ+8JOuuU8tR68j8kVcEBZh09bUxAGCSBrnoX9f7Y1Ja
GRnEzn18UwGhpQcopNvhfN8EqzVWM8YQmIMJ5GnnxJgxO0q/s3tQCL5GP4OVG3Yo
BPG/BCTDOrf0HemkLdk7LQJd69vP5/4Y+qlWvMrpwVIF7PVezSM/uNTaqMTC9Hcz
9+qgYFaAvCq3U67LyjkDDQFPOj7T1ryDFum8d4Bgss6sLFZMQIyIPnSpy5gWFc83
RtYj5NuBMVArjOpBkqySJYQr/Hx5IVce4vTFZyFHoIJ+KsN2eVwM/1EyeCp5AIRM
t6qvH22fqIXey7O0a0D0JaTLT3ETadTq9l0Z4vwqFnJ+mvhapafkMr0uZyzC9cGz
QYrIOa8EQ3SFuoil6gkRmqXojNW8VhAqpGtCyj5/1gCWlJArFRFYRq084vL1YT1k
kwMbgsW9AGUNqHIAhT2R0w6dXI+ClbNAbVdTvezdvYmULjlMeWe6491qlE7djkeN
fLyvIks5zvJ3Wd5DotIePHyRA7hx8d+TomkU4j/zSeqTt7KMfcACYN6IUlYk6vZm
tJpLuyrkAdCaNg8+QhelJwUfnbHtyUTMlia/zxQEFRQVsJFz4BMHTCpve54RndMH
R7riGPn0lBQ7X+dfFrZiUBI/Sk2vPWFBaqBJF0DVh8dx7JgtGOC54wqTOqM6qMbc
uVsXmunZJi+sDepx0MK0PVsOaMwReYutDXsYC+8YbimfgA+SeNLO7HKn6JHGAdki
fzBPy9JYsfD9DwniaCCQNY5YosFP0dp4AnIrxN630xG/FtZK6qn+fpMpoMF7/Fl2
rr2qFM6thfK30yQH5WyotiXe8qASDY6M+rfmeqd2m2r6EthbFS+HNEkKXJcj3dxl
1Hv56IG3F+0llewvlecfUhx161FH4ijA8rD4lX5EuvdFQWhgSidXqS5SDPu3qkX7
a6A61qEZ/By9q1I8hxB5wH001CTwJ1IticDQQyac8nL79aj+XAN1o0Hls+kHAd6l
dbbhSnckJLB/FStJ5AWW2Te7b8yCJ6H6gpt9KXs9VsgI06EGFU5F4NhB8rhB/JHN
zRVUO9WeBmmEXf4ec/IkkyarDUZ1EuEfQRRj0QGJ2Jz4P35oJ4s3AzmumIJ7AwSn
1zL6ft5O1d4NmSBj/wy2rS0LFNH8Nz4x6zcBlcTfxXFz+89SMViEkDGLGX9F0VGW
foG3fTIc2ClEwxeroKsYsmb16PC/OuPo4mDQQP7ScM+BkQ60NEBvko465lRm+Gne
o7Omqxe3x/uU+QygWkr6W2GP6i9QRx/7pi41aevm7zEZTy9ImJkWgWaLUilZL3qB
WyqrB0cnakWmuObpBWa2YTNgtqiVzl8SBceMQ/9BarWigHq0VMzCxwoegs5NttVE
WvfsiKI0hXWtbO83UsUgZ4O8/IfHB7WOJ8PBDzFkyeQPVUitF1TnWK1faPP6ntju
vO3YnsJ3BX9w5Jcuov3CeS1mKn+R/oF369vHHVUpsST9JPxD0cpK74MljCrlJLz4
fqo4AlC+r1ZWLFlDkT61Y9QZQjhpkKiP90JGthoH8GkXFSoWCLCrsKEUDzZEzoQe
qmZadIS+7WjjMkLoDsw/qbi3L8ZEZlYjAukSXS854/ehPpCwlNT604AJbYBiY/nL
VCSSil5cz7vz7MJUSBODdZWKGgcsdqDQDheBVR2vSETkQsLNoNPkWaJmqI5PotIX
ttBU/RMvVISbQKkR/6e62b2kJMKHY18/zgBDOCKG0aHh5fT50M6/tGnprOxzdSBu
GUOzuliVk9qOaTqQmCo5NSypfh0dZym4n+C0bYmqX9L0ZMeqzHdvAyma5R1EqIqD
91jlDY0UHFTOIfCRjy4yckrmcUCXDY6NU5Bz+mO08gA2NQ5oXwvQJRufFD/mSsyy
KvcA0gp0hoyNni8bokolFORVhqnDeukjG4TRyy4FEDFxaJH5dFBIX9yUe/8TumEi
LUhcRB76PwfhFni4dv19Pw==

`pragma protect end_protected
