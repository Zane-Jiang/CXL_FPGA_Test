`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Wdmkp6fwv6CEL1ysRl+zulXCsw0WV8HMeFkSeE6grU+XwMR402QfJ5BmmHy4FUft
VYvqCnKUDjCASU5rqnCPyrVDo9DFASmbP1tDHCirfml3cZzYspc3uqBrQUGUrCZv
3x/qWBCFLifBEO9ZLBHPwGHIQ0iVEpzFKYwXI/L1HQU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 76960), data_block
CyxtfvieSUn/gicBkdElPAJJ/hUoDRu0c0mv6CRQPtcem8YWzFCpy0sO3wlzYn9X
rMTWypBcJtX5/MC1AQzVQ9mOK/8NDA5dJQTXkaZwbhT9q4TKB/55nfeLWeP4VWoA
m7tfqygaTR60skBFwPFaIO8FYFFeMcc/Gjym9r/ytpP2lsQDQOBGsIPG0k8bGf65
0GusnmjFrvZyHwieJMHLMrm5y+QBL8fs+MHYls8cLQDDyJzjBNo/92CnPT/5OvOZ
GHBCaEsXkvRhI1yr98d2eQbe8DZvaasvnO1QQPxDeExfr1ohzu6SYGfSUlMfpKS3
YpGCH9jnoWpmphQJYzk/Wc3FCGM53fGSZ4DRXUxxyX21ScnWpQZ4QwvKh9u17eLj
0PofkcDmQ5Yd7OHy693/STa7AWf7FWdwsJ1WB6ut/O9GB+BIJQOBmKy28Hd7k/ul
TfD1B/szy8m+GXarPlUGRPbPCmNj7KK2A3tLdKCSbesWYd8YJ+d6MPuMYPc18bs+
o3fx+bKK/MZZXet1Ed62GLyH6k1wsB8bpN3H+axSkMQuqcDsH9qtLbUERqx0aSwz
oZ65YkrAO8ZQto0myqVazE7nNRM878J3lrwYsVM+Zjx87nZFk4xOtdKvbriEbJPJ
MzAeC4m8MGnIxNMvZ4DkVZmkEQICevxgIYZji9yCaLC74mADNXD/2BItcRYhCmSl
0EFaPV4csG3gtAv3b6sGRgULU3d8hBiAX30VOmI11LhEdIasD6UI2TgSpyRaTaBn
ohFHSt99Odp0WEWgLchcZoxV/GY6Ngv+F56tCJmA05m3xjtzFWzMJAxm/Nh9swVE
psUDR+x/w0jH1ceECxWBc0wXNY9sUJrJuE1FWKQ/AhoK/GPe0P1Wbjsb88wjoAsk
7/blQAlty4hLfH+kpabl7+XzPsGJvsQrYsXNxNnsKYIuacsMgoo4tcpTmSUhazNV
2tl+TLQuRx2mHbvbB20tJhhQhPtkzfPWqRG5FjMq5H/z5kCRfuSWfFIcgZBr2jpy
WndWvK6F/35hCl8deVPsobGwd51m0Y/7N1WJedALCGabN/JCeVNgvPThnQSLhMpV
7tNVOY9h0k05smffFRwU3iI0oKE889tyTx5vhPMuX7d7pL9qwGQ+RJg+tbmyvnan
LJKkXWdCzjnYX6JecFOitQxPN6sfGFsRgGV39Qe6W2K1c3oesReFnsPuShh6Ldmq
6qTrz5+iriGkJpusLXN6pwlKBgy87zUFVfUdhINUXOa5z9wS5p2uheSpwjetk7RM
MTgTF5LwAuxZyFwga57JKZRDsWcBj42J3CTtCw2Cq+UNdmURNdGgFfNL+rQXgR8T
8+wWovNu/YiUCGw2jaoHLmjqU8cKOi5rRTpKMonPzy40BKrIr3SSPZMsytW9LQDm
IY8j+r2O6Z3KEovuf369qF7zgJVSKvEiGX+B51uY9cBGN+SpG4q3HdOgPcSwcFui
k1cE/968Hj7r1VT/1upZgCwJ1S6+rbn8EMb2jiIXYpICS6rPvglJQ0GsXC9f4jMp
iRTzhpOoIf/FAywEiVe6N3ELpltwrKCdW4xgE3ZV3FXc19/0s71qpGpje6/9Ua0R
etZm0OH/NQqpTLXR+1OSm3SWWu3kvVxv3HwqgzsTTJWqWWrV6cLtedoWz+XFR9tN
aXWuEhtEzInwfJ7WuebUAUcI8fEJ6XMAp9aiEpcYn8Y6G468ZQFc/cc3lerK+A0h
2olzPvP/zW/m/HLQdR1RqCtWLFGSKBLypFVeCgulmR+82j8Obuxfn60p1kBkodmz
7mynVmtnJv750GgoWu6vS7SJbwHxWqgyp3zSHoBaMTki4iixBkriuUtrjssdDHZq
5k70c5cRuGUv2f/dx9foh6AANmdZuQ/4iiH9G5lmOgh1LVcIfvCGKqv5LwF5o5/D
btAsBavo2Jc0SJnNZi6hr4Ryeh4b2bpnMitEWJ9B2NIt527O2HbL9RDRxHmOG5hX
od8Fl+UXFXzoSFCbAJ7GophXAU5/31T1Ycz0NaBop8nO8OMrTLyqeNTKm8iyEvmc
4J6i8GAfS2sByyo2xPWIIH8ORxoH3HWOFSz5Q2qCHInJEBMIN08X2I/26RPFguE8
IMDehQyRArEkcms9U650nxtgliyJZQb9BrDhfn3PSg7EBOGfcyojlRvHN0zG3Tvc
aP7pnS06sKAJ+PQoMnZ2KeIfBFwYzLq0hzMMmqQi86jTXwWsGFsxyhfAsxi61IxO
OO0xV7/LAoAVyOEULI7Nl7QsCcs21S322mLEcBzE2oYBlJRV37DV9XKoVbYkPAoG
njC1vpsAVGj89cI0pKdW/CPNk0M+tPUTnRCIANvljkMN+JHw86tLspQCSpcGcc1Z
j6gHX8dAXEGqZW+hrG3QfqBPuhSJqA3t3cOxCOTKwzbuCKXId94PXSXwKutURqRB
S5g4qUY9gmekkff1+93D+E5UAqk601nFN6E6xnQ4QguO0NOJ0ML8iZi37NvL5hvO
1SREZulIed/h+L+QylbBQuP1Ce04UvhL2NalFUpM47+uDA6nrNhNhgTpkqSxGu/B
+L8UZ1DgjxumXVYBT3AL+xcAA4Jh1QBKhQsEIbbD5TOfwyH3+WhhiJCym6xhPVZx
Mx1p7AslmlICJU+F5WANs05DdGVX5UEPbeGrKhchhY0M/XpypyWqhpxaDxWCbUvV
gvgx9S6dWn3S/GzNIFm07W+BIxXH1CuMM7BQ1RjX5OSvagJiWDmGRdQYtMuIW8q5
iTACzh/QhR1IhjA/AUBigG5M1FcEaTUVyQPMI0Zzr3aVQrsnIlwEohTDiCyA+bRh
v7CQkB6CMHtmL/b0pchaWnpz+XxXxVYjEX3EgvddVt/hyiscRXpihqg70q/tM9vY
YtUU6cXgPZvMnyxtK0SelnREIjkgXLeqeYObABy1SiIO1QHUyHOMBLPtca5yqMYu
jALet+F+SafVt/2iCsW3CpU2FG4fczVS568fAS6WaAMwREwvytnVGaQABWpVQlz3
bGb0NVNrt1XpAZYk6G6Z9ITmlbpImF26cx0HwGgcGGspcFmYqGu25Ym2aMYlowdu
BR54D5E/gAq9W44zEutnIwl+qcpXWwspZP2xUWZTkRvmDsOVZbq8bAPPvXzqNCRy
reUnTGKXlvHdf43drKlti0M+ib3FZHXs1cFFiMeIbC8OKdw7XCKnPD8mbfaje6ga
MDjZIln+ErIx7Se4LeHcrx3EdAcjHWMPOIFO+BaSiw+dxCmlCbrkYcL962FkYmC/
XYTpVxGv5XMTUF/zhmqFawjkje3qeRuQD1/VZojUcIkoaY5pRY/DPGCKmMRvuy9I
Q2nqHwHurggHu1/QKue4BmEc3z75DCESJxfsQdU0YeGDZcXrEZTFxCKGbXlvUV/y
oF7D6ltvKKXJeWZPkEEYhnxW5gmdjjoBIrd6WRxrB5Oh+RY+o4X+3+FaFOvTFp08
/wi6Ihb2LrMs85LOheJqWfZtiYI1z7/4PTJWD4eJwC7/039+R1JsvljOT+pL17eo
RXgn9z9Atd94y107hYUok3dSDyPbYnnEf19BMI0TxD7R8k1c/e6f91/OzfBTeGP0
Id1hQ41O/BDlCGhMNifRdoS+KlirmQ6HKtynF7PwmSNSqHlHsYsjlawYrKuq0OIW
DNex53OeleI6I1ebd032VXMtmkWoOr7QMuhrQ5+KW2CTyFLhSPpTNSsajT62Dq5o
Sg1y7y58nokmiEW8qINC0YX86IUOkmdhKZN96ZRUxBz2mzrtloKtHpXm/VOXQvDj
UCLFdJHpBwkCqGcp/NuLGpPPF/JgNoKZg5AX83/cpza4zJ/GB1IrLn3MF3Mg/RdP
JqY1HD9jkURl0/1UxKDWlxr5LB0ziOdJPqq0PJ46ZfsEW5Ac4CH556apFwR3RWXl
OK2ZJccCbQqTYrJs1r40ak01MMjSkyhoK0zV1B/5Z9lEToveSTIF3Akz1IZdNXR5
FBOqrbIImAvhxcKY03n+6qWnr4vI8SeF+ToyZybPQWkE+RdriQhUtPgg11VyBiST
SvjQl0AtRS26w6g/XsxkG+5akaWMhLWvZ7/nGjbUgKmMVcck1Kem0xMjw7sVL8Bb
P75etcN+8+G61pRymd7avz5cvL5i73y0ePirmyuY3rab24Q5GEO+aWqnDv6wUSdB
4rzkoxm9oxRfuPpHcDuRZxd2TSNuspSHgcegGdtBS3cz+lYtT4xf+A9YNJTw+af8
YGNQSv/e3S8z9+lisIfgPzQETwodDFlbFr6YZEMs+sGCCtNBhIqfuzWGMXvADbqD
HXP67nyPQWla5ViX/BGBemJOnONeMI99jLbnW6xshDOkIs38yGtuq0KBu2agP2c/
rgUFDIyGyWKYIVqG4Wf5xZTwBOs6Iw/0qK8yxYWfTfRwwg20FHx6FNswufhg51qD
nPACvJuchYk6gXfSuG80swfYegOLdu4HrbkZ4dkDIPhBlkqyF+WPUh5JU5QkelkR
zMFcUFWxbZL1j0WU8X3phKPQi+0qazisYWxSNvR6fO3ZTezXx/uyTJ2CcEdZiTvl
vljiFOmnFGqP2llc984f/kXdPDj91otz3OTp3XyfU/qR2q3qxdlX3lYHpWgIKTuE
d2pwCwsmpyu8PJuTlyllKPTP38opNDemMaETzxfCApaWztExWqPwgUEyiccOHHao
YpWKYbUZmNHRGR1Z4+88TJY9eBnjVAzurQrguT0Khcd5PB4vz+ur/YscKz0sh5xB
z/LooSrjlgChn4FSj5JPjB/QJaoObt9w0Ii82z40kR3q08NNhF0W+o2SeIDJwRi/
YYOmK3+gfEIK1OG/MgoCyYmiZnUioiQchCuyw/KksY1j7DivkOTg//HUTzGaYYwk
mmmuAGABDuxdZWNRC2Fo40I1QLbxfNE4bV+X07jiMmBAiX7WFGsAKTYRVN77z9AV
WVz25ot+W5XtnC58f4/1rQYs+P00fa2jey04GJFeMP6BA1VfCMu5f2VtXIK+3bgG
JhsII/0/IyWaYx+a5dDWf7L9Qnm1ggxACfpLuAJ99GkyQk2lDDv6HBV7/7TsIFDF
I6brqvf7qpkLXoByKbV4iTj5vbq0G69uYexFcWGdM3PNYlb93Xb2+i0PE1p9E+xA
f+l/DZU6fW72mt0jwQqVKfx+pAo2Lh1nsm1419aYm70fVjOuCKFw+/sihDW/89yL
shbuIOYrP9g4K89rqeLOxh1zDjq/MEjWs9pk5H85ndcMpn+8k3unyAm/EABI642J
oagg1Hjcx4SXnGH4J4UCGB/KGDqH0sM4s6spAUbdpFCYgNp6Y9RZ9wi1CCjlF77l
tAwXGQ74jaOhTGzKiaxzKTHEHjvTRUGmLP0hVC7YO0PoddjY6VjdPFZtyocdA3s1
Lht6ovYaqh+N4u3XpvwXkRJRodwYG+aBPeiwZVj4CPrY+oMD6qPiaRBhpiFAqwmn
FOQ0PCYic+7KraO7mbdmVh6jyVORgHWlPcvgSNHpAATxayAS9+pSD8lpnYhGkpwb
5a8G8kyiCbY7F02pDpElmt5X3TOExLtSndSYndUM5zgPBKXYaRgNh+JOe2Vvd7GP
zvqnmh0mAJvdA/8vU1wIndgCPRbN3Qf6VRba2MtnU7QAW5VQ3VNC+dnIXQjEjnb6
hVdg+H6LM32PQP0Lgmk/J9B0eJOqwmZkioa/DJ6+HZite9OVcTciiZTHwTQaVMse
dvTTxxLPZ5Xt2Q3G+7lyBhy4czFr/vK5GqC0oVVCQBoAfhMgFSAk5IUe7bgsd2tl
Ej05cAP+2U7GITAOWIIHgDEZh1gnLrxfIB7Dgbmu4fFlwlQhTTF50HK+B64DkLJX
AKbOcwaODWZPyaTvwAjjRkfrYIHF4VeW/D+QyJFNR8IuIOZMlDyPqg9XdwcFwcj9
/ik24Mm+5iKe2dYLraaBjMbLDPXHerUf6NDML9mvA+7SF2E4ACoJsc/astinDnBF
LKDVlBecdxjQrkwAuiX1Yggx4GDF94AiNjhUu4ZSVP9wenmB5uk4BygO/Y7bwBUX
t4Pllf+OUSssQilb4ocxaPrjFFvlGjcCLvKVWwZZZw1ThhOXr8G4E9dju+LeZPwK
oxigx0a3cYOfgvVF1ahQrDGiZjFx64HbFQ/envgHVKGxv2f2uSlV9qNLpwf5dUnK
6+t8yjn9+JlUZU2nrLknonxDvHgZ4gXj2xzxxBoa8Ic961Zu3JUf8E2ndDEbVmP6
s0cZDFQDU08WpeCkDiAwlXqDUfdCVTdDTEaEzEeSFXANb6E1+pDdZj3J+uLTQviR
gFsI4LgAar+f+xPc26VBjBaWcvFkYQGTXX3iWLO4o6x9QaI02CtztwBqUEFfqzGQ
Sm0/UQRgp/MW7RHg9jfkXwCSv5bPfPrCZJxCWgyoXGPb62GOR0ifdHbhs0dGs5X6
sm5MZOMCMWqdZzy/5vUBLQQ2hy62OUYvkylK49oo2ENRGVAt0USZ48k1PZFYfLVp
4J7Tamqz1auDaxX37kBcoAv7diIkPWP2eURkK4TeKhfyQbDnoZ8qxwyg9zcOwroE
fOj8Me0/0ANITIfpfSLEcdq9pgM9jXMT0ZpfqupOG8NhxNjDGsrvw7FMw72aJhTJ
wfO+mGqr/taDNxmya9K/6G03Ufw3oDeE4nWd7L0CFNs3qAQdbXHZ+6HtpwOD1cHH
wgKiQi2ZOPKO1nhACGUmV4tlb9HG5U5UCylibVpi0yqllwCEYIvuKRhnXKwrBeiP
EDi49wWPGTSIgehTr2bWORWaDjWI/LMOYaxFBldKZ+gFxoE5ifQXk/WPl82zj+ia
YDhOjoESliuCCuyliEQj+R1obJk4DB/YmPYiOwBLEQaAApDcx/KiOoDMpl+q9Evs
mEucuLOp6c967jmMlO+6faU/T2Emk8SlOymYuy5QWlIX4tm8hev+E3k8YKHVAE79
R0OvSF2Ttxy5SoOpSL2hQ9iJZEt2JJqFhbO2G4PPn9xZWSVCIGSdm8NkJ9K0TuJb
XLXMBR5BW6cSsK5IEJN88vqRYdJBsBHwCZqCq9E5P9e3Wc6LIvdWZS91exwORvrc
dkhISFQgX6+WTZ7PyYkQX5jAS8RPUl0CbFuJIVqLlEpRqXiIzmIXVMTMHw3QJIRX
dnRbn+ZPrOfwcqgxpfANVc+2TaNbEtiT406vnRSnmFat94boDXJuCxD/R7ofu1+v
Jy3h0eTOqR19tmBkp375w/KlNG9dn54bGdBkUvotiXopkGfZFFO+365+5tVspnn8
yICrgJBY0RMztCWs731n9AgjYrshXibo/aBr4JiSoucXWC90AUwXOguXb4IwaH1Z
L+xYFvQNgDQSWOnM654qn1syu8hQEGBdw8dU6aHcKdnRQyH21t9qBTilauvYKcFD
rT4CneHmesRauy1HDRaVmiau7CmuQcx+kotunk8TMYmoALfwDh+TwUsIQqd/7201
CVZqpmUfFCwL1/PN30rnKeHiN6UaS4Hw733qavyN672uX3qe1hdq6R25Cwn7FiI7
kp/0WQWYYhFQFirhCZ6l5nA1tzElfJSf0/mCksTugjvRd/JbQTDXSmpiB1HcUFOS
KoEx0ZFJq7rf5Iu18vtp6UmIIJVG8J3sShctKKQfgs3412SLc5tzFvSxpgTBbmvn
VJ0bgcTIanxV1rclCOd1kORhcsk8hYmSAJASkVEXJeCVPf9PHUG8MPi1CxpGUOpA
Zm3WlxaAH7YziLvfkdWV3kLoZLPUrurGAi6wjZKFnAq75W5nVQyz/Y83wXOwKuoh
obA80E2MW3KQOvxWKr8rmn61DMe+FkPrQeZYJybZsIhmuHjojCDeW9C5j/mp4fmN
rZt+LM8ZclEOQloPoIlVxgV8KVCsVHpW5y7f+X/7wNMrIib6SelejrgnPaSeenxx
6DjWM0sgW96W9ZPAxz3SMn/vl7POsVN0HLredoWlD58fRifyHwqmvaQKF3ygRM2i
CsKXUpBcMjEzDQNHrwIC9SZDHlGva7NEWfXMIbq5zrjg3miRqBSSsgUHNffuS1RK
DTF2fCs1GzRChrnbUYfuZMHw8c2jFDMROnPZU8EF0VkBDCKnUS2RI5zUmWiiBkzZ
cSR4JnnlD2+4gcasd2rmB1Jlmiwb20P2a7g2xKKtdLd2uBcjh9Obp58RmrT97X61
qiJHn56VzhfnRIeFEr3LeTbnPz/igSLaHyVcQc+PnD+IHYIH9fml/ToKzd/m+gZD
Av6ydQddGZIVuVW9D0JKDDZ8zGXiNyO2Jx3fDPYmO0sKjSAGkDhIMdeEq/+TdbtM
4URKSoGpVWDTr1F8chnMqOfCq5KPHNmJ7c/imEI4pNiStLStJnIzKU998SmbyW78
NegzsWqeXSJB5Opd4oSIrmBffDYVRuppZaZwd6TDqTrNH9Z0cxNtTBMyBOVx+dG4
BKR6a54oxNSGd2YHPYK7S9J3sxf2tb07tcUlSQfrADtBN1H04LPZXpXOkCM5Lm9v
arf+TBLXAp0DVBHrrJtKNzLNkYVAkBwJ+wbbQEO5joQGdb1SSmR0OghQksNZCkP3
vjOG02zfQ4rCXx6zfLUNEdmMtW4F3ptqyIafznn7KHVgy7R8MxxO2zrapl49rdV2
dihLRjWWdAKmOaSd+NljsJVGjwcw6YiN4Xf1IXZ40ZlXQh1Jk0zTK3tUjKqJOXVn
rvLsZtKkQmsgtZQ326YSQd9HYYoNW9kZ5I/vzY4DLSyyo2N+eu0G3Em6q7cEO11U
cji8q4+t5jTistEybJau/lfFN+NdTlcFJ2yxqVxIjbTU7gzKjqFt8qVnCnaJlLmc
wmEbYxiWbcYipclekHpme+2ae8O2iQsnnK57Vc2fNVLlkz+kjgA3p0trMSXnz+Fe
e0cxI2lHQx/6chReBTqKFGYIkb+v6H4kA0d+W1Rl8gMJr7kCyCCL9lwTm9uR1Fvj
hfbxW1rSYc7Ct6NPH//ju8YyCcNSpYda9V3LzItA+wckyGsoMBK98pL4lkRnaTsk
8GkvM4jo4OBbQhxPnQ5M8Et/I52U9ud9I010oooiN4nTFh/FXbthuWZOr+H/Wtzw
apQw0fQ0MekgBDBxTyTH1xNzaUIYWjLIwmbDokH2W7ReTtUHPYS/QPEHaNp+3bgu
YRz9yrjFKcimacmGVudZiSRkjM8l2oEU4j4Va5K2dRBsZrrtKfVnIZ+01vtrL4w3
RIiamAppEW1XxglvUw25s0xRkfMqYjoJfxN/S89GXnB1UWaqzNPF01gZm3eBIkcf
5ZVMnqwQrgRnY919OY1N0PXW1FVEaFGGwBFmC/wcs5kOpAfehZqYi6/44+Wosawv
Ah9y3imEZdQ3iRmHYIeLE/l4jSz/IajlW3pHufLZU2garuz7PnGW2ColPtGXHkx5
V6s5Npw70eZDmHHVNw/95dmEHK7Thypgna7dAfd6s2QssELwOvA++jCS4HOaL6Q8
FMVvSxSaftbF7oT+JTXLlxRz5RjiQ7CPDo5w+W7pGJHsTC0eCztnSWrnjIshlNDb
A+NgKDB7up2t2zYmia39PtTFjs/R8RN2vM62zJqC8SQ6TpNHSCkAA4aXu6yAv1MI
2rpM8G4J20RaRZoRn32j5xpRpS9Ur22KsPp3Ya5RhKgSPW7Jp2DK2BbZ2kx4m8Ca
L/7KmO4kaD/LoJC4NdFr7bBcVGIP9s2V2Hw0mr7G+YH9nq+C8BFuhf71xsjidxnu
0EMvV8HexPHtcGgsl0lqHJ3+tRk74C4WUbi+3caTK+hGeWjPFQsPvvn8FR5h2LvQ
2i+j8wdDCXbKrn7RHzOej6ZHXBVghpM6p443xFFjekclPrbdDWvkZxeQM5mq4+NL
YB+WcZq/xE3dBmlSBuJr7vbpH65fOvS+sPbR4Bo1WEXBdSIlZ4QpZ2if4+WxnrH5
JCCtiB+Mo/7cnMCZMEb4VWX0VpUCO2WotHkSHvv3bRJUpYMeY8/xpkKcZ9Kh3TBT
4+1NIBmMA1yiBySahO5zJ6GP9SKpTDHG5kdnBrmBbhrtDu5CmOKESwZ1f1bhy6U3
SJdTpksV+bhYDXPRiHaNOZK+3TMkWKuR2g9aNIyLogEok2Vf5zUnllDIJuAbmTIy
wBi1EpaGNfancze9NVOE2XBLgJ0DJl2j3scJInTNZ1pqM17ZGF2KO66gnh+XLLNm
m4M39tMpn9+5Hhny/heenRG+LxJp6rjYuhnFC4d3udoYJOq+bB8/8wyznx92EqHH
WcM+r3RWg3DmxHSpxUU8d5IUSUBG6TV44bs5l1xJ1LLhQ3O2Kay6ovgohFIS2JEC
ciVPjK9eZPvRHSqIZTlvHiO8cuP4yqLquPNl4bP1TBmxTyOGYTUwTxi7XTizdFXn
k3/Hd8kQ529e5hohMVHGvwgc0WFguSyAuetwxNGMVVaJog76vpOBzX+6Ts2JaLA0
6Tu5UzwiL60KNBqSEDNmqYGgAb4PNmSfmLiQUzO+8V/iRRM04ixfjr0XkKxp8CzD
YSAvRKF4/Ag//nVaqEqOfBkRbqEImh4tNHnkCYvvjVkOL+k3y/eqq7NW/JReDuLC
RLKaSDE1p9zhSv9hLnSkl2CxhDbfSyqePb5kmofsNNWtuJmvNoB5couc7JlGQ8Ov
8BE3lwekOLiTNzHPxYm1JwdUOde+DBjSXoZ7u6Lt/o2BCy4DQfgW+wW7XGIwZvq6
UhA9e8in0riT+2ICcNEaa7XY2iEYBE8mme5Zth+SKDVu/9tFqbc+IjYt0ln6APgl
J40/D4Oteha2jj/SDvR9EZAAe6dpnZy1iKWMZM+6qQs3QWod0Tvf7kuWMLkhF8vJ
nTanCMuyinMuDfXMhUktlqhHuGtdVXLX4bBHpJAB5dWFwHfx7zFfnVckYa0EO6we
ZtEeE+NzzAFSEQdYr+1gTqetXnFRo9Ov3e3gd9b4+aPCMbk4Cd2cl5DQF30kROWp
a34Gr0WrSPbq2yxl0SDcR3BVzSeiXtlCcLl45Gv5eTU1zmOSZhrfoMzdjIeWt0KU
nM5PjkeMkwvjYQwgFNUyMbQsB1fkeJJWGyIujtBQac2XB6GUdtP3I6pZAVcdQ9UD
FwRqU29MqUxAcF8qmtR7rfHf+i2B1pxJPJ871NsLDJrZeY66+ARM5JX39T3JhLc8
4OHKKsPc96c4AfJEeGqmZjvFUN/z6aIgZCBXMZKxZPrD9nIH4HOiT9BEpwt01hvl
JwK7YX2DU5U6EK486XSaW04HrTWqYo04EuoKkXNglDDecT1+Ud2B8ifTtOYZygY7
MGJ+TJ2LfU8514TciYSi5zQJ8Ln1piVaeQeSt3bE7mMWly7yPCqWvlYTkQBEx00D
ia2knLxINEMTDQ7JuI4Uhxy6oWSCdY9gFOBTfX8s7BqyEwlITcwV9duTXALmLO86
XhhWgH+uYxAtJSmbXY5ATbaxMKEenO2um7W6V/bJehDvgiOt2vWo30JhBab2oZG5
vmRG9twO99veqCl9Mqtpl46aUnGkg/saO2mCDEy6HCSWOTGB0KcMk28A3BRAxTD/
il7+6xe+9UwNw0RXI8tFm2sChmU5aNerxOHNDzCojOc8fQEGJuhPekVLYctyLWM0
KW0f2kGHSN+v0wZL0oCa0D1UowVhW9SvUZEEaZ2bvvcszoSs01rWOr4wvomSPpn4
YEn8uUn8NYQChIqnznh0InFZ4kvtznI+dhsP3Nm/Q2D3UIvcn6lYPnmk/xy5996k
Z48gwSOTnnf95SD/AyFV8nB/A/8DN1W3Gr01LtGya8x5PIzpdvAV9mblPJJvNNsJ
e2qdGEC23es8qBj13VUdBD6TsTB/UICCJFZKnt3+DflYEodh5KLX5QIUkZxgLaGv
vbdWqFHHP4QhBGzMQORZM7VEyIGOtoDFcucBSyssENXaFtHqRTHj+pqXKOlyeAIa
H4TbLEZUJVso6OdAoKs3mZjAKDDgP2jD7q6XjL6Vl5+pQJNDk3YTfSDOiV1Fv8BG
PlXgIpvEP8xfuYLI99IgfrgL/Ctzr9uywHQVXjUTb/2ied3hTO9f4Hf5axEYm5j1
PolN2DvjAeSvCNKN1LPa6PWjw5EJRiFJ/wf1+SW4ExbuXAJCZwHQRxrKvIHCE21O
Bmtag9nzDWHd4JF76qczneOqWV5U2zocZUOSdKIKOtxGNaCY8awBNHDBxS7WKJpb
3Yjppg3c5xzAPw7zPOuJaAw35BBTzT7cytrDpurRnaf6y/Hy/jLGQz/Lk8Fe0CTO
lymLffbpk05ArEaNFKJAu29UgWfYfqlNGMqtZpLi9lO6dAW3oYx+DcBenB+tD5mA
muS9tQWm/WfJj3JP/CSqWLBU3i7CkfmoZpGkDNur5pFXlG/+1y+l1kVjAQrcQlTe
3hZNNU46crMQtf7x0h2B53mvoC+CtqpN8FhllFxYd1U/DR9Wv3oe5G9V96txoK9S
+ZcUd4fr5DKJQbi93S6iY+eBt7HQzNeb8Xl3tlhhHturR7dxgBj7rRwrpxDOryun
M/1QdUKZWHN0rsIlNLV/fqrlxFJDMY3wpHruixzYt2WAkan5po1cg6zqwQMJLn8z
exxXSWecSiw7FnnueZPNcQ01pnFXbBJnj/GKZ40NR+S4pu/g4ijBJ/yuvx3rJcPt
KYgNPMpkg7hAbQLu371KjyYXipKtZ/kV65/qzX7zEVKpeBtMB64gVsIh5K11SihW
CoEAxbTBaN5ur50/3BQKbti8RT38BcpdOzValh9cT2xz/gDxZbAsxXmkTPRY5TUb
OFKpQAmJsaCEHKONnyWGlk4QxfDkWrr80ga/ZJ8si/o4XQ+ZfhLd/iMeegb2/dMA
a4r+RTfWZrOE+xKumvDbQusOZ9oB5fuEQvGejdzcnfzfGeRPFv9yX6jU/zOAVRgZ
oD2lxMqj+tH4yl+3CDyTrij1fMalaX54thwqGo4WJRdBL4AcpY1OjiYGA+0+o/qq
jeHb2u7b8SAYciToH1cFVTJ8QtpMEEwyZ4LEATS3fzQItkqf9/Ypm/TF4I8Vn6j+
G9Us6aY4jbNG0ym2bbET5M4YnQ3VQBytjGQnzCHKl8OOMxvEF2E3NKbY/6JhGeu6
o/SKwd3vmfPY2BXsLwWwAQ8BBOcgnMLE7X0r+5dP4KhjxPq+ixp1XAnYgg0ykU/P
duS4wsBEddJM3sqbpwtLSRx8105RH1Oe57VL+Ef7b99abdW+5Qen6oHXno0dfusA
wX6RP4Graz/3Z0gmXhm6BSKP96l7nREMtouxkU6jXr02wCHM6JNH7vHqTqoSpRuf
2kAqGoKgjwQ/7m0ciI6i8hJ7Fg8AjmuKb2ATGyIve4LFnzp2lqW6hbkAGXGizXRU
Jp2OyK5Dwuj7WCXTutZOQoKedAg6bKDRj6doBJ7ZVwbjKky6zak8MO62r530B0Fb
lgK04lSCTIcQUooNdizr3pfVBqGUJo1Q0X1ihrSKbf8YD+L+/DeGMCXIDBtfaQx1
mG4wz4IGs3V9jPA5w5gj3jA2y5TW552iJr81JJnLLyyKvs8vh6t6mPTnEAYqpHqm
0tLGuxW9mv/2sc7R3mx++TlkMVOb/pAxzHB0VQp6n3g/TpalMRahiKcotHRMyvvm
vwVPXUbSh5TMY8JmLCOw5eTWhzf0diaY1qREOI2IQzX47GC2mO6ZaKn7vERUnb2a
uDDoywDk4R33+dvx0pLPgvg0FJa3y5Ff3YZ4Auwip5VH7I2aFsWIMYAqvZ3JnwHI
QVK3R3kbzrBNtLxx2op2THtLNfy8WLsUR6PePCD5+DvTqk49FkYkSnlaBAOOVS8g
3XJUJDVnnyFplBwodLcR1ArNBwZFqY+lsuOK2bgBznVXCxxk78FWCB+d3sejtnvI
S3bb9lmftf9pCSvNYseJpv2vwTgIncfn5j6CW7B+xpJaoUXkYhX0tmQDKa6JjUIy
sd428wl7kL82t4azzX6QTScVZ9oG6Z4CLGG/s6Y7qpbqBCePBc6o1eCDiE1ECa6X
YVXLt5lQU0/imnAQTC7diIOfn2GjSunKz6pdw6KsLlH/rbgNkRvbE36H2Opyr4NJ
5a1yTs1dvHFq+mXkzn/tm0bgRygiKs1P0A0jWvHpMZlqCizUcczc9qQtfIFZLja4
ouZSynVwIv5E5o60ha16XwMqXCykKrtg9N/8TNsM89lDIrbf9/PCRPfVyN9ddaqs
cemIc+GyOnXX6jFLlyTe0GvkjMvUaUCAvBoSFvMpDWjp8El4uJ5bcYGIt2QUJ1D0
i3+cTm3ndGrJoWb4GCkqyfeUYkg1/lwugf6NafPaZUIRmtY3VeriNhhL+JYEBM7C
O6qmzNUMq2h2I2orly2SRV/mc77vpi/C+TuV7xg0ecNj1lyvcYZsLLIufKGjJUlQ
fzMPSdhk7gZ8co+s/zAeeLJ+a2dNH9+tib20LEre6i4Y1yvJoa/iWMIvc4M3CcPi
cSmduvoEwXVCAIiezLii6yYxZo259Ui1ZEjUdnc/QkmGaEptvjiqtFRBHaUX2WNw
EFYSuVefrrTQjTbCRm1l5S9ALpkGiVVPwPaGlq7zlP70mzvZAgKaIqVHUyLyCQeX
0Lzpiwl9ULPda/J4V/11GCsfKYBCo+fsxCZgGdPT7wsLPmNbLYjY1hYM1IprBTYV
ZLFX1d1oQ2N9vZ8SLtuPM2BfJ66YDxv+1bbtWPFW18jiMEikoXC4UvhSt4ntgVNQ
1j6Tsq/zPZXVirgF14eazfwPn0p9ZN9MhbllSLoTtlEQAs1mcOBaYc06K/a4ti0S
HpaxDWbCO7coj6RXjpUUBMfZjRP2XUrWV++YfwY1YGS2JXzlvRb0YVjUK5V2h+me
uM0dnzDjq/95rjuWW9oJn2QYHR+Xv2YTz9JfhrL25dVd9PSoli94Ms9BPzscWFvQ
F5KxbeAsaHUsR+G9+rSIXCiPUocj1FSPym4Fh6zvA9PQI5R3PyVboWFa0LRRjJdB
7FFyJUOenZxoKVkC/r9BrN5XGVcFvg1HhLGXAuWZminUL7J9IgdDd7A3HYd5rIFJ
nf8eu1aOKLvRSVb+Z+8qDA3gSnhrp1P5w8zJB0c6boNVoulzWYZ9yrBzUbKU67bx
EU1v3MRkIn7Jii6/SO6WYyhAnyZDZUeyon9WvReQtm1dL/RCr5LNQ3alH2yNOcCp
yQlPoOSEB+jrL884lAfWvrI+eJAOqiv44XBVBAyrjoMPStYvLeIarOauOYFh/CO2
pO0E6mNstyiqbSz3Z+o024Y2JtsjSPQh4RDp9KC5hBzDQgDx/fStxzivtMZvZ779
t3ixU46DuhcjoPX7DIBRSyzrOWQjzJ3B2Jzgidcg0s2CQOfAFJmMfzbbRpnqtABt
MUJsrUHJXfcX3tqyI4nxTcfZsNOQ7ediWgX6uqTXEtaoMMwVHJ1Wwc9AN8j9LJoq
JOnKhi4jmqnXQty6F5T6Z3oarXUS4t5XEynAf5jyyEM1X+6JIADj1e4MvDAW5bLq
mIBLQL9yYJhGNGE2I9MjHdkO8CUNaMjEL75JCnVyqV7BFiVxQk/FIMc9TaRVObRr
30G6Nfv4+0kjl2vinwGC4LvlycRVi1aheYL6YnGynTHD4f48NOBFMrMYjPzRkmXE
QJHrbSM9DZPNzFGmGUH1cLnX/6oI5v2BDvANf7mjb6SXp91kTVcDiLnhpEOEBIPs
JudUjxsBTluMQy/TnAQUy5zyD/NbX0PVHMN8z74ThdFGBrjUVLNPH/gkjhE8DWn5
hu2WDeney4InIRFtmEHCVNQuLrJVNfuodBND7pTCECOra/1U7o29zWrcBmV+uUPc
0Bl9hmyh4GwRO+FN1LhLJtafUC499edcQQOvn/xVPTmlJzbjp7x/z89x/mPsCZZM
6NIj4+IJgG24fSyLrprA3vgIYn3vjbnz56okbPKPE9PSAG3dIuQNuIkOhCI5wlSz
pRhTHxZrGaQMZvfcEjLrhxhOsnyCsNe8kxoqFhiyT1pMg/n6io248HkJBMbEjWy9
jOYqBaxvCktGwpM/ySrflhklOUSmAOxS8aZWnyP0/xr9f2iFPmRuOgTkQwMKo7yO
JRiES3Z8xsAehvXsUg1A88erpYJlMnT7rs86S2lazgf1+eyYUANGyRew/ROfcKVr
Y90EgsfTe3Cl2BDIFFU/v9N6d4hnfxOY0tSPyc8cAONxqlskrQWkSR6nFKA+oawg
XUhDJHZLdG4WtVUbFfR5SRY3b8UjeGDgfGiZZUDBmI6u6AmtpCKAEFKkKNwQBJqk
n8QwcqV14PB1VTk5WYh4AbHfaxZdO7SsYoKNnNkYsF2W6mnJ5J9nlkO+jy9kiDI9
BNYvKsCO7SClCZlnBm9fblurGNXoh/NBbu76J7tOySXkjdEXi4K2P2LdtrHFgiQk
BPbHXXd4tQJ2gQG6oBG86GwjD3aEJRpEA9M+RVpiQDIOMxd8ZoIC/mI0VJ1mrRw1
gOoPcY439ccy/2kscGc5quBRK+dA9fga/DvkHy19MfcuYut/DZePu1Olwy8F6GH0
stHkXqR7GgFAy2jdIhbpoySecP14nJ7KqnS6zlxnSGBdvQr1HIjvaGqYX7PV2jWB
L0zADZzVzgR25GXy1YGHd376EMgFKaCzwI5vqEOP0Oftb1+hbR/GWBtZZowQt+r5
76BigVFT9WG6zS1gaFRIM+KrkKLeJ/ykEBOn9sC01gry5lhFbmD0WatUgKGrN4Kl
IR6ni9585pGnApOR8AifFcpy1zjApTP+7JjbAtHcpz41HgwUZIuXq+iN5tmhW+/C
8VBAXS9rXRyz6sOC65UkAGdonP7hKI/H+D6/1UPnKVaWtKpHsO4UYqTZ3JcHvmDV
z9p/Zzzy9/T83iaFgsmrg73Zh3RpKrziO/8M1iIIJgeIn2Uwrjng+ITs70imxgEm
hm3aqguHXKxVUCfBkxEXhmf1H/bT7tZsQ8eYnsesOIh2T293o83FURc9FxOgO8dy
LrNXmaWz6rkNaX6yzkSSbQXIjFtXQfN9tNCf5Yql+6EzWf7QLU+wHzsm/CTSwI64
5ZTaR8+EpeeTLhyIbHxAD8sFEI1K3jBav2R+aYky9Dp5nK7Wcfedq7GvvbUL7izu
GJw5WB6QmODmTkFXr3W5QbxblrNqwkjvi+Ps9SIO1vprtt9ea9jQiOCcdaLWHfcZ
OgttFCaUJ5vjTH09SpeEDmfl7NQk4svq3oUD6Z9wuB8yaxX+dr2lwIVcajQ71Tpy
ourdOKC8sp4OwyNDMtEI/eKTYpowwc/Lwy180IjHUDstwLBJEkKja9Ozri5Dd4he
qTCTSV1gCD+bbYEDNeMUwcBIEjfONRjkiP9fXfrtCmnUSy+J4McQZNKUlrRfy9P+
e0z616EeaVvqqJWipCc+isDpFmDUrTcOfyRH+O08/Kw1k0ZULx/bGk6w6JjVsjMW
h5+M8rtwprquFcUJjd/Puz9QCvq+Ro3MVXppIMsEQE+ZYTUvtatwb58um9+Z26Sa
oR0W0/91VRQbkolS/GYWqOiFimsPEqq2oj2cJVG58HqZiJkdHpIvOE5W/TzeHHMG
s+bHH3JPUscxb6JmeaQUDSIZdFU/kmmku6v+qFQljvqiP+/Gxjtf4KBH6f37xJG9
qZaTfEiSOWGUe+RN+gQ3l91+EdY9jmXTQtaDwxP77oQY1qQCO0Rv9jydkqsowRnV
E0ZGNSuaDiF2H/5rYpGSZlRBWSIZzMj9zasRfXwV3ZOca7nzIjepwSLhn33WIj3c
IOgXBSFJXnEgKrehYHAebQwKaFv4EQn+0jmaiWZMYtdRj9maSoTp1VB48hvvNE8V
3wtHV67FJc0TH1LxwnwmImvBuq07mdqReUIXx5yEUVKRR+HSba0fCk+kne4ZLDDZ
jOBExvaJ0RaI/YvZgJ1o515sLgiVG29DGNxImc6OG3cCthQXwwiiPNbFd6MPCeap
iUiy5dTLw3UVOkuPMwhDjueT+nbGprzxcfMij3b+/vIMBgXZ46l1TcJAbxA98VgI
H+1Tj4J/vH1Fe4qgzpJ09oXG1AZSqfpxNhOUYBSUP0SMF3MzVo1FSvjr1/tg83ec
Y6WXGncsYCR71CgiXHtB92utcRtJjPeZtN5MFyLkVXnQ8f1P7yFbHNENu6GQO2hY
whE5O5+tRfLXtpQobXLFQSOP+wJ3CsXjQl9vvF7ODsAI0Y1rTFkHpWpeKI5SW+oa
HZr94a+SOYq6qGhVDX6wL+IwJIJ+mYXj5PftEgGe7YO/AA9mOJaM9+gMoiJmAZV/
UmXwv9UfP9P/0CIWk41kYGINn2tG1GVvtUFoegcHYNBYCCjM4w40z5KPVR04sKrN
yrNMwj3exXZX9YW/nwXJ9svcGRbswdkfac8lkz7b6EKthQWGjiH8MCQzQRYqXF23
poWInghIq+S7oV30vOzc7Byid6LVQHBOdn+MyHv0xtV2ScsZsNC9+oZmGgc6uZ2d
OIlKkvvjKLiFLuHsgLSsGtTJFxGgLbe3Y1LXf0eHtAiSOEO1k2UgR4uqU7lVZDrw
B/hfkSLLbQbk3GlWVkeHTIIWv49YL2QSE+6P94Yv7NWccVNloSK5kEq9kJEnzrHj
Nvj0GilLoIcHvCsJJji38wXm1qLKciK6zF7JnDdvpy033KPn/jX95+gwbSXmugMs
0XSmy58empkn3tckCsYKOSuR7TLPUKV3bz/vXJ4tV9dT2PADN22VxdWofzJ3Fhnn
1yqKe9IUNg8ubfZzeI5w3pETKWN6+xDLd/ngLDYgeKDz4fHzkP29fi+fLn5/IHni
aZ0EsZLynncDOaGTKmSPYayKlMFgTkqoG3XGjvR6ETwdbTcMHqKN+lMAdUSAGcXR
tWVlSILlw9lk+5koYcOT76KZYd13L6sgj94z74E/7gVUtkh7ngA8Gu9cefxneXwC
NOcnwnIRAV9ALYxUEFl/ZDg4LMrDSI332FzSE2uobz64MTsCQeTqc6Y9UX6xitb6
10EdRPU5gSK8fjzOlMHXuxZNP7PT4q2pMonEvoJSZZXqNq5G0oZL0R9LFLyXCT00
S9LeVvOB+RjlAH8YeQISWWEFjGUXwYReNN8LlxwFtsmR/GoWJUtw01H+Rij4ntXf
+l1QwHxQxENoTl7Up6fRraBWhXwLf7nl8WYiJRY38L+Tv47DtLmUAIyQkac76UjV
QUqG0AhAl+I/pszI5Qa11Z52rZctLi63xKnP3iFT/t2wtPGnAoA3fwxdTIT3jh8m
FF7WmuJMGYqI8uV52zISmLvdPqlcW0HbdebUozXO59A5KGF8u4EmN/dy/26h+hcD
ptTwzf2grhKgZnYpFSiDDMCkMIGNNEY6aod1+8MND6Bv9u62y42PETl1ysGnsZK3
t3jfZisur2Z/anuxu6blD0tMnahxJNA/N85YXoixFZ1XIiWhPbw7ZnoegSPE8K7O
Eff/6bFrXLZbFEV6ABho8UF1MF3hdvII+fm6wipIF+QREjWNufVCzs1b829NhT3q
ED6U4eUb6jbB457KbbNfBisskK5qFzr0zlNOb41ZFOLxJqZdYyZQ5tBC23Owcc3y
N35o/q0lj51hBe49lpmSP3abSE4p60fYu2n8m2ricS+7eNZ3JD9imjUSxVHvWpVh
kg2kshzzBI1Ykg3KC01SpKv3M6KkNNcbr+2+cTP1SBg9KQOtnYylR5E2dMUq8pnL
fJQ0UV8Ji2PMzZzf69g3rBMTeQQGEoz2Uews3UjVnRl19ebhcDBKEfVLt9uygP4L
GsBoaAX2h93c25aQLBySlSy7wztAFaA7LKbnMb/VZau9hHwD1KX8k04kKMr5YqAG
nNLXkspc2KHOpXZmDSOpwaNAIgb1tUnJiC8GGrMDHpzekwp4S8+7T37Z4lhyKvND
WiNvxYT93aCETJhPs05YxLGWtgGETENbW4kkMOhn9bnVk9qTUe1UoQiDmsXrQjR3
HtUCsE1chpTd1xz8e4eBWwtE8lQ+o5JaGd3GSPWYi+1iCRCXZly31qN/GEExYy6F
OfoeYSsVlI5JoI2BPM8QHa3YTxqIsqJ6KjpieJIiNL4fSFfw1MpaJvn86ZSYF//g
W+oz5SdL4vcbP+7KPRPgvk4V50o+pVDuAC31yhWCaAApluYtd1CQy9+j3Tq671HL
lD5xiuEnCsYd8OpmPm6oKMc1W3dXmKNAGwgT9a1LYKZ8ccOavd4IOMCUJ4qNTLmU
7s6EBWqC5QQWJ5FsmSavshkkf5EbOd586tDWMJfZwusxGNyouz8pdcVHDbAvTTfd
ysaV14/bqmwC3XQlkMTY+yNxSLenMbNXGsV8dvW+M8yWqN47hlxXPfJxjX8JzFht
21CX3l5b3pSI/uH6H3llJzTqzQDFZasB2QXJtR1SJYCl2AbSzOQJR7sqLz2ZMmGK
Zue7GiHBslxH0u0UO1IkhliR+5oYhAHoqxHUojhOzabAdlCHfJxXhzgagwowWvM6
uAJgeHqX+Fq1w34Ti+IH00ws1sVB5GPs4g3PF0voDtBYqLeLc2lzMUCns1h2Ac2s
K3nQFi+fkD/HkPIxsHKfmTuP287H7e36Jk64X9mOFk2RkluO+O2U7luMFOqkFDnz
aADfLUJiuoFHegkZQuxR8O1ynnND97OccvyXi/b9z5J2ePO8PSCjUiY/Z5YuPqDW
ja5oFhuT6+Qn0DOYTffFs4Tq/Ut3aMdbZxA99Qj+ewAiT8HFEwZIbhh4FMR6MbYO
oyXS6RF6f0J2zPEEEIFpSrqWmr5kW//B7xePANdrfu6UYqtcVbDvCdg801vsfeyz
S8qS9O1dmJN7JoQq1nvnrQsBj/fm+LLD3KdsfQhGL4ltm82hZOiD3qT5PYfFBaD1
jT2OIkBC25XQFN2tP02czrr+P3uTKR6DYXaW8zKj9T91sFEwA67WleTVH3Opxv4p
Fk2vcutW9Zi412cXJfgnhRD0yCGkQ5jm/C3LeSP33KuVDWOZIp6wGgV7lE5XVKXD
9flIrA+1ANH5j0Fxo7M5nTeIwGY/HZSHTT14MYcF5+cAJCL+hUEq5ZIy1BOGyQDR
YkTfl+7cbpQlVvTpC3lqsWT/03d26DSWRogS1sJYKqYPkM/hP4ZL4jFGycsaQaH4
Mivu+T/wjjJwiQiL0q1zkF49JC2LBxSggjl4PvSlL/ZDWutvZlTJghQEM8Z3wHfp
6fofbeyhJYpCJImdIgffZiLIxhqZyVWlzvO6mJKL2Wr2ZuuaSoyPhaaMjdTUUbEp
V9fEN3RN7f0icFAzh0hN6d8DmmRWQacL8G8kEaty4Mg10OTvG9JVgYV26GgTYIch
9nNOnHyya+ivjyCi4gghZKam1AMhj6gkwFF8Q0bWHrDMYaDGYeWpBJ/Sz9ich48O
bo+AmYO/6yiceeInYd2Ip3LHQjb5owMtpRro4P/C96FlpzvJmSpqtJUacrzQSFGB
3a49h0WHkmIp+9By81fDSoCeutF/J6fhYXPQo5eNiHrIZ39DLyWhz5RE6T1Po6fE
pq/i6BlKo1u88YTB+yJLXR57XvgFmQcuFNp4xggMIbKRMA8NHLUSFPZ5o/Pz06Yw
Yf2k7EE0YjOhHi+O/597bCVyLxjFC8i+/mzW0oFF0jBP2/hyJl0efZEEW1KbF/wv
7mtuG6Oc7SdIkpUOb21Gln/EKg9rtXVVq/cx/MmqL34eM0MzBliHlc4iFl/8N3aq
FFYHUPCUeR1AmSjX5UeshURra6m1zkuJceNOT7+pYGpjuxGp+L+M+3r0Ihrpw6qA
lQtWg83Olg7IH4yBJBH0NSwgmDXtJefO9L1don9F0uAmV+HDNl08R4uQc4OVhxW7
2N/Y9cVosVUXEFkIb0q91aqMQ6QQCex4gjKayUVk/Au8fMUvP2g9jKz462iPx6Fm
FCI/rWBaTsGOYDl7EJyJPGa/9m1dvccBKYYmqPhaoTlG0gp7S+fis0irTV67Pf7g
JcDo4f+L6riV4PRlXdhg/qG9arxRrqXujESIEr3RxUMC/6SoH2NANyARxvjW2o1p
H24QCjhDNJXDPiMGWgRmBObxW/fm/sLdWiBRP0sa5YXTIb5u6uKsEVtFGOYC9UFJ
h6AB499PC1ZL1SOwLfFxy2q2APmPykcx4+0gUcSVKgGgBdt4Qj7hXyqwZ1HCS77M
7f1PqKA5RV1IxWnbm4GaHtWxsGFA4oGpTsqOZQsMGEsfyPPyYG/pgdUAJZ8kba+u
iU3pUIT5sKO8l/ksCpDnmOd3woxjpYFo7yQjgfawCN7ifyMN//5fRfVgC5NJCZLq
r4sWv8J3vUgjDbTvRCg2KFUdrIwtOSaq1YHmTJcXd/UCUEZB8Ns3nSqiDYffGZvA
5mGv6MAQxCmSbRKVAJ1hIQMfNGO/OSJblvfiQzFN+tgwiJmmqo4qPe46yT/C6W/X
ptQc0sprpTyDYiGBBj4V6dRJ1ASeTbpszof6N+T2xIKNt8IHyp27dD43ssonN3kT
zsjpgybwnc0POVOdwTCi6iRGosLCNUdWFsKlkme9/sUo1Li0KixqU98o8Fc0LtYf
9upFz+tyTM99PKBi/Xt/P3KUCqmQhqwxfevMU3ioyufg67Rwx0vVUTGbqwTodXTe
e/ePftqRAfV/hTFSkiLyIS7pzEOHwhk59CdgajTfJLELqBr+KxJNRs81LsEOTcHp
1cQigvvpNlp9sgzLXpG8vf1nE8ZGvvNWfxLkcUd3TRNl+aZkYbBE81A4wjfvGEU8
29AEwl38xcMintaBpRV1+c+E8N5XPNfqYT8HIwkAEczxWtWXl/Yk2OVw9nSJff9e
/glxxSArwhwEEqbMxaOA6hBaKYo2IJWMyJZYhGAF8cMbq8PT+u1S2BPYkb7N+IJu
+eY4eoa1uDwjGeFLmw+4xBNQp8FXJQTWBghNjb9RxhI5Q7lVRkntqfW6AMeS3Dx6
EpsX9ZDV20MpAoqXTXFw5OAiD1wUZumFMlhy50Ni3L7FUJAtA+cRprMdhNzr3/IV
VYWDKTz0wPxH6sgbcP4YGU1LIbBZKBNfSLbXvjHazuNKWV3yn4YfomepRx6YD+6A
ZckOtVtW1xovIEHiOqjy2b8OCDVOD0yqnJgBEnuFvMRN0Sz9jX5sx3v9NiCnuTrn
D4zAuuhMlu7mwhCgJgXSroO01bdSO+8P3UthFhXlpD/Cg2Z3qpxJFA3LC/Jkh/sX
Bsvmtt6jnfNGJf1WiLC7CNuI1HpIXeileO03EOFNP2mT58f2n32XVEEjkf5UuqFu
kpn/H9GQlbb8Ja93nbzVfujFPphwtwsM4mpYmfvFfaqaVUqkAxmIQ5/tRzNsrH4Q
X3NAUZDR5GgbbkKuHJwKk943lmjIB9ux3ncyZ9POAkhUEL6ImsI2JLXSCzZ1BLdV
p+lbfpqjaboojt0qoT2qilE/4kwvA7JochNaX6QEFZcK/NUbs3zpSeF9eZ4GMTKh
moqNK34oO+9F2I5iAbDHLTfNpixBqB0FvQt/xWSwoFhc13HTLoF0k/TQxDc6qjZW
46BQ0jmk2erVOY8npNiED+9gc9pyTIBt1GvoNPZl4Do+rimQMv3BenK64LtXfDkY
Gsz7ac70oxrzVBUHkreVVA8LirVJT8aVQVoKDRrAcgDRfbe9gqlEz19Wx2pCPc2N
x53f9pBNPmd+y8C6R1+ATqepf/9Y9HDYqROXD7PF9/JDe2voFiipD8NH6CrSJMgW
8tAfimKn70o98Sb8kjdyIAqTYgi9hYSzohtbpmrICegYQEOnDYMNL5/fJYIPT5/8
OahVI7AyrVdVI2fJh7Vbnm+jQAx5IWlH75hdgnjnpPC3xwwIXVNdA1XI5vOrdHgk
SmfV7CTV1LnMhoZm23UZV04PDIufE04ng6DNDV9haegJipBohE2PxPY5IFJd84a5
ufETLRaR4+0yJP2SlEvfHtTYgL+EwlB/Ph143CCKBVL/6itc+/fpb2tv73KRZus6
qxFiSr9tOVF2AWbya4PkSxyo8heKfqYjj9miSBmJ7XCIXs3Pq3Y6AueHxEeoibNz
ZpTA0q2ozjcetfNqGltGFSEZym1OuG+Je+NMh3NQZF0xbOa4CW9buIHg2C5Q5Z6f
jWQXFr+leKEKaV39vbz+ESJFNKLiem3Tv6IjGpROgICpKma8No108EmgtMUtUqzn
XgZQFV04EZ/qMc9UtCOGnR0O9vG806IkM5zY9mYgAPvlGW1zcz2/MNFmei5FMxCY
RSUSzMpoTjW1+GB28f/Hnr+Fs7CAzHGmrKhmNxnd8y8O+D1ThsSCa2q7UnAb0d52
JqLwBiNuur5Z8vV2k1UXLP6anmHCU2i6k71QOFB1UcRapqeF2Yn9u0TGBRewqTaD
VWpus9gvwm/760EUq/XFT7wfop9R/aSN8G2Bu4oP8ppB+Fg5uK1XGQYrC0xvsWRE
0Lx+uUQcx7qXJzFBwDtjbfaQWMJEkWTHq1xSC7YS8km0EoVWRl0QIw+Lgadzjt2n
M1uZA2sSjbxDGo/ud+hLL0fFEY5d9aa53nnC5xFURKCoNULHNCG5bWWr8T9FzpCt
Dwr81+qiOaHOW/GAWRqtAUr9HhuLGsTdJNkV1DuuxJOC7phA2ejmMdjwmpO3yuZR
vKx1PZoATRDfCapi2+nJFPyDQnvuQ0ipfkoeE/mBkROXwJC7HvfYyxuk+Lk+fh0u
6B2rT56xEni9A2J0haaQfteOdZPQg1VfVwy20rEY9bsOT3I4OxZWaRgEs1+hJpSm
0ShMxfIwj+G4Pyd5Tr0Vn5uXZldTYOxBKyqEUR2hUC2TxXMUJtEnHP2x1wGCG2C7
QBsfoRUryqNs2ty0JTmC/jcvEhxUyyDFfioDDUf9kvVji00aJYU0fxGzuFJkBkpV
r/FdUhXLc/IVZSYFMX2sFOkppk2AN/F9UY8tC+4/WF0v0iGNMvhGJTk9mWr7S1WP
rGOk4Q5sacze0xSCgIkLCj4UGNMC3XE+7M2WhTNIB3Nj+HraAOWhLCxoXfXygFEK
G/VQYPQRRFZlzEq+NYylVGWKx3z+QMpA7RW9CbrpVeI4y4WyfHsQAsoQUmQCP5tx
/zi81MU5mKpiKLCZhYi0Fd01fC0Zl9fXEJuRri3vTn2v39PcxqQ8P3Q3Ak1WaqiW
ATcGh7ez03Cjcl5A2pvrLrvPMNhJSxO8TTtN705aaOu4vgR6qGlTeKGwRcbtrEcG
FOvAfp0BruILQ+AMARGhW/HEbreHkZ8RDAxffS02Ht4yXLRHlh7/dQAaGymqeEcO
nqE7/HvzDSHnbupMvPmGvu1/6eHNNqSfhlG/1gevSMMYS0sfHc2hBH2Q9e9dJvUF
yvYr713bVRzK6qXPWVeYLjp3WhUXy1XVDTAhKjPDfVBRZf4l8mbcapXwuSg+XePY
7THzfCB6+5uGtqozHM4m+mb1ce+9lTEjW5ZsenKU8I2IQjQg/cZ3uqoltlQLJ2Ho
27hPsfYrRgxIWVvIgaYTYe1gwbJ1nLENP5LE30v0xr9xescdg+Y6l8HKSws/nW29
xyWzpDEDkdqGxR9E+n0LAVh/JvkpG5YXFBCFRcaQEdwpbAI7+Ois1sexFX00iMtO
W4/g8TWHZCB50f6bKbpSPSmZw9/2aOuHeIE8V+rXeY6dHsUR0nw8OdSrgrjO8eqI
klZB4KRVSh9pe7g6KolN8+31bC+XhsQ5eCuyh4gpeIFqa2bwLa+lC+WiqVfa75Oz
jUOIZLMjQY46a12eoFGzRAs5N3itB2sxPsGNnWB3SWhb0Pmoty70wd42Xx7bNbY9
Nfzf5UIZ1wCMuUdDHEau1mlJslZYjGniGg+DudzDIJETBeM5FWONMiZYm5/YCqBC
2u0rv8p0/pewNF2MSIpMwPHXKhNAND8RU7llzdmr9yfzm1OMYeOTj3xZyDfJm9mm
pY3qIFoBJmfNj0rUpjOlo7PxbGb+R9Rpgu1gI+L3lhsMtooHq/8iAEWoKK2GoNf8
pr42Gnzw+pmbuwGtZFyLlkmzJArzbSD7lhYaAPJXipBIf5jVa81HW0DF59v5hFxP
ITq3i6mf/sArNu+Pkr2gnIKm+bJRVqRqtuZ8sGChfpr3k8leDsRO+gXsxi9Gp/H2
FAMU244+tDKu523Dvib5NXUWPpQMVw2WJmJ/Q6j8uNOjVYczrWtvu2tk6Y1Va5jx
5UNFfbNGrNk2ccrxIpDvu4xsNr7QjtekOwvz9/SZL3ep6wyLalF1X1qR4PVIA4A1
WdnRTGIdfpWnDd0UBLimifr2v+27K1Exvlfc2gIRqqO8nN/Uv6SWUEp9j8mE+6S5
vHddXSPcKHazka3HEAbqNLp2MoJ1c4Ic/90UrFOXSXesSyBebKfYM+QE4GfoQzk0
/zcs4Kqi2Tudh3jow/uXsxOaPL3/avt+UAorfEO/4N7lNH1IbFPFyHltd2LpFj1W
VlpqRRSBV1CYzh/kDWObbHG5HYfwOlFEZTslpjBPtzN0/YsZNIJUZrurFiZ+reww
sSw21oAkhhYPG6ITL3cGk0B8v+IYRl0FVvUk9TrK9u95Q/3dRkAT2yCVr9YbFf78
Ky/BjRsXWOCioOdLCDum37aIv22ObPlNf6ytyK7P+n+R8Q1MAEIn3IA72VacDkyl
WM9l/fNRpICy2J8naPhUgYgCBDAV+i51ty44cACB+tFTaFXRWSddfNMdxjIuCESy
hkFhB6GuMMqc5aY05jx3VcGwjFFfPv82jv4irTkuAwAFBeT+0548wA5ZGpxBqFTj
BgxHfAie6eQytmnANDKhBhlYIbnbsbbCoirSgg0TlcN+AEQO2JDjmkx4NRGD7e4f
bi7RkxxynTiNQut64NvrFk+bZSSsEHepV1GB7nT4wsGarcXPHK5xH00Tq8j/Ozgg
rId0xjmN7/xd5ANl9d62lOwaqx/T+vXHFlNQ96tgrtyjUmVy6WZDFyUZ+VYzFZBG
ZIe3sSCbohiIEO1NGmnMIQH6owMv1AC0JxFoyHcWHKmYezRCVIM7YuTOk62JU+0z
8s1zJJom9tyi5rv8VZumTCIKgp5OgtxDAw0ojzeWIki9eBZIYf6iIIqAxPtt823N
qSADSVIZtQ+kgFSNQMH53PY8aBbRQilcBAs/I+YZHBUxueRlcVxdRKhDV1Rty8G0
Brw1rsKn6smBT8IdrLFVldTo/fG2Uknl6wZFNWe2niVlOvjqN6RQXYdi1k/gVk9d
SEOK7PohvxBxUxWLvW7JorZ8nZwFGtAr8HoYp835ENfMiZS4u1H5igQokL8iV4CM
BWcbaKBvIVsWRHEHnJwC/AdsIYQESyWXLWscacq3wbDFlGI14oN3emM/yOJdekgp
qb9sgn1yjS7EaPqCLdAkFpo1wRkjVPe5SbtTVkUgyjAxDSQQEkPm4gW16MHEoaou
KVl6qfgEEDMnJOIp/ecthn51v9SAbz/QRiKcZXyh7y4nT3UUd980OPum4RsegHac
zIpJCM1CadHrFiHkMC9tQGY7IM6fx/PC2tdUpR7HF6gmpNbl3pdVhOIF5UZ69owv
cumbEcnKG977GnfNSFtg1JlXCWOKbbBcqNxCcj9diaHRQjQI1bUyeJIVTxQHtQHk
CmBfI+88s3lImnQOo8v/EGp+snUBq/FQG/zcY3+/xpfPQf/nwiTp3SafFGbIkZyw
FQOVeonZvoQEHGr9+CZhwfHSFu4TqF/Jt/F3D7b3fphxFgGpIOkFuMSKJjn4alew
a9RTQsAcdIXAt2glYNaCfo8nXwyNWPBLsHStaeM0Y0D+IgOo8zY/wX0NPH60vRkW
EsXacV3RS0rPfD+7h8Yk2cUauehEfk8PhZTHBxfa+hs9VArWMB4EevdV1xbVxieG
IrSMzVVRw2s3wmJAMc8na1d2AfLkbTKLTwDEpdnK9NrAzyaqijIXxwSbrzNF0e+W
8PTQiNQffksaWmLpTqZhqFYSOFvwqcoGqkdHru+H4smQ2UucNzsYv0B7togxKTo8
Wxs4T5ZDpdvtS5OIxV3S1Kftj+tX+KQF9GYNYgq0DyXXhnslk4dj/1ZCgJByoUJK
F/LXf6bXNEUcIJOXPsqgLYGk/cbDe+2LwBjJ2rGwC99mYjGAqOSHbI+1SURBTqUi
wzh6ajawcnyGgUyAO51raNsB2wbiz1Mx1HGapqs7cXriPBsZsPbQouIQRB3EnXm3
iGLzTlCw82mf9gEoi6BhfdMNoXCuPDxeK8xzHCd6Pa5LAPDOyXzCGlPFU0Chuab5
1W4+iOmpL8/fgI0X0nGPM2Vmp1gVu27RFfWQNF6Sc/xSAlBzE+Z1WUZpW+l72yFx
emPMsRiV9blyge0EKUosYWHnUNWLaOfBS3Jny6EuKvlx1Q3p/5tNmMCxa+znZhYg
7hSDKYxtjyeGDFi78/GADO3boc0OlECFShflnRx/7kqCMWnHshAAIwSdotogkpnq
uwL8rtNY3N8R60LO545v/ZEm7Mw0xqqdanqyYN+/9Fje1DuYv/5LXkBqKbKkvjEy
cw0+nwyfF+6ZG3h+9CYYcfebsBDKA9g6t++yrgLtPwFk+juEaG6lc7zUb0shPMma
vJCM4jwTKU/Nto+UcIjqyZvptpxeVjHRFAKUVdsHQ6i3EfXdbNNXWt3mcyToeNFl
1JLG8ZvrG4gz4TZpFx0XS9ATnXGMoqAQSpeKRPWIkAyT5cm4JClVMl7EYnoOG7U+
lNAjWlHuWzfey7kp38YfhC7aUtopSYH2W1c9o0zo9GKGq5b3HjXcTqOaHSbcrWMF
msLcX0DB7QSiJ0YW0irbMJtu5Rbv10nzq4BfnxeA5mmh4nyHR1bfFSmsrJ4v6NYe
RPVUaXm/+p7uRFBmMcsCRgmDu2wfJuqJaMQOimcu6CKsKbbrcsVHGvlTzOmDhJ8p
VFEIw/HFJvFhdwm7ugtgYvFamvL/XXTyidyNW7dZmJUJPtUv3JeKh9h8krDmT1aq
xCKJYzYEv1ja8GbzTvs64ZZ3zaF9TiULO1O3AFtlyZMPmC8bAJhUrsU627xHM5WO
y3pu9tgewMdmzY9ji0/KJoRN81AgPVWKbJyyHkTEsYNwOvPzcWKjVSMZqRvO/s9U
mVH/8CJ1Z5qVgopa9nJWYIn9OjEhzVa8uVkpGHDKQC7vnC7iFRn2HS3XyS3WX9pN
LuOOzjv+J1uKHugjxu17clJ8rELnOR63bbY40tyuYKYibVlaTO0R6nIUTpggrThX
NRg1AlP+zkhy6SlGBi9HBXBDBUHSNVr8jg1PZO5NpeNrPI3rRmANP6gxLtVLuD0H
SIFA+JmIMvuVUso6YlhcIAoP3DP1edJzj4vYc7rxIygjSLVqVDLCY3gHpuYIF51b
yz3JOI9lBBVi6zgbBucC+tEsZxEk4+ifdOxW+X3p2GrLv5wBZtEYzEIZASmP4vWP
RJYPLX+oEcEpTLarTtCrIvYrTxtCW68WSmz667N90XxVzZ9CG+Splju3gtmhKF+/
21uEXBilPxwavMPGVoQpduLKJs0rJqHZHLxUMTdhQoqgWdXsGHqQyKNH5/hCAVaC
ioWfY4QXJKe/uydqgiM+E1ED+zgNDiCqRappzvMnLy9/hN7jq1my0AwEYhFegBIO
WryFOO3GJznzSDQCXk/GVoXXze2+9Jfhit13BZORub+i/WW1xcxzKd5I6jGhtLl/
UT0LemCM/O+YGE+nM9AVMkyLArsxbzXk7sgxn0FdCwFeThbxpmTgX8lpk3hWdsb0
BtSpOF3HAr9W/uMA2oCQjpuqEo2Jb5A14rHQpPEhsOTzxV3RFx77MAhxbLdx8De5
YSLWdCT17avly0aqMMSRY05trpddUFdRDW/q5IOStIH4I6GO17bHTcCd0/CK/FTa
SvuMnNIWDaBL53/B1OmfL56t/eIaZ2WWq53Mmgen76Wi69ZP+VP5lhkzccHr5cOM
wUwcGls5F16gy2oLLy2ZveFn1Y/ZzNd2FUzpGxljWS75gchVrLBr7pIybJyThSzL
Vrz3TuCaLOCbmG68VyeMoO3VtDrqfvexfykaBfcZOLkWS7eFhHe2NAs+lGZzJsQ1
rPTJiBmpvdB+sgF680PN37YOPtT9FsCfQWq6YWdJztjfZT60Fi0MHYwig3fT3rRf
d+RMErQeVnMFLpuh3hE9fNn3AnvBlzE+Et81kFzrpjCIg2eHjLSfU89OYJtJk2bI
8OWEH2hIJidoGMymTq2y561DuoKumIrMRa5Kt2Foe0uw9HVodMhA61ll21O3OZky
xuXYZelJxlxwkmCLaU54FGLlDkQqBoE3FEyOn/UXRZ3pdBursPShOCYhpVfzFdsM
L5EKcG7tg1EW8ql0u7ZPjIzuHE4cMjF+BLSrud+W6yHwCZNyke0PaFN+yZbAbT1r
aeM8D4gLM7Kg2fLpooEfKz6ewZpWVoFDvs9VRe63RgnNlo/AA2HYxTKlGOfeRPcv
ZBMu1SG4mZxlAOFtNsqubHj0BFWn21BtSPt9epy36fDPXf3f5lNygTgdbujocFDZ
Jt3ibZ8gAKhBHIjAKpZMCEx4fSNFtOuefxjwge7rBQQCchMEh+WLTht7kYEdVSD/
GJVDT19Rf+LTcpwmkcnBTIrrc0jcHSzcZma/EG1OhNFZ4QtCllg3xdXB6ePBbfcI
uZOS7XWsa3Nn7uytoj8X37fL9okBsXbll243+oq87S/PS/1BE0yIcg4OAK6hckvd
W1oApJbY9n98H6jI4d6369u4hIhmgFAWGKHiTmPmVuk7GLQ/U91ZS0oIH2Oj41M5
dJqQthe59NuIkmkyaJXSJiIDPqvGMeVsaNyF/utl8uX//Gds4XCsPeA8Pw2DpuWJ
7BUjTIa7LkJdgcDIdxfe/dTyTQkybemyEQB9tZ/o/S5wCFNqx7cq6Y0MvRJAgoXM
jUnc4wWmo7BnnVX9jrwfZ4uoRFgOKyl/3jfyR4Cfcp2gKbcxKojgiK+XP5e6z5a8
jCJvzMrfzqwplIEwdrVEp+EjB+y48w76OydFiOUCtQeDqVN8kQtjHoovbYYFZQHP
5HvHL64VXBF2+vcf4g4ma19vc09CWznbGTi3bX1SQB+hrJ7gMs3qhDsjyIAzwefs
WTPX2yb1g1DjNbpw7f3VRckIDqAqS99yI9tnbwcoVcFlP2Ynfwc/blW8UDaoGxqg
EKMaaAY2IF89qs5ZVLAygoztzt4zBytv/PZ+xqRp2XNfYp9IacpUqc5kmu92iC73
DhZZuMiFwTaQu4X7Mnv+kzRdKTGqozRHyBljshuPGGZxHErJUwbl8SNRl4CsMvt0
CZJ/FuK6bhEBkmZE3TFYYn+O4fPAz5gG+cWEY2FbWsaaNlmOpvuubL+1pManu2Jx
N6gKPPG5j+NroOnn4xcf3g7CqN6LeGraACifVfnvo5B1HQT0JlLHsJ3JdL/qy8pK
EyFEBlqliddBPWH4Rn4psB46/0gUTg5D0z91DnBk/qElYT5blEwhRS1xmXK+ZLtl
odufn8a1ogCzSE4CmeMpv8iM+zo6sD64/1Bz0gR8ZkQ1/15sG4fleCgGrt7Yg2hE
wuTLzid86tfEu8nDncQ1Z76NWfNgd0pxKD1Np16QHCW5Qb0cXOMMixww/v3PZ6tt
4E144odGzvaP4PGAxAtNB8U/2AGJRAepyo4ovJV+Cj1edMPy713ZSmM0RHlF13o/
opFZMPVaHRTAGelxSy+a3UVTl++mjeAtnu0sVYKxiQl843mw26reO12vpCgYrY8W
IUGuPM0/T5bNROJk+ROmLndAU/faKtM/eCyXsj/TXDb1++PdUzIzWchEG9sQQGuA
m3xAvy0FhoxTmvDocG7ZUuRnEYGzGjLbb/Jvg9n+mbE3GRFy2FfhB+Mz6EEKkHBt
o15E/jVEEAPTGjcQkdtt2EbhfH0j3xdSCxTUVcibwnBRmSGzv9ZLFP1+/Ws2Dbzh
58y10B7vtX5IAc7CcQtNvBmMvCrYaoXq8zTz38tkZAKBiesyXtObFf8YZdkhb9gv
KM8FJehziOer6ZO13ciTrg/2Fi6CYxNLqoPOgeWCoknedVooYl0CR3p5c+OXDLOG
dFHuzZN30gxwQW/d/2vrMsm+4iPUXqGTZbkl0qKe2H3zcO6d+m704ojJctJs1/s0
CEl92DfhMkl72j3gjK+18mSDEuiO0kpciFEH/G10lQ0w69jhjR1Pc+JFTTqniWI7
6kgkwyT6bhr4ATc/MJBei7JvClK4KzRbTvjYqfoRuRySU998SnxWdVpDgANALVh3
9koZEVlWZdj1l3jtKnCtYs6fmNsHeS7n0DCWGaX0wPE3dDiZ5ecCOOvgh5MUI2yy
p4ab+w7/OOPJ+m9nrOTD9L9jS5d4P1kZcoSMifWYTCeRc6wGhX7bfW/OPl+ESpw9
V81ta6TZq5dbg/o8Nrz7Cc09qIymBBjymJg45uU3hkBg33dPSO2WWv0D0nuze11C
BdKNTMSaMqyAN8W1plyZmHAvJFqWFuUk1vnvxrXNqHjRQZWBd3CC3Wt6/Vpleg6B
ih+thB1e6u5VAWIQP60qnTwwR6/ul5PkffW8gw5XgUqXQVhAGxk80uRLkAjyEgBI
oxsZArfByQE9lJLlszi4ZW87q4FnpuhWYUYrpe0O1S4PpKoqRZ/XjD2XJM8s6ZpM
8x0ATaXuvMMhuM+Zs8v43Xof0FW8BCbl1sLpBAbD1Dkr5FvKeUpbNkUZkn/fofwm
CG4EKunUtS4RUqFvWNLkA1robIbJlurZQN/tJDVFrChDWxZF5b4xPZgJubsTkx4R
eThAWmyJuunfVaFF3aom/t3tL+Z8FYgglZ7m312LN8CdJE9AGpcc7oD6Xyu267aP
eBeKctO9MiXzvRwiTyz13GSB7fcuPoBS+51B/bPKrwaRktaV2haQDkPYAZC9xDpo
q8ysqN24rq7x9BRG1XTJVVrTVr/Oyx+7+y2zb05jVTrgoThAxRhQ+m2CR8e/ldBx
g0wrC8/fp01ZWAYrzqzZkpp372xdqS74yUUTrQNcRP0K1C4E0j0Qm03ZQEZrvkqO
Fjk8pcSKr/R4UJoKNTsJCbEdZOqzYbtx3FjWXZrl4N6UHUDR8b2bSqlIlDDHnRHl
66qx9jwqCvi5m5dn/NAlHSjtBsg51XJm32jBQuUoiHeR1RLeQSmQL/sewQgQyxpz
WUpN0i87lkCpoBS+HB7AAQ4VsG7BJr3CqgHJpCVyVrw4Cpx6EudEKQbj//S++vXr
xtL5JTnYg+1WmEyVW9+iWJ2sNQSS7QrC/lMwcGPn8CYyBEJVRJe3DWlgqW+Rk6vx
TJNjYY0lc42sDvhfetkKHA/MQAUL8/6Qit3DZpoh94oqHY2p69iw39F8L8+a683b
nWdHAgFhBcaBQWLQt8Zf7JpKBhs6BZyezPgKmIVmYWtXmS8K3B3KVrIScWyoRYGZ
yZhzF1a1+uUbNjnI4XgH5q5cKNF3BbZYsry5Ip8XFqEYCzGERWOJZ45Q69H2P7AH
qre8xB/fJPR3PXoOoPe/enjz8JXcw5wC5pBqPR5MooO8aAFbtWuQMSbAG3VVVv1m
TJLeFHtT84q+1XHpHgwYp0q9GV6RjrOOv2NB4Z88DF3jmxW336jaLanlEsfpxgwN
LvZZJ5JNsGE0qXHSVGQJT5ymwYYUOhZa2o4pW6roxa9vDhGoH9d7n0Om9pXfdWYj
Ej3MeSCA4rMqBPWjSXxlPHeZkKFxuZZN562sQRyTYoCVxp1waPxPvFjAPrSshYPX
bKl9cXiIMV+8rCxRDFj8wm4DibPXtI6kFwEkqEW52cFKIjSoPIJTBx686EnDXm6T
TkjK//Yl3rjjy0T5TSMeAbFTKUDGSk+yWhFkGSqM7eczHsfHiAlrZ0aC60r7cOIS
yV604abFfjVpfMP4329qw4r5Pfb26GS5RZ1aGyVbL3S5E+Qwr1NjKOFA1BOYcRmm
rbCaFw1tjpqtn4f2lCPhrWpwgu9yndAbXo2DVnci8wwpxerU0yT4JAPkR406pA2x
okDgrFfPZVTRhRnNDBC++q2I4oBiFUcaVLZ0c6ddTPxLa6q4VuyP3O5cgv8O8V1N
uLvNIQebtvKuelppDi/IKcXHZ4FWVWZJmBN99cxC/Xf5Q+4Igm/I9AnpTf/3DejD
Uq5P0Wh+64PubW0ET4JqSOqEeOGfMdx7mRu33cKu8D+kjgwuvlXhbWRgPScS9wFS
9z803oh71/57xwPNvMLb6oVxQdmiaDc/gIN1Y7kTkUkpAYvID9FVTD65AN6gfOcB
oAnY6PKy4k8GjgqzOaFhcHaC3+BHMKYi/2j/gmLYAXaDeUcuD6SlcrfGuumL14LV
izv3id1Xa27jywl3BeupwxwlJ6KaA/XO57OfGpGpjNHtQba2Ff6PUikETrugQGM+
CUeXFbsvvgFGevB33zet3IQIiA1wnc+o/WEjuwFrkXYat2TYut8awN6IgxAjgbHE
P/ZHnFm5tHP5kuGK3yG0DOiLIMm90l1iIGKcMrngrVKIEs0ZYvFtoYObsZVmQSh1
j0DdjZGBzWX6BNkya++OF+AUuxB5qsPVo9bWunPsysnhV2vGB2c2H+OJMCRQyUMW
LlnDmhkg586O1PDOIUCU9a9eT/5e86B65CbtPWr9Pp4XKL6LJ1x70Kvh9CcDkcg8
IKYiRBOsDFQjWjJ15tTyxvAKOFujxn2r4ChMXUKvrczLAepwRQgY5QOzmei1KPW0
VorNEOXLp+f/Hm+htSC/a+6xYrCzgU98Y7ZKSq1xzt8yZbDvCTUB1fslPTBOiGGv
ylZZx1JY0wKdlZm5J4AvvqxtA00jGau/69plp3cDBaAYIeD1WZ7e5BHifWZyXcPb
8YpRYG/SARX11GEPTDFioFG1E70krMowNxvvlmiV/g5+27SPafFNHBC3ugiv1sy8
J7FOT1G2z2yA75ryF4IslalWmqDiZN+NKTPysiHqQHb/a0wqIAKVHgbYGYW3E05V
m9rzDsbdMxryMKFSp0rOnz9+Xy26/a1WJzzQ9DV2GuIxEYN5jHrZeOVKkrTaSRd/
Q5gSPEh0t1SCVJ3AsLC7vB9zLN9Ppx5/yHJD1L89j7E8p/AAbXQ/QBfQ++My30iJ
FTsI7Lk2IuhUa6mLO8Q7LzMpOi72xcKblUYvjtyOJ3XTIlsq+YFG8XMxqHItGQVX
kaS+7Cm3IEZnhFqJk5kMtul35kD9LkPDZ/2+RPXDsxfLB4iKQwAZxyDT5bXjcJ1u
YGyiXGw85KWd2K/P+1pO2eYxow8pUXO+ZmVST+sUoMzLhTbOYy4EXfb98TrxUp72
DjY6dzjvHCQzJPYlFN4JjQRXh3SOrJtRkDbl1cibJ4zT6xg/GlF14FkgDkS9PzRj
NkosbzSfBT2fncJN7SswHmptrgubVq/98+wk7xaMZqnjgwrpxzGiYn5cURtSpPXb
qiylsy58Bxo0Hx9Uzk3zuDcUPpGf6Oi7TaHTOHsNFvwsPeNFgSqJ1ZDV7mlQ3WeL
QqGWXxE8yw3vy2m6SdstE3DWculL8DS2EdOCveeic0cyCB0tfAt9cxMB4O1makuV
ritzJnKmZTihPgBQ+KRCz43sBzOC/1HAX7fQjJlVvOHYsBLD1FUCi34RpnfDcTuD
3Bw+oawNny6zJ20B+bsfugQg0/u9v6hsZhnccI5F15yKKX7Zbb7SngOtkpjNnfo+
COQhawf0dcNE+u+GttKUwrf0LzhFCTLdsbS3G5CP+X8c3oTcfYFguaCPF1m3ctZx
G91cXxb4BCxAPxiYEmettXseRQ6rcfH/eJlDngKpSy9HOme02pnX3xCIQZO2bS+O
AtHDRiAwMhzz/izoPAMbm56dx2u2XogMnHnM+cJryrrX+p093/zZa3V9kXnYsNkE
+OVaLxOACzjzhaUqqyaS5TvMtUYspGvflcKm0bflgFEXgMOoJ/J/6IHEdzMTYbRr
cSdwmxwmZ1nq29PnSKsuX+prdxo+2y78weHpx+aTPs+RdU2Ngr2nwI5j/K6Apg3/
KfwMTryAo/hKpNNbHcnI4b7vUtRPxRlaH7AOwg3phiex9yuzgEPC1vjyVRO3qNLx
ndTUXGbj6uMPQsPdkKRC+zNyYwnd96sQoaR2BvpO4hYnUcwKPHDsrPwjnDABwWWE
fsiAtqRLlr215J9xkqo0X2s+O1gai1kI/tHIzI2/02Get8aY+3qixwCuRqB/fkQq
D4EqhTXkdRZAFelgS8UdrPht51l8WCLMchPZvUA7SJZ4RZi3J1Yo9A6Ik+H6jtPj
Jy3nmjjvWLUqgMthzgrbWF8eZcnqrbDjlEFKK/8urvlwNYQXtuxk6GiNgTWkynsg
k6TzAuFcFw4Zvgh9oxvEbHSqrWphxhmNyTwqvN+ajtMN11vnVD0x1NoRf5hsdGAA
J6CI2DPg3yMXCYeo1l2gAG3qOL9MXGGmXB+QMgihqYGvFWHkK47144AK0n2hv7Cj
vyXVEyOEbl9e3p41ISr7uBZjssxuHM78CgGtaOt4nguI9AxWr5TYTsYfNoSTYQU6
/Idz2gyt4wkVIw96QBj3YMGptOZetobzBfctdpKDfeydSeAW0xc76PeZhLmF8US0
hZonLQhMUnFmPikmxLv5e0IBTtPOTxhORCKnZGiAp9ujMa8PpXkgxOt+CsCTRWbC
jc92lbyWJCe3KrtL3cKGKtDZCbadqBifbRe+Gatpmlg0F8FwNXfbb1Q1urymIvPZ
2iZuuG/8Yl7f3G21hQTKAOPjLxVCEc8S6L3y/CyJs/IYgl4BQDYPWUqhfUPYQQo+
odeJVgiP25lZqlTT9rSSK0ZaoWHbCUKARast+kaqbomnkZLd1cA0RNRJ7NzE8UF1
ZF2PB7j5oZtpdTGdQ3odGzT2XetyaUql6OmqmovNbRbDwiCvl9dxqNTxAYx0iAaN
UeX60mRI3Qt98PZIpKOx9gDlOPHbxfLdNlEbZOgHT10do1xQZ6Jrv8YFp1BFMUzl
r2oZ87Z1+A7fcCrTisHuNI7/CSmmTDhbGltZiXzRugEIjbYx99hV3zlShYTUGu/6
8W3fUDliEJfbEr2hHnyF0dPLucrwnVjxDt5H/LVlvL9QiauRintBtGV/19hmbKoT
UW5QvPXmh/+bS+SlLTV+fEpVoSvM3OmeOet1oeT1g37EEu2unlMov8tu1OcvBGpt
EAx9LJUnpgjPluspF0ffm4q6b6jcKcmKcbfZXU6bAl59QJ61Bh5e2Az4fAjYLevw
cRtJZNwo/qOBbwSvsd6VRPmIGw8jEIA40r5pj/5bIQ58C/kJeUHKl5id42lW5cj2
4UIbwkai721d4vxDzjdHkIy53jrXbcUOluYPof9WxFmghUf3rU/PCi8yLexLbY3a
D23Hj4MJGXDI9SKq41eGnSorVr+XW22kxBq1vcRVbg80Hp8v+ACddVewOgITWjoA
BteWqy4GhHxeeD2OPVGjibS8gCzfm/EXwdAMGcdGZGfJ/1BYOVQN52AgFHBEYgDv
kEbKbnRKuDs1jKbrpS/ROS6fEtoXeh48eA296b7RNdtOoLV+uQjO6KuYFJ02fczU
11avnoqJxZILYe38RNbGrx82tqWlbELFQRMNWhQbfdLMl6T/Lv96Cd2HklRrZ8Q6
ul4YF1ZFdhu453R0LA9vD8+64z8uncbZexlnbrxAxGGKa9iqB5AodGeCB7K2CCnS
ICMzaE1sZUsHIRLFr7igCIeyl/BagQT+QTlq9gJF4Vj+NmnmAWSl5Zp87Te2gXDe
mOg2+Lv524wUpIaMX5Y/ZTTdN+vXQKbHa8FxwVws5InAJS1mCf/E+c4QpuYCWGqO
xBSo0BgLaIH77/r/+FnNZlW9gjso7HhuUVV/SAv07lIjkHWQt7QLza2Th32cEPgb
dC613V7TSGD2QDj9gY03SHdTq+6bw/UZVFnkv8z+iwUIdiXUwT7S/jF7SsaRc2/q
BldZuGBA6pAlbQut6QH4gtTbeDNmxGLSJGY6wHf5Y8ZqdSt2yUBrIjd2mekWIR6G
znBG6NEEYZyg5fyHp5Z2+F8Q2vRA47Xy8PjjjjiJFvuyybL7qvcj1wZ20SUmderu
gGeK9EHg4uyCw0Bp7rM8gjjGy1aOI4ur0GcJUz/mWhZOy8uE8mJPaULH3LJe+zVV
bb8mKHrK3bSqGqmetHz7s+TyulGArevzJKM3JDp6eKIu65IyPE84stbEKDvIXTws
hEyexQxiXQkTCjMjyq3k66n9I241qDQp0Lzb+fyRysVjmTfTUdIuNtI8h9W2utH7
lFOyhng6/rZsql/kJsPzEZgmB6DTM7gt9WyHTW/l7fLmsDJx74LyhmytrbFpSPc0
73sFOfF8XmZaJ+QePkQBztXM/cma4R/dh2Q/O/jfAY14G+TaxcBSwXO+DiMlgIYn
cb779wCFFS0gLpAv03d8yT/C5zqrCcU/gG8NHeD7cwPemlwtWIY1kjfvk7BJnobZ
pQl9D9DK3ceAVxbpOj4CyNHZJb3QAT6mG9y2dcoLzT9r8cfRzqhyZrV1vvSDhxEA
pj2CYwkYGjTzQoU9gBJeI0s3yvrhgYxA153883RZ3s+reThJdKN9yKBV85bxsPGY
WM3o8l5ZMQeJNUF/ld85LrkoZdL54Ofpx1W0xxppQJVrtcs6YG0s3yaWJq9UHnKG
Qjky/k6Hp7Q24H8tQCKOVIUzigpobY3b4jnIZlpIc6U7oJfEbxjDBFDixAFT4amv
j9Y7C6s0uX8Lcik12bZDfrUyJacW0ej/8V8JuqbMcxMULKAGKnl7jzqeSv9GNkCv
S3tEOxgkD8LjD4qa1OeNC3M6oMo7r1iVEmDTSVz2ce/5Y48j9jr9LLkc42oCEfY5
9SdemrL+hxo9OB7JudSG3e+Om7NTNl1AYmDU+AtMh+Oo5fEDHiShRzXeAqrfhIVz
eYlBfd1v4Rx+51zuUhP+mV13VQmN79o4cI50opNa4kJhU6u4Pvx5Nfb84hQt9wjj
l+C4/ewRfcgsmTGna6YcGdMDQ7Uy8ppLas88X5ZMfqu+tVuaISKX3azCZ5uleeHM
7QFrxh6Xb6kQxOXs+4LCL8K3ngB9VWsg9etHsZOaccgLdlCnnwFG4aybtARdQe1H
+NkkIck4M8m9khORgZjiM3PAihqtF7UUr5zOQM4g18dAdbbP7ooaLkmAHybWIIGD
pkExbyOJTV04lp0vNXrfmQBMgZlXmNYujZEpbVmEJcPN9yup5K/IMVEVxQsnp1dj
dwwSVHu85exbJabqrACnbxl9nn6w+OKs/C9pSXbp/tipEJHOkWSmJ+2p2HuZ1I6F
F2LMs4to3DPH0auU4CsoLGP4heZCus4vlSw3cQ9d44G8Sv5WFzf/WgV9vE3tY9I9
DuKM2wYdhK/FnyXwLJPGonXqxE8QskXL5VWTY+qrtzFFVUwpK9o6tYV3ybKCr3DW
ULHBTeb6fjxqPXbBpgXrc31O2DLpqZ0lMuoW1Jn7yQB5SS7h9Qm8n3qSnHY4Tnhx
MoQEYWr3U215+17lsCZxMGkBOw2px4gNKSxi/RfLmzlwLMUNBZV9m2VUT9k9p00r
krJNOJ9Q36Hh+LLUgg6DnHufdLuJM6O5gy0RpALYQE8VNkXbWDgpybO0xGKWzc7T
CejWT6QYaQ79IrRZhT1clf0b5Fga+bJpTubRzW/PkPl250twlJd1QdvvIMidPbp9
eiTNLQm3BdjHq/eiot73pdm7j45C0WX9WjL0NrLNPeFV/P20dG5/4TQuUPOkPpDm
L2Cw/l7uISeY+A5XL2jvT0CSx2Dge7IuUifAQbSlzKNSKT4GaFU2RwrsZ1fo03hw
EldD8MQCNWUwgl/2YvVI5nvp3JON/U01YMZAjMo6Tz4sZEgPqk+9PbnLx5mhT36M
PJiKIb+L2dVXA5bIE8citpzHs0xKqdp/nyRrdQp9PUj15YBEa9wwWTyryDo+YdXZ
aeS6KUSDG7+bDXNv+gO1BFzbhjg/pG+y1YHpqGEX+2aP9IURe8MjEV3P2TiAw4nB
Wi3Q+p+MlVplUw0vsvr5ur4sCfg9VkcTLNlQwbs//rm6PfpU8kmGRwMMi+SKHOcC
+Sw/4/eNUp5I4anlzNCJkuWzCHmlWLSwl8Wi3Qywa4RUr1YxEGd6QkKXjqO8BZgA
nSW3aTCKN0b968QkzEZ8lBwTZhcrMvHf1aD/Aq+s9KeaZxYgo8sd5GCpUMagDcEO
R5fhO/6SXbszZx4q0B1qPrI0f0G6u7PNwvCPQ/RoVkeLU3rrlluGMmgEfFopy01/
vKWVqy9Gq7GJdPfk4AT/ctEkXm2Pdzb3wDZe1HMEpPdd3MHDnopnGArkQfcVB+kp
qdd3233hUXez1bJOY1062qKPvOyJ1PCyEKrwwD7KsXytyZYw9el+go6sWh/QXiyi
n9oaIo7eH6p9l4m7oEQsB0wTLc+JxR2NrpltX3Ih8O+XvKp+HjJ+OTL0iWpCKcHn
/uE3PHVbIga+i/DQ8pQosEiNSBmbdZXBf+uj/2dUKJfnl/penL5xhtAGVli1JSD1
aVGWQBgs5teQsfn8CgHWuki8h8yXdXbzvb7hC8xf61NbgucDOXMV+XfeDfs5tWk3
2B86Vc6n06X2KuqqwT281dyVJITYyX8JZYWcC20bg+pMoCNWtKe2zqRZ2xP6MmBe
O2UwR38k1w3ObrNtH3aP/2BD+rZTvNP/39HAb7FPFZkyjqV2+jWsJN3vsVcpRRi3
gMc7BiOtFSTW/0EpEXruj6R43n15OsbYtyKKrVTNzNbjsxaly1tMyvOeC5eeG0Hq
7pnAIV1zJLYQBWFSuVeO0fQ8Fs++tmS9jCYTJBhEGJwp7xjHOVwlx9XO1589qHKZ
VOAWdg6aPaQy7zc4OGPbo2c+CrbZyog8Y745iLa5WcDJC14blzrLL30q1HHeeVVq
zstrunQfMn0RAkJwRwvuW43UCS8QqCLC1kDGdtbwkzN00wcl+QQ7UF0kylOmC7fe
IkADl1YwTI6lQugpm0fCbhZsmi+RC+tdjWJI12fWem0bEr3GG8tEJggTpddzPQo3
nAAhvCioC6GPb0d8UkxkbdtcB6pwmhBLJWxf2M5ZiKyFqGRN5N6qjBoc3/5yQym+
1qDbNi25us80usVEUssNuA6UjzpwVdzVAoK7hghxN+4UrL+GP37P/LDvH/loraVO
XIwTdp6ue4tNvSV1ik9qGcT+JAp24wjF1Wr5EnQucwMhplnZzlF4DrxSUweoM2EI
glBeP23VwTSBadMnO2pn9b7o0dkODhqYQtDbFzDWW+Vbn0eC/7fBQKeqe0CLhBfx
1Y6hnWkhjVqGToDMD7ITwY6GgdQaUvUdHN7wjTZpxFi8IBGURgu8DNKcu9O9fXHb
duFziq1W6WnZSlAsJQ7enUkdou5OIJkAzaFXjALv/2Cm7TbL1NMAOICBMhDubWux
Au/Dg59VVRus6ZG+NNGSTusdi6xJFt+paxG5xHFa5k/YJu5gNk+HqeSX0dtjsEWl
i2/51/e2PAarTrCIjaB4oj5rErN98lvscOi3Ed6S+cGR4Bh4+j2u1oSixsjNCO5K
cI7FLOI2OnxGpSwcfQrRcvBVJMlk3qckFk3VZTEj/11WAXV54JGdbf1RUEpfWZcI
LorGRCRelNewn8lRV4SN8vyWNURKNhyAukVDsFc5L3EUFZM1IFiUNQCOrAl3ZyX3
oqrxFTWp+3EBNVzw32cArlb98IrcFA8y3PHDCY0ykVx25QF7TpdDmqYstmozMWcK
td7UjsMx4R58OfY/IKxstGmfVBw/NAbd9jbNTWQa7qR6CCAwMh9U7d+DEMMvaQWy
fnCRr33/xm9gFI+zBhgIyCaAaAdVl+KECATnjh8PyE2/y+e5pta63fJCyVINrUhg
AsMfZDMGb9D1WEYS2uoV/h10AbY1bgt2qKqjSPaEKa5iwoxBsxuBOKvav8xsTgO1
WXuqFHBvYcdDgRzRehKppO2l9A9GLI8nGk5QcGJLhNLOSrQE/fJs4CEtwKi/McWq
N6kalAo9ywklOYRx8kb9Ih1I30aD+nHISeds+fcMhdDhgHaoMg8p3Fu0U83Ad/Di
Rk+T7bS7HM2WaQhl0g59khLLwaNHWPYC7C30xwY7e+vHolLDVkgesPEoSl5ZAgoQ
fHMBU2zr4bSDQrKDFmkcRtCv3Cgrgt95cl3zKanq+/6GsbSvmce2mzs2sAB0g994
zH+ZxM+YdngX+igFDKracRevZGl2rKHhsz9rAYawat6xlIKfuY20uz9gqH1vQszn
kDlIg5/VzDM5+MBys/c8HNFJB2sz4eOfvWwNtVxgl6U7BAhiczO9Y7BPtm5oZuGu
H1OB2kOpyYvSbjnzo2zBqAi0Fn79GVAvoSptzovpOZywZQTQstzgi4K/XW3ml9Bt
/iNnu3MHacVgC3J6w+d+3dKY6MfLOsrzCq7ccLWLmXsoXMUHWggSWeLXxEUly4oa
HmHvwnfZ9OpMMq0i2ucZpbmVx+AsN6AzNKD1Qio/6BYIYipLsuLNC1LpBEqwdDin
bxbSwdfWP/3PMEBAXucB2iG5nYAkkMh/AkxpdtSF5nJeD9oW87n9Fl897Y297faZ
jjLY5el+q2Uf6lmSLXLwjCD/L2R2mYqTw+m+1vYsC4XDZQ9+/efT/2gukDN7HcS6
dptHdhwcm8xPSgy6dSsRpyhBHf8grNmns4273HnqNCafIERQTWkt+OYP0kFXm4Ro
7r3RAxCYmuu+c7t/Dmv3mDpsLAHY/6NrFiTdCYk1oDc7GatSSn3qv/TR8zmHqtd1
r1l8fDFXAEYeYzNCJJTr4TAVlIYbmWzb1gEf1IRslAPX7B8jq4o/MWo61pQdov22
dptR2UBLDfCIhH/+0inCUrGQN/fqEppSL+lMD6GjSqyuvVYm1pcyVxxiLLA4D4VP
qwQZZoLv+GlOobnCOPKk1DR8+2xEJdUCjyux38Ll7/fJTnE2fEgz/wgIc1HX8F9k
IokBGyfst62DE/sfYUVOJO7ArEz4WoOE1/PqHVNV1jNmn+VXbkgIX2kp5+zVRQcU
Fx7fb68FAIY7iTbncLXysCElLbYUi75voHt/uy378Nzb7zX/JFnSQpCKYcYV9uza
DuqfZkFgUm7olB9d3xRR0yTu3KmPOlEaFcwsX4bdg5MzyY+1zGJ/9zHnFY6+fFjo
0P3z6Hy3NDbRtcrNCn8VLARNArvsz9yTSAP+ut9DinNfpgTls9J9dJ6/VMTSltjp
dqJF0LqCQU6OgxKniR0VC6zw63cKJYF5umE4bqyvVkwYWXaMA/nT89KXfTlC3zm3
TbzU+uyx1VzLRxoUdTv2iF/CvO28mjd3tySciEVQG+tN3lmlwL8G1VThUH9f+nxt
Zwj8kc+qIox76TB6tbuK2ws5dbLtUXHbyFXcEh6sLdLkNZ6khpZcKfzM/HRMghcB
zlah6csh4ZtE9pn7+fQ2Dbt12ofKsKz8hOiPTo7pUtMZgbT0xdozGnAhX0JLnTII
18ge3tSLHTnxXt4ZcM67bzFGHtxX9e6TNPZWh/aFYaFQtzt0O7piTxnIfzuc/Tdk
hdOwCMkPdWP+nneBOYVQ+UPtrQOfwcraZlRh0MU0t5O+sJouh0MgBXH9moijpPWi
WyTfSEzODFSn1ajVvwHVz098UZJXdBqLlx7aZmr+KjuyaD9aRxhASBYaHCMJk2Qb
6esDkGO5fbNAmTNHp6tGO9G+cH2VWIO3lMYk39rzBygHLow/aGwYoBZ9p3hCX848
5Af/bysO6882YpeWH1D3WWLynZY2bLXsD6wgxsdXxeG9iPYXFLmiAuDDDEIm44SY
BzU2sLrdJ30oZFkzmMV907CO38RJ5nvGHDyOLKFhv6Eas7tkIerl8bW7HSOlE3Uz
olhsRWdj/zajVKVB5rFNY+8eTiTpBw35LwRpVsZ21wLB5MQKiz4690nRw0ShUeXM
pOp4X2JImBVzOWNgwSDy4Nv5rwNqVrBnDWOFUZwnnfBXHyV5bKq2HQDWrfo4/bI+
TeLNMJjj28ku87H9tgIz/zVIkAjEg47HZZXfeX0YeuL7PVeDhE9aeRAPSK66TVzg
yQ0Wxj92LpkKGSvAKBQzcyDgzAP20bIPFmR6p4f4Uc7KY92YynT8+eh4qcdDdZjk
jSROr+eS+ZxcCIe2E4P6cXVQtuGpnr8ZfmPcRyXJXdHUeqUlHI2pKxTfN0lmz0J1
XHh1nZMHVAxuhV8rrAm3g0IwY9r3UfFrKdqvCJW3UX1meLQIPyBIgYUf87dcqLst
p6v/THnR0kDbUVFqWiJKJLMoZrlA1aIb8ae7SpVZmxWXjM1W63CEkxpPPdMhDWGF
RbZpAeULbLvxHHijWWEDGUFtyFskjn7Tz/5PwU88mRbwOtFmmHPaayVGJziNlEO4
3MIyPwKeOG6UtEC9V4GmIdE+IN87kRKSH3I3FDjsbUJZbiBnnl0pgCLLDn1Fm6Ca
C9ACd3HhHfdyEJChqEmwh6zIiSf5GZP7OsguZ5z+Kq9rro59QJaG190xPa8YcOy6
gQKvMiRDDovJbLGkN0tvZkATJR5IOkYGwSkJAProUik2Gubckd+JA5Irvi5ucv92
TfyqiJRu8O/7mRjxeTLsPNOW9FOHe0FU2BGYh9JlUcmCDz+txH8z7gDN3fgOQWbO
iJn9gSdD0A/UsInvURwMZ2ad6DeweI9SDeYPSq+SKdGhcWT1clZH25pfnrTbqjIU
5GKzK1TsdHTMKel+qf8CSKTQ7cZ9KbqqAso+ZkCQeHcsPerihB+n0+9JJR8a43bS
SyWOFJJSDapxJepiV8ETy8O4GDqiKYbhJbDHrtTWqil0lJ9+jh9njHsrVN8eG1jJ
9szFYsoxMkgQX0zpv+8ypem+BQsI7FnGAUQ5buWAN+dhx54cjtXC7S9cyoYq92kO
scyagBf0aG/cgGTmbrJODp0kYvlOb5dsE/Yubv49CHZqjBet8sDGHE+ww0GQYOZk
j3u96WSgI7F1u9unDj9X6zliSCTeWQs1rMa5M731mNk9B4t2bOfyiuHTXnXhQ/Ku
2fFVg0t255Y7x8kS3T55GwNQjbhVBGbhtua6putN96OtBIb9OaJG0IcFO6f3DT4p
8QWzjfhZ6WS66mjwsH2/hEQsLV6VvamFswhxJog9UN/lk/qmMmeZnZITJkqSw90X
HyUTmlHn1qc+/+W8tQWmi6IvPrE73t6bDdDnS7gwoKgo20Tc20Sq0JxDS0vVMKw7
BC5+TRETimI5cKnnqS3Vbp1wR/kehLeLsjHxLapeONxRWRQFSL98NYvRlvqqsysE
WSVOxPgwdg4Pb3lw4IJyHj7stcz8a75MzX/khnZdJ3jGvzKJfl98ySw/viYqaCMJ
t98i3uUHxdA/tsWSJ88/RhEqRm982A8FbkdXWa8tV3xqqoVaOWNRIDu4L4eW1kNz
Whue8jva0+e+rhdKYdbcOEa/ShTnLXHrulQr1xabKyqeUJYvgZih0d2o+x+Msbfg
uZamv8Priwt08KnASbBg4LgGXVbTXD6Kmxf0UMgPlmj7yMj9yiU7ist/4rh7AYNx
Ef8gU4dpE6eTxIT5z7prKj4XtP991IYqrz0qwKbUXpiMgQ9NhsvITRJDv2BoRJUq
zCejlxs2PeurZlhMVwGelBENAdawXju+biUb0Vd51N0kTZEeukjVDPbMbFPwg3VE
28mbFRg99HEPzzOCKXVHcB2MitJWoeqvWYUc8DFZ5CagDsZMFHj241H43BWWKFAo
CuZEV66MWoys0pHBK4omc6v0/ymL/cU0GCg3VEA+rukLnDCMZNbu8lQSoxFr1bCo
YjEm6BCke31z8PwkaQxsqsJafXnzD6cRgVa3vZP1b9ImXtd5U+LT2EuyokPdVa/W
b9b5pz7/XegR+PwwQVUvJ4xPQCyEv16XzVSoxAOXJBJuDhi8xoOXKqYulMPt4M/1
qh8Qcv4CZLoSN/ApXf0aSNctcvukAyv1imr0oELs3Fn7h7x44Av4QGRL5XqE93nY
z0NtQBcR+FGkcqBcokhs4w6o7Uv/Ws2Hb27LZpFNWr9NNZmR31WQhIlJafzGAKCG
s+DWFvLzm9AQbdjz7yeoFTDXXA3ZsYqxdN9s95NSJlcG8JEugSuP9eXTddBT84Zk
4K07P/BkIq1LSzu8PKmDSewNXCOdLFCyh5ARytkoFEDd4O1K+0vC75SnsDwqo68i
2SGWfUew7Abp3+Rh/Vy5nTnFLMYWTgY64Pv10cOK7ETMLOMpMhYbOEf6gQ7CFolQ
PjxYc5INrLZmBCZiPkmuStC8sbkON1oYAS5Wvs60w1MfpoxTyD02PsxI0XyR39n0
BIR718RLt63aObZwknIf+rv6vIFvWvDThxp7pG9NTNWasA69YqogDoJzfX1pVqO3
EmQwh6dnATv8ccehL+P04eZX1UqJbEgeni+kKnC2WwT0Q7wzWtSxybYRulssfLDv
LzpGtj3TVh2zkSQnkfuxMJ+hj89vifAUxJ54Fq3AyQztpUO2m7zpqoil1KhMwXlO
HjtrWF+TxzFOsm5fZ9cBn6dy64aca08HqpVBjMJTNvggMr6PJoY5NSnri5hWsQVn
jmZfqsQGeuB4aCeDfwO5un3ZVOE/I9owrfjNQEHjFPXixcqdwUNIdki/KgY2Z/HI
Nyi67VwztLkIemktjogju+1syQuFwOuK7O0DDA0ptG5u74TgLLrTZFJiwTjeUwwM
Ig51V0JFSksnOp9TLU7dhe9r1CW9sOwO2GukeYECJWc3pgZZa8nHp0q1PPSWCnRM
h93MJolxVL+ZZlqhY6reAjC8VbOh1aClQeK0BN4wZcyWLA6l9zMA8L6cDQXzYsfV
RhxNBC0bFn53+dc9Zo4/aAeicXzcbHrNZK7K7uSAHsLuPnZFGdol73zsjGhGKUKk
3mxcR/MilsKQrsUdHajeBsqg/uKx/Mg760hyYE+s3jFBi4xM+2/fvA95JEOxCck3
eWKf5SkMGw7ksAWVcbaHztpvY+VGCH6pu60IEuTJ1ZVcTRkofZHh8+RA29WYBxnc
wv7PrBIgCqi0IQ1T98KQfhoqEqFO9epqdc3V8NUQytDB9AgfYyhwvEkZPx+8SDAT
ChVF20k39bqwdrTyLzSr6SNhV/wAyQyxcuRHpwknwu9tqDDJtqU0i8wR8uIvZyBA
0zd1MJscTqTiABBB7MV2ehBqzXB4FBrmC6elEgr9og4MZceQBTbOR8fWvaHHYw0L
TPQgVxDne7dxuZQ3j9n3GcRsYEBq5sCYqjVwri2LkpUwsRPxa0zq4Mt/7ZowYtg2
zaNvztijUoU3Mo22XFu+YMS5H7Tv20HdfFKey6Ipn+c5MI+xhl9z26ZVhOhlsdIY
LSRxkqYtyiMTUlk2NiZEVtFolii6IRo8cLBF6dQiqciySax36DETgFSlTBir9dp3
e1Q1/uMRFrLdPvoFPYq6oCiytmN5g1YRWz4+u43q+B3PXjxlC6eEVIwtE0VFWY5L
byuqwzlbf9Wx00EjYJAoD7+LoKs5fRTi8C6QM02eTPTTr5JP6zRB9xEwN7yi83dU
gKbwOxr54dGoCykZhw2SudRVvPQK9iRHCtGTZ6ZGY7J+8DLaczYyAk1k289Arcmj
tFTA33jH1Pxba38bKTrqNq++pNPrfbfKXy+mNV+s42ZD/qaj+nP4k5C/SbZ4CjMo
YysB2GzOMZIm8hgzAOdhpwffdhmIJaRExWYKJkjzRXlI860OrgoyjQw2FuP0yTnt
SlsfQ6YDjLdjhx1k7MUObuG/ojUvCyLrNrnyA7Lu8TN0hGexl1fGGO5EI5LkSatf
Ki9O91S+z8YfRxZEiuAOqNEoy6v3pgZpSm6qabA4wBPWaYS12mrj5S7IsjYPJ97/
D9VLHoXcIWbkFDDFjc/4DW0Eqm0H0tT76KditBg8IRxoXsXgY3Z07BQqttAVBIA2
zMbH+KLDThjCj4c2NJj9iNfBn4V/3k4d282SgZR25eIh7PlYQLt08jEDgtE4ZYC3
dtZcydAilAa0uuo9cNdyHDinR83PJotWjYDhmaTiMgFwWkdWELmFvli0LZ6rY4u9
2muK2fuwpYdguCNQXmfPpXofloO27/Sdj3fvieHdlX0RUzsdaLfzoxx01lpTCj+6
+QT+vXGyFs3QD49WFUFNi//XKNrbIq7rpI/Xyh+O7hahjd7aCflhW/s2eHEvyA6V
qZy0idS7HwO0EH5XS18NMCP5gQPhmNBMYuGSB4inEjehpIpxPp53tZq1cMLYukoM
YLn4Ga4cpx34NYVq3tK5AZQbO2Gqfz1+G9hWJlo/LxDP9dROdhflai37wIKYUmuv
SabClh44stahA1tXzK5594Q0BvLtDpgdiviU06QxtKfHPVBd7iGTlrHXxB+SggbA
b8hh5HVEVQN1a72G6mBiE/7yKxAHNtSFt6qqRICStSHrgefFmajCmTvUZlze/YAj
DBLtElZyfE1MkHnTYwoyPdyj1sp50CInzompoIdrQWn+oE03tj37cxyclx15384X
zMtI2R6HV1A0HQz/qY7Zmfc7/tuB9W0k98pAuoHCc0b9d/PFHgJSmWkXvzUsWVU5
Cva87spl8cwYAkmnrW5hHr9WgkMZsSOWgVBrFjdNQOqrizTqW8ri6JU76ToIukgZ
uBxCnB4pi2sl8sSWebL9VVuLtOG0xfhgCRv2saD0kPBBgWmVxBFC3jnHPsEp+HLf
ABLe5vK1WofM6JtXANx4+RLr6TORNuNQZ88DQMGtjUcCz6E2z62PJKZIwmt0lvrn
5D3RgvzwOtcGrfzmqO305DwWCx4/DbjrVM/QNuacpRbCc9znUIMl8LLo9/l+vb0B
qXn3GQo/K/upbsrnkXP45JUU/GR3dHQfmljMwgu7qjd9qnBOdPXJPv225kyc5/Ad
uIO9me35S65HkSwmEBcqe7wD5wD1R6NgzEljdGCyk8uzBLneNFyLEOSh1KBxAUZQ
6RobDsRyLBrwIZSoxmNgxRTB3pha1HBfEC3BUI8nuUlhJQkIH2+CPmWlFXknItdp
Vs+tv/99cIf117z8mC/iTkJyBlP0dsAswF8eOV2Pz3ILHWqAHOT+0F7mxa9UVzzO
cwkorl6t9mkMwA4n+sqC3aDZ7OWOZg2wm8rAwrsCEsh2BnU9aLFr10bHJ+hkc3c3
Qmt2t3OPy8L+yi0Gn1rDKyusE2+J8T87UbG1izEvvJuiIJK5Jc3Tyf72DdBZyHAk
SOUcfG5Lq8okQFt/I3deNEqWqHYMQC0zFjetQIfvUUKQrCpReyJfsvCXV983gMt3
aAiLQ804w+u5FbJsPtaY5y4/ubvMJcQ9TFPU60Rp9gbf5x0K7YLuHxnGEPa/vYmr
HQ3ImMElp8nq+Gx4NdYMSOnGLiyysbnFTBnecrNz4AINkGPiJoUFdyiA3NGfpcf3
YJPPj4d1tWi3F+pOGx8Y0bhqmUAR/SQBdZZZXqIUlcP39YU9eJMvZvmE6XQ3EaAs
5C5bwzYkHGgAxWQRktxwfp95AoEaBBZh80Gaj6xaKBI6SX3hBUJhKDXLGWpUO5ry
xFvjZQNvzInf1//TQdeih6thbBlAxJ8at4/BFPwi5eSLX2pb3v3+jZep9l2+wSJB
LYL0oWPUsEXYtxRF5XkEnmWt63cwTgU/xLVhgpSIEW6JjrgvCgHV6ef7a4yQu5oq
CYeG0wRjya7Wu56hBXYFEapWQdnfOOs7YwvZE1ydPnNGgsNiIrlJhZFwhAzEehkG
tlkYUxpp9hDJ68RcrvAR0ZDQaYE7oHd03SJA61TUqHO2ajW+AYrbC/C/4IQz9J60
a+lDWLaN13nEVrYh/hE6zDOZCesDrUIESwIryvX2TWlShS9hgRaA+d1Ih02PMHNQ
FzoaSYUheRLB67Prnc4W3atugufXOd7/UxgEgQ8NGMfYv+0BXH1SLroHSfD92YTg
Y8aeBdUANhf/kOWJrPptQ18No2yyH5JvTyoXwsADhrqWM1XkNGlAcek7KYDJ0T7B
cFnSBuep1oIAm65hmE6JfumL1x4wsUNwaKEL6nlPClXJA429IhPsIMNld/CpUpEY
sL8PR0hD032ABDFxkIfQtqgmxVcq2o51TFRAjs/5PKIrpYZrENCCsSoL3l+od+X4
US4CI5ReoGNbUE0TJe0GidjmpLBOiTU034sE4nfVsvAbcfTxdB+FTNHQL6pfbGbR
uifMEmh4g/YNvuEABtf2Z0CAPdPl06QMY2E47GeVzK6rMzpXVqGbAmg8e3loVPRM
F5yNiW0V886HK9MKwr2oDHgvrX7lo3PeQSFN39gBPdIG7/hORn6NBrzsQVyW/852
kSONxeaVOApyYGdqfnny2h5I0HzwpC9q6Kj5laGmsRLc7hutQNEaDp2obLpA5hnI
MBRA0DalYqOp576JL+dlDeLrfIdl8hpAEAPitXuXjROlOLlyBcyJ15N6jxtzH9t3
29P7b155qBeTyM/dUf/Js9iihUoraJshCcC59TmKFP2IgSkVy9z0FUTcI95R/G6a
T/+CBI19e0oJdSFIOlpH/9gH8utj0kWL9qaYGEKCgx9lg5qOJ4AdrhjsZin/6vR8
iB/5mj+fiTv3Z1hhT95J9qPWHF0Pmoq9SfzQj9a098WqdAXxxJtBzR15/BKkc9yd
4Hx1NbnmxIXzXw0cQvq4Sxh8J9Pxh2/TZ619aAaVRDRZ3hGDuwIstSTUM2qwuzBF
cD1X19+0A9qUbUcEkEfn7+hq8bmxc+seyhWdFDM1qVtHp/Xr+eAHiSK51qcqSjLc
SCLGNgVAeks2ByMR0XZUuoQHLr5kIQiWzcqLV/rX8qOUG5pItSHjj6CUOd5ndODB
mOfEE2Q19mLSdT41qphzwrY0EoDQ2iUIBvt9d3HsDh1T3yR0rVbseWQkxPFEwn7+
kKM6UqW6ltRo3s+mMQFEva5tsMFKckW3/YdS4sConYbyJPhJQvvPYzvTdJ1Q89wR
Jqorg2bKOqcm4EF7xZf+gkwpwN7wMVVcke/t2Nhft0ANYt7SrU13vUbauXrqMJIe
952t2jcYq4SIEuVqcS//oLg4P4CSl6vftA3VfaaDOw+tCXsqEjelcPv0d3bOwYQ5
ihkmIuIAufE/lTyurNF8YHvPn3HI0ZGPfXcksdOKCOadUQgGLq7eCLUzi2www60r
MCD4FeIDt+iBreRNINwezjktpOqTxaOxUCHpsHKfR/0yV9n6G1FYM8rVxl7appyF
n2deQTuZwSRT/IRV0CmaTbBRNSNVrkb0hloTKMA4kYioK4aaEA3GU+7aL8SSsAxx
xGmKrF5qmFPeZfpEMmucUgP79t34a9dm7T+k8U/DzeQFfTpWpsAtMmitYCXqy9tb
9HWBXEJLGJ5SAYGxI4uKD2eUUAKGiFQvrV0V61iZvxykGFRUittfWFKgqNFdpE5u
7jgC+aJKxcARGXENZdHb9NVbUnXwAboGoCU7UVRDNwyM8upBc2QQ8rjZPFtpfT1x
YKhJ8QuQ2u1u7vCS1s1VtHGKnxDi9OPPvq9M0EjugNgIJBKxx9CSed/c01+pfgMR
4iIyD1p8ib2XpP6DBpyE/CYW/dsfBlG6moC2hUIbnV/oIRAx1CGa5z/79mAMgRHz
Irfd4hSGZeviJzRtcEXOWiw+s/SCQ/FVytYNq1rLqItiYSL5xvCSHnj0ilfx6sOA
RIB9FkZyjXCyTjrjRD7lCOlINb3PvM8H1HgWNnmhFIYyEyGIc9jXrUFHgRqwglfn
8rY1R2MFEMgppZPZHCL2cUeHlHz93liy8dPFBkeFPQD8/ugfkUDnlg/TMLlZLHS4
mQTL4SLZOVzKFKDyfLhBLQpG3/VIZyI+N4/wJ73PC453iyN8lV8oYzJILAKwADri
HvQPjGrXm/YRROTe/JUYiYTYoeZ9pHPNnGqjjz8UELcKyQF/feST7h7s0cAV7n2H
i0ECKUzfMSpr2j2VXIwWDsateV9sjMBXAKfh1GjO+87svWp2Z69UntsgaMFbDMtL
IWu2foZgFOu5zjS6BJxBSSDdZRYwS4R6eKBLvNhLNgEL4JXh9mxY46iKf9b7PGUZ
njZ1Le/z/h+FpCC8iVL76g3snRiYawuu/QwoYZ7le/SyorygSqv3LSDuPJf04TgY
oRrwRzix9o/UacySbYsKH/jwc5J6MTQ+pKluDmO5gz3m8/guDjN5m74fz4PRe0Q4
Ze4QqsNGL7fIvhbfCH80H9VfrdSA2nhrzvbhhhWhh3DBwXGxzhNpd2X4Kh3Wj99Y
cYpC7y6Dv44mVZF5Za7p+KEKGk+04UZnMBKIO0PeEAHWNvdyfsdCKSg9DRIaHnGT
fJIsIuzJ/ZzY+xlo1BcLRu/S278fstnWfnno43hO8THew0QMJbtHjyzn6HL41Y6E
wmz86JF5bM4sHdSy06vfczwb30QaRqCI+iA9hjpAfYas7Xzjfto1BNy17vozTG31
xiVFMg778Yd7v0ypZk/THxcnj7XA003+FSIc1n2G9iQa+P6byB6Ak/Yko5xXcgyh
XEosCEtiNSE2tsrJ5QGHQId7bWLOYjQ+ic2bn+/kGUb9dlQh7Tjsh2U2gR/AyXak
NqVr4AGYetxigsvXdIgkcRT9T2pxKX5v0QLRRXVK6Kju5i1QWzduWIEMwy/ZSnhp
RRQN3Lu0VlG72tgZGFtwb0WwIziXHkohMuidUfI88qR9AfK6VmvUG3RgUuy5Fs8P
jftII6Q+v7kvsIWA/DeiuwcLc6lxGH++cX7T2269J3x4pgir2wLT5vKjNOykc2v9
iYg/c+/Xz7wZWdouNgBVksrQPl0mwTRFvx3Q4sALAh4idB8VdIv4Pym58jwWR0o4
35dPPIuO1F5HGY98SWbz4dP6keCQm+wVxlDAue92z43a36jYcvcabcjlD0Lr2TN0
MDqcH8EyUlHI5NC3ZK4Y7uZcKdrH99QABrzwYMmXHsgNhjv6f8ZnBuMjIS7c2Pkp
unqSdE7+y4QEjnJuI/7ttNV8+6vFIj5y+wOKyVwiqbyltV7iikibBK3GW9cNx3wF
r36i++S3YcYNCP/Sguue2wCH0QYMWpJEd1vWesalCwA1BM9czmSGFTaWMgLU7QpH
R7Te93Yy5a0LtQz8I4WGx+km6Tl1oy3H4zQz5meZ4KSnp6VPGf+sMRHAf29Y0rWt
uVbFnKxBShsT9iiVENSTCEBWlrpUVL2EBec/3EHbtiJ6CYnFW9hcmXF/YeOgJCUr
ATSuR3K1owgKlDNX0sDqP2bTpqJx5+tzMozEN5N0HRH5Cd19baFeWX4LasKYzNSe
nZW8rXnNQnLT4W1bXfyMA0SRjPiVor+YobQUDRN5IjDB0azF2jmjJjWCE3n7HG1e
O8R+Jv/pTAMhfopDbLtUGnskhA5OBOTwsflb7r4UKE9D18OeaAltTGL7MKM+JUiN
hWPxLEh/Akf82djTXWp+WAgW2WAaXnwyVt9slATpxfct9k0fyG0ZHCvKucECTYX8
ztxJRK2axGTp+66zUxy5Kh6v24+wf+U56MltcgooMZw7DYud7OCekJsYa+8CxVeQ
KUfy3KgF+5lRVCJdcsOJkaBsHazmugSeo1Iw3RtjAIxPBcSKX0xruGHedC17PKa1
WDfQFXyDooAUrujvqcAFx4+BSMMNZ07u+/Fpoh+eAy5taV3QppWjLKoDBMOJ8oXP
xAqZiQJ8bzJ48Uho/cDCt/50t0A6q9tJm7tR+mu+fvPwmLZrxXf4yZyHUzNOYku8
qYORynRPK2iS02zdYkZZQaooDnWz5AIvlTQdT3ik6WSM2le9p3cZg2TvyaMw/G3F
5aA7GUAVrVqPo6GdePWxjehTiuv4P98uKviC/WJlybGBYPOvW85rN32kMxfNsY7P
Gmx4cLgY+4OrLdydE3TjEAHz/GLu1CgWo2qLaOPgFvNlNtoJ0gInDjHiz3LLCzO4
cq9lFnWgBI4gH3ra6R79J7YGoWa/Csgw7WZo1XwKrOwr8RakOF3g2Dr9wjl8/Zmk
0Rm/tPGp6wQ/YOHCuP+gLn+k6MIWB63Q/snNe4YLpqqDAHYscwjutxr79AvZgEdM
JQsVHeozA6ubtXx8hBjyJDm9Z29Wza4pgqSyBvk61aTCyd1Ar2P0m3f2AJm+UoMQ
ey8BxB3Y6EI6NEKK4Te5W5Aqy57nWjbMMvbUYvQJpbe2f2TwaaOM1gfg5WxYm+dB
RmfxDsi+oH/x6Qdblj//RUsgspa2YDcDA3KH50aVn+UZPNsk7VExArKZHCpQOfTh
1eLEaECmAPi6iP6Xfa9gtYpgP23qk77FjGKYpjaOOQIePLM9D/zuuVFM4Ppemrmo
sUVYhwlaeXADNfJWytHljqCU2nPpPGv+zjkC3Q+hEH9zQ5aEC2uxUKm3s1lLBb76
LGA+8Mm5Cfi8NB8t4q4/+6C5AdQ3IvXyU43aaRPfqXcOdqp8vdUnB65e7FMjnwBo
Pi+KsynciEhMSi/6Un8pSn980UCxH5VHEC6AqYpktnrmQyi6OFpa5UY2ilnoKNLb
t/RpeEqNfV6VoxrpkvYJ0lBflFwe58wqWkeDM4H39Y6Rps0L5AOkFzvMfo0pQeyk
ldO/CkQD0G8TAX61Tu9dw1z+8orHawdyKG2wYozWQF9HeFZjVzRA+s9sV2aIOcwS
cVBuMSoPxeHQtPq+w3oaw3RARbwXON9UC0MlcnPqo24Jku/Zw+GOQBmLB9DvX7PG
BonBik800N08q6Qy0MNC2VQ7O0uEHSlrDXt9LzUDcsaHZey5cW4Q4tE0ZVuXW4U4
SXPApxpPhcuYuGRA/8H+13RrLWUjvgMU32s0HyOxd7hc5+a3rJQ+F464pgg1nUqk
TsXcfEhVZoM86HvJN2IO6lo9j/Ubt/yVXJF0x54xzBDqKhBRKH+WC0kLiH0vK9kl
JhBlpFG+apzwYHDyei2OuWd6g2jZ1R2pUvPCoHCfKb9LUEfymUyRrc09akDCNdwY
+kDmtpxVFZQGuu46L9blIAHqPUcytb6RlaPQJgMSEjHXhg8iWxPhuC2tyVRiznqz
SOpfvdNOwaSNO+ZglHjJ6/7OsY9xFLI2/rVkZic41yyS1FifGJj/O2J6/xX0Rfdz
UHcY2FLO4w42ll2hIgGd6W/DDl74N2Fgl1dqUtGFMTtRtA8fuZ5tMxl540rXV68Y
+YWaf76UlcIH53PIXKMPN2rXomtZsdh9Lu/3vPffROZ6nch1oouTQIcmRR1roftg
rNGQ/v5Zjs331Q1jPVGlrCaLTw/Ils1QOwYv+a77W6r1z5gFHgn6uW6tm10ttAIG
LwxGddco+wQzyeWSNU3M2nUZZIm2DB20VWZ3OtX5zt3xTThzgUbXIuSS+ImIZ3rv
ZQsc5u65ns6VS9f01R9CJ6eUu5YEYyKdTq8FYrzvZwuqFGsxjPkxFtOA42ILx0cz
4oHI2pXH8N57qFN+k8fc5sim6y/kMKg2G/kgpUaKI+pExC5wt7jjUWIHEDWTDi1t
EjY6r5BoF/j82iT6ZRuPYv84bUe6AP2YK+O/cfDOqHYuGxIK9XNoq22HfomC+LkB
35cDjmkCF0lc7pTKJYFrM0UEMywpJhgrB5LDoyfsPlQS0JDBEREuvYo0AVnItT/F
7RZb4B136sVoH4E7ChgL6vaP80WwEMzXMNxobyRVwHReXu1hJUFZ8O/ekKI5meP6
/C7EJJQDJQTsyrPJn3y4c+ktcJ+phsUUkBKjiyaBjrD1wfQcdykEEFzFRDlrEQU2
ew12xAFDuBdGKB4bWF6rCyOvAsJKQgNdRz0XkAE5TZlbIkPBjBfyP7nG9+IqLAkM
eLL4+6rNEnehfAqN1CeMLBODGeReJTiqkOIes0TSei+qqSLCEVq1OTHBRmKR1u/s
aNTMasiaplZGhdcn/pv9/EfFLtoXG/Svdmm4EMNEdW2ysx4FTAcNVeKvKyN9fitJ
511HFqeC4/GRXK5kC7nfDiP1Cyv2j98q2SO2/mwvcvd5qd8xPIssJtm/bPCBANg+
LXqr0N8qlXeg4SoPWL76jnplVdFVp78UYMjWC2bcvnbX/5YvvLLpdtjShpY1+jIt
WttjUSIQtuPnGv8uM7AnQnBGQ7iLpj2aPxg8y4/EYPbGUutBHbXKst9UabtxS0lU
8gpS0c9WA49uOljcSCiIE0Jo7j/YIr/GoUsh0dZDzJDNCggrjkDF9+4br/GXCc5R
RwnWx2/EQm6YQ2p0yacjsRPke00fcSDxNRdbkMVSGel+Pf3LDNa+cOpKwRPvltJW
7uWNciZScrSW0fABpXX1SenSFDLxzP3B0i+BOyaQDvm7Rwp4h/5qRpw/d1TtkpGY
tyJAyAWYBDnRAHR4hDEdoYRaDZRNmNlms8CNLJ41zd2Ol40FtSa6AnB9VB8V6WU9
RcFNWmcr5n4dJQK5aX5VABwfmSFuS5jal96InM/pI38/MbY1X9LJ1kqh/GWmOlHv
kxC/4dWq7Rw6sGOri52g7wdVwI6Sf8fl4UkQSsbqmXvweKIc13oUkbAKfD13v0EG
JH1tY46CMJeFJKYCEjYQKos6NJIhlcCEDClt5xGmtNM65gwcIjp6Pa97BipMCBvB
9INbDi4AzdT6+tq34Plgv3be3v+kd6eOQ8v/Goy7upqSU7ghO335UyB12WaX/2P5
xia+L/zI2CvEhuMDM9BcdOq/uIXN7Q1jy+obY5Fek3LnTAryemjR/3d7Jz61dLpO
Xgq9XYG7yalytpDHAIJLZy11V6Np7mZs416Eo48rHN2UiFM7A1p+vTlgdSdu8ejc
UDg1db89bm8fIzqRz3XcYIXH9wtakQ0X7e464cgDPg0tEzY5PZ+GfkSX7cB5b64/
PYyh28hGqkhU6gB20znVjKHIieD38Jdf1XL8r1J1Fpbr9GrIGbZrCNdR6xigGBny
JehkTp+ALNnNpshPzGyYfuf+5j0iT32YBZCPSCEnT23RxDm0M/di8EfhB7drETEw
4dIxztbnTWWbdSm11Z8m0O9MHNEEYbwO+aSJqbIlOOE+9EjzfpHTPmUC/o+x+zZi
XqDHHsNRPIftHjgCQ+K1Hv28C1b6HJxaAQbAKFasPjY8dTvaxxWQUvu1STTRkkwy
MxZ4o9veLQ4eOG5exYiT8v66IUDLt42op7XYbjC9kdh+4pIxjX7TlWvy9HtYzb4H
p9T/sFDdlLSGoB+PNfwXcNwo9YcwoH/CpLkZccgDObgLxtFu1rDnKtbQNCN0PC8L
lug6ZeuIkyeoF6TnJVPUA3AZhivt/yz0DUNfvr8f6euA2+uLby7HH2L7reenDEKk
iueGx4G/NfteGH76iQtQRA3Vdv3eLpOId8WWiHjo3oW7D8FFzhQTBRzQUde5oT2G
+QhtDy7E5jMYCQ9AC8/oappgX/TuCiAO70U7b1Q0PLSsFyLPm21KWh10vq1nOLtV
yULC28U0IbmEzzSwFBPYvOZ2zBv3SCJmX8gmVHbBrHi0Jd7R/A4nXH99u0TwUPX4
a73swK1j8cxw9yLgnEHNYUiULKZhYnsRLBWXgWdY3GGqbppySZ7RPwYww9bbcazq
noMLUIOTn8FWKFe/1np5tn/LJxQ0VKv1zhYhvRX9YzX9+xvMQ222EE/DzaamgPB7
x4us3m4hF6shPIip6JIuLHhKPz9HXCRHERmwox3m4FIkhPOCxjUqjJ0hzmlECiFf
ONQkAunFVJqpyFYpLDDjvgtzhoCl/T3toBeKJnbzYtU8L7Uy05bi8CFLu3oHU6iT
8fXFkZuF6efPsa68cH8d3Ci2tQ0KaNeLcELEphdw6igbf8EpMAA2BhEC+PF0jHuV
9Leje3iVaLM1Hqs1tbAX2Gc0ivdHjpGPkCw6vGhxLnqTELJCPK/J94neTwxCGT2b
spS0ZJrPthUxk5q0cfbWnZvESYRSQRFFEdireiot7JIiGtDC7RdJo5Mwk1VYTUjO
fi460Xanc3J+LxoZPBxAslQTFI93NUImorPch2erApnj+Cs82lYtqYNE4BhJ5UJq
8GzO6Zg2JnZMF5bxWVm9tVkZvFK5DlyIg72KKoDUJ+IokmtlgfI9xpu7rb508DZO
5x43teE+GgVIgZ4NTXmdOswuZQ2T8cDUFlSsWdZXWvDHl9DxqP92e3UTlrDB0/i0
i6hwnmISesNVi1Lzb6SC+LAby6bt1TaZ0xML+sGZ3R8kp5O98Qvxi5TreW//ZaHW
Kx2GsBjM77d/0SLVH5oEb7QK/UICdjSdPt3d46FSnqnmPLtvj8RV2PPvhgheoWjs
ChxJgXMjo9pF3aduEllKFN6ijiIv4sWZi33/HuSpT+J5EB/HZab1FiaTr9pdAiDG
Wylplivf+OP7BuK4VTkohmeMB8Tw0/Rtlv97WoemLICefSFK6e1Z7YXKOX+6AaEB
vt33ztix+BiUQl+qShkA5pUNyLqgajQfhCpGZjnbUjwz5kBrTpuHeYStluEm71FZ
dB1OeixXzqsi7D5QgEDMKGKHmBLI+UHwhzSJliwnJQmXBf25rNm9bXBVa35o81w9
43plxtZNl1MVxywLvADKSGJtxZsCjUbx7jBElBjaeb2M7ZaoHkezvcQ2+7kXFQJ/
dlQKXRiYkJcezf6vnmqVF92jhJO5ht2p6NgTV7IuOtz4eZ6oQrcR0jvCjC5EPFaZ
EWKmb2duafI4tp2XPFXvJsDLb2OHvP/eWkLt5YeXa7laFN01qXqFNXwvvOYH71EB
xuSVZYXMcb46KGmMQ1I7SIkHaZg03I2Iz/Xqe+QeTFlETtxSzEvS+a62P3sYuBQP
BwTIMpQAuhG+Oo6TbGQzUQAelekwlHrhgWRBs4ZXHvZco1cch7MLTtW7dgkkgRWK
X+RoUoMRoYlQsyY/0j8d4D7ZPWpg0F52vuJ5sy6y0nrIFcM2O7YisD1s/p4p3T4w
No6gHxvycmMOpAnJLLG3ZZ+mwXQlFuSwldFrRw/KvUxE1KQSK78JDpBwXxcXTvSV
7LeN6C6i5fwS3LrQkRdE+dOnIERpUjSdFvmrGuuOgTG7f77P72fqWemRWzlw0mGD
RwpYwbBLr9vctT4XRwfvwNJrlJcA28nx6nJDz8uDruGp4W9GsoFEdQ8FDIKr1Isw
5XUwAKqNe5bQcdHyazQybrarfZmlDl6WAaZpYzOIE9RhDbv9632NxS32zq9do9I+
9W15c6Eed/K1oQAzYHpSjyqNpxzhB6FKq27xvmdlDVJ4S6ygIM1/+myivESG9yYU
R5k/lapZ9cYKYAzLvVz+bocn/H6MvMOJZc7l01P28XqmlpGuG/6pcBYGZ1RKKbsn
AYBGSauZomsqUqOFcCBMKshXsKYo/mYFkKNA4Cg+As2NI6J/6qmuBqqm+nbxAd7C
ouuNLE2EwuuXkwu+DvDdO0MeZpN0x2V2G60d6ERm4eJeUyy8VXDjEHQ60XpGZzFS
UAubOK4Fu2Z07wDqrASDN9PY8tpBFs1LPEaDQSs/hF/uPbmrAXtTOwKtsC4XhWam
ZaPJfKCEPiRszReG9Z6Xs9PDG8f4HjdRWGVI929klLNepHv6+7z7TRQAhFu5s3k6
okAm67/t7AEtLygQeOByYp96i0rQKwjXV1tf39txbmNMrGy6jXF/++uz7HTSM7RT
9ke+G1l8DJ7rlLxBOA6PM79W0bkwr513UDnIqPYemeXmE3NswzRr6xzrG1H7eL8t
Y53vNwfBfMbNixIXmLeHU0m6XgKINOTkp5wvqzhrJCK81UFI/WmwU6w55b/Aqy5b
YYGIUroSvkLSI7p3wYMRd14uFMMuz2mc/wUW4YcZUcNsZfGZ2MPedmzRcGl+ywTJ
xyNQZSMNGMzBL8Zad1h5mz71MBetJIkNx5H4C9zG+AIZFxMc9Mwbb0ZGguzBk71x
acWncfebE593ScsvoL6f9vSfnCHc9/F/LLKavyoNFPQzpAEFZ1RHrKBLCfudTrdW
OIOukRa0mO8g8bQZaoOPpGpYwxIKjSCU0fZPRhHO9T6WicOVvgUaruEgX7yzIYnb
lZbDmVu/L/YUBxHUfhcnvJrhcgbzMrAHXY4HIUSJt6D9vJbGYwzTa2r4hhxXbmpc
EEvi3ugsR9C0uqtejYmz8LPftFFKE6dZTrcK1fntUknMLLS9+YIZ2biEboiqdkV3
B/PUKD1FAtuK836ZuDkSBwPyjVEaYJxWvbPLrEOzrDVpRhj5O8Ezrt+bt9JduduS
/eNkwIQey9Z0AErhfbDczYWtr1yBsN0fzyalwL60oZHIeYeXWVTgJLRc1CEj+U2i
g/r/75NuGPSuleCi2xP3ErL+KmKd6jAYtsGndUtxFy51WvQew6TzgP0xFV5BsMqO
kBzUJT9cUW3nyexJ8vYsVRKsg5KEPGVPUgmdWo+XTzfKG2wjovWRmkdODGk9Ly7o
8hx4HcCKRrx+eJtnB4IdLqGNdT12JWoChIY6QfkA7UmnjBHc71NWqzGpco833XUP
8RICzCHf362ci3BRLU0brU1qlUVdPnsgK7Rrm7h3ooeUxfLMJOi8JZGxXgfuyF9S
aa3Dmh5VyDQ3t+EDgsV5TheDYfjBX1+1vRC8qqpvlZ20W9tJ2ygqUcjZvvN2Q/9C
oVJasED8mT7Jh3KrjW0KMXyvSSDcyY+l0eNlVGkmjRQfqmMFT2ySSfPoNLJMSYl5
VwAsF8KLE4GvkFZ8xO4nd94KIGBY3a9BL9cZcov9OmgwIKhacqQC8U0ZhdT2jqp7
QoeCiyhZwXoJ1x1w+X4BjXZ6mzSpXk5haz9zugZFC1DobrfxfGJltCxP90TQ1h1d
7acJvAx6oQGwX/x8KHb+ZULKLg+3NkPZZ9czX0Vmmv5KRnsS1h7mSqJ94jWbSSqO
6zdAIrsbl6nm1Pn8eUXBljDkrWnsFNN7tPBQ2oWDhioLnIDkpdAS8iORN3dRLSPt
bf++PXpgxmQS46I85CmppAIR7cgeoTFkcbcBy93sfw6YZcqZxWDuNMgz+jf06nuM
rf3spyENq3UpuAfI/jwuey/17dwanH71JcHEUnDnaDkRc41/rg39rogn+TFJnhRz
/c6omkUaalYthy+KKT1GxQn57r2026OhV10Em5N0jxqhSDiTojGHymdq0emvWIj6
KdbS4kRvV65MkZYgLSyakxemZ0iJvPzqKqyGC6ZXghtXF+maCXmmW72ocWU0f57s
FvnuHwmL1quhT6M/KPpswFYU3lxOiOAQqqi/MTnCwi/yI0n3nOtQc5dfyecawzW7
AdI9Etp7TiQ9dB/V+xZ/YCWrW5SzgQC20a6XhLxctgJ7f2klnAV2l33e5s4tui+2
I0KFFbWGkwOuOm66HpeXJqAvj93ch3XCvrc14lUAx83TZn0VMYkSLY7DwOmjM61L
+dcXNX4CRUQm8q+zYS0h3mGrHzkY8CrIls8y0UCgljmSYtj/GaMT3Ln11E2hHNB8
0haIvP+Eolds+t21q3sBOVWkVOBM56oenpjhTD8mCd98zwBoKi7ZZQiV4xSITwT6
5kN29bTv8Gcejd3iiyJ4EFxqd/6R7v2Ba3JkjloNDhfLJZkWKSDE7LU25YYtnUd2
PIxVoBaVsSyQ7tONlHH/JRuDhDPXQ2255gY1v1C0I/ko/aY7cRgd2bXKD3u6Vavu
MJ+Wbs2W8Vxb+BwVZ4ZlIWdZrFO9Hn23w+NjBORYPkDQ3Qr9Dmi/bgLG0K6BAFLH
SncSFgx8ETDvgUg7zXVvtIIrWp+abhbLMiEQB7ZZJ43xKGQkrTTsOn1qcVr0u7Hl
UbF3JrDn7PlsgIMnUOR+TLPivhX2T45ncMsjFVkS7J7o9GL8rEeMiDxuoVjKK2rB
YFwBeBCxjjzC+5eQvP7rcY0w6YAkliYin3ooTqjejw136Kc3QPPY4w+nmPXquoq/
nof0K0JBHDKMR0ylcIfPrUI4hhc7qtGGvi2SBT6/P+gNCfFHgGFx00GhtkNB01yi
2wrsmk4vXKjWqRQqN/H/RkP+KN5TBTrJh7rENKlwyC/yu6ULBAPL+s+YvTZ4KWXW
XAS+GP/qQ58xTynFk5Q8JLugRVkNCj2BL5JcikyDYGyxqpk1VAIx0yptC0UUFW/9
HLwwjT/uaK7CSmBCTh/Ib9fzONTBRszc9U4ydyF//N6gXZBUua1Z9Dtq2tcCRAtY
yGlI22k9F8byIjZDUKUvS2KAl6oR6J1MXKSvL6alkFQsaQd6ZZ/yYqBA15eOpMRN
DsbLKB3Kv/OqVmsrgq/wczJEJ0zj5ktPX6FXX+bWjM70EIGOZxL+sOoRJd6esla3
to3vM7XSYCpEvc69sN8OCBciWA6JNGpDHJokdV74OMZNo4kCX5BR9aC5eBHvxp+t
SwweDFHNernY0PJlDShRjkCHq4FvGg+7GoRfFmbUDGKkSLS7WG6ePoXafRSBq8SP
PLqpAOqEn/mcdQdc+xuFUY2x7h5+ZOqo5SZtnroBg9+SfQEP8dL/WK0RSQiuUPr1
t1naOOsKNWr0fQnBOznUcei3AbWrdWQjMQl2kbhTve324ffJh1+i99WqWdEYYrGf
I45ZAAO18lHnqSEDhumMNd5wPcUvyvnFos987/bxGPPfCSaz/cTfYfKNMwyuVYMw
dR8k52g5IFABM6wW6Tpoq3M4OxWztoQrUBUtQb6g98pMmh7OzAPEd4A37lKtVRKi
nQR5MlM+8OOKCNapBO5TsSsiFDHC9uiBfyuMLBrx/2pmyn+3NuyR1iu8VJnwu6YZ
zllJOKmGrsn5CL/t5fmbzag+t89a2PM6mQgOaQEU+1u01hOK4UdzwAqEilbnec5g
HbH9U5ZqiJct5VIfr/0Ymijn3HafcVYvwMEHNK1uvbn3d8wIY2W2/LXbpde627pP
y9XrZZFPujRYNfisOxyl3TGB4d2ck8iEz5gGhwLol0v+D0pMDic87iOlQnHrwpnc
afetQopBhy9tF+C/73Qv5ZAv/wY6zGw588UEhqfCyg/8jpr+c+1e6P4SGo65ATyj
H4nmA+o6+u0y8R3fMpPP223I6ralgaLArC4AeMuMh1vzGP6TRKMMycrlmcvLd4aE
ikSSyxeQTwFOjXKYHibQftro0SN547b5yBs6J7yC0wfVLD+5JDgR9SHZAfbZXKGg
flwV3ONTZP7sTEtb72QHIDXRsxY5XA0pzLaUIfFd97oWjR0N3ZtAgm/y8wE0mYws
MX4FXDBrDr52krg0OyS70/tLjM+gv4dPxyXtbQPpJZ4/wpKLfpCecFHGIE4Aeamg
3joWlch0khiv6Vm0ONjau8HJhr9gfrQjAqVzzUocmvLmys4Mr9+j4uJ28lghgs62
t9WHBUFPnwb23G82Y+nqWRoi6l/4Zm4a70s3stFpxOGauKP8KP5I+S19tsmvXcs4
Hd1d2FIim7VpYcXMsnClFLHvy0hKOq7srrdsBOlOX4rww65IsupnwtSmxTk3jL9r
1MEd9tKmXTCPIW0L/cwdiNXfAMjsbya+QsiZrFltckZ3JuWAb+QacUM8xcm6tgdS
HO+aSHunX1sExm7+e+XljBO8bQ90jtB+kVfCcnXdiuBwdFfrdO5v5Gn9W+dQOF02
2eG78WUbjWZ8Qj+memqMYCWpm0kzGOUwZL2mgWaBNtQLqN7f0gCvX24BPatxb5RY
nhA9KEzrKCkCU1OTXZ2lOXi/uCr27IT1ii1rK2fws0Pa4BH+xELVkdMNMxsPz14C
C88jqAFSLM7xr6wh5SJ+SzoZqD9IagFUfpsY0M+oIR5JpZV+VMREO/P5gOZvJWco
ZDWo6WBqbU2pDcOxBAvru7KDhyfQDuyrODc+5R5sbB2vliadcine+AFB1dKr+ZEF
tJrXg6MzFmlV0e73qnzr6wQymLKy2Xiqqsx6IQudkn61jus3trCcxcd3g2EBPZkJ
GUvGTjtqm02JmrIk3rWdYCW0kXkIBIckdsrJovvsWt9RUoyds8qk0pIFcr+nKEwc
F2vp8PO3nrTnVmHX71QFn8o/vQ5PFkxCF2bFapBHFBxSoIaCxKLI1XwUmoPsHO8x
WEaRG6BR6uCQJbYR3lQnbiCL9LWfIWJgfbyHOq4qKTS9Z/pI/39EzoB05WFeTPOG
tOL4MeKV+e7LRxFqgHo4j+cp3g0Dxz8LgfOsFZTHFzMZmj8DIlFZwx4dYTgj5iOK
xP2cwrD6AYfq0hRMgvTRXyiYS2Qb0VGPywLsTu+FktZYSL35ugucFkoG4BCUy6lD
zwWlty3y+sUvYkziMLZ6NQztEainRNl3dQce+sAQHEzvgMkfUHbR2U3afT16n6JS
HaCRa720avQJU1eypot62sjr/5VRS7oeKXo2AYF8uQp+i1JP9pmDcRFRNg+plXkB
r4Y2Eekx7IXH99zUmtTyGWOxGipglpcucksByQlfBozOSJ02XQWIo2lHPvhbg4kL
LVYH1GedrLEvxPY3E4OQfatl0AwgXtNL0kMyFfMHUv0lpCxYtRXtxcFxfpLxljgq
AWztEf7Wb9LqymbmQJUKC2vBdxblejkUlhQVLbg5aY5fPEUOqVEU8bxvu0mgPBAg
cl/zkrY2KMSW/yrCX+7es0cxKZMqzmTjup3rY5x6EpM/xqQZuAJhEph5Wf8dfrZq
L+po/V1gKCh1/MqSa6a8MajhbGFurwz8t8kbfUz+Cie4cahhGkRwmDvwPAxS/+Ar
6Kq1ME8fbi1p3Ip1JCKs8XNM25qwnyMv1IXwB2Ufbf6KEcjaM5hy5Jn4TzJdZj5F
NIJmaQPAw0Roa3Gf1hJw1l4zKRUysH+ixb7r9DGXB/PPcAbvxEO2Cn7h9bFEQNeo
/qKfcq/0efit8ztkSvx4nAe76bxgpu+zHYdR8rx2G5l1B0tlDrXKUVNmNT8gpIgo
LhwFiarj/7b39D4X+rDOJOK4v9EwUQWjfpqQf6eCTbsDugPvJJrB7rsgnZtZWUY/
EkZvMXr8tZF/4r3y/rJcPYykf8WmcSVHmbydgVFaitlVglCJZRMCROHajHCRoYjC
Fm8aV+bqGPjPRgPSLM3F2J6ZFmMlt3Ae8GVnvHv8/2VZkBrAvoF6sJ6DwsYjCfgQ
6VWD/btGHrnnt4s/d4it8hCO76L7MpS5J48mWfv2N+isTCKP58WdoP78qHs6a0Cd
Fo7d2P/C3W8mwX8Vvha8daB2nas5SfV1eAyWovBZGh+dHReeSYgxMD7PH1kcySon
JxUycPQVCZZmXH+sYppvCqtHLMV/cKRL3etVQsTk0C7+yzS74uQXkAfZus8pJEV7
lXbMRVgP6M4nRRWr78gBjH3pbFfvEnz0XhIMi7+NuktjERE6SjdGmK5hfpv55SMh
hiXiNQRM1dAQuOj6BZUxPc6f4k4d6JcQDBnETn1Gj1PA9Jc9gDp1nXVOi9tCUMgy
SdMid60xWpz3SWdWElnA1KWXREUh/aF2yq4TwnAQ2u7qN158dsbHuBZBmEl1z6O8
+iTt0TInnmZdBpEmt+oAz+vtnBfoXWr8JSo0vx/oIq8CXEgZRytYo5QQKWULo83g
7OVyvQxnfK0eKuCREJw1g55+enQ/YbkNGI4MK6gzjtwsyZHGelxZmkEmwLvw+KEB
N5YoxkXB63/d4FXQKtaZihbIJUDBrL3W9Lro5d6l7k9gHas9O79TLoMCDZ6hji8A
nMaXaefGB2/zc6jU51QncHDfEgYlZuIrNA716Xv3iveVXhMNdfxCllnhpToSiFld
iR1+1FkM/BQAw6J6REuwZ3oL5scYPSxhPHPyN0/c1VW322wOGuEuBwDT14R460bY
pPRL2Anj1xxymZ2zOIrCfKOgIG9rtArazAaNAOwgGH4iFOx6bDTyfnX3euXOmEHR
agJPemRB+8Go71q8JKhlzLco5hY3lCf80nwhFoykBtvYy9q6WM3eY61DqqNhzYy6
cEDMsHJUfccpvTcTAJakSWK+alpSkVgIFWV/YiRu2wwBMVCKNGL3dwg3L9YdQpA6
JAKKUgSbA+zRAJjebScgppRQ9N7Q/+V0cu7fJcFdO+lNQViUVB+sJZAqj65JHkkE
u9d2hYGuxS0JFsJ469TJLPXqqFm6Y5SRjSinHTTJsO3hoeHHMnTJcqgG3HQ3DJHv
EYn7NZwGZPGXF6o05BtjNQBIn4paRDi15pFtKpDvk6ydvneyRfsmm0f/cmfk+yDy
DIEt3USbhPYgFB8W2xCeLw0e4j6t7jDuNG/2PAvl2I1eNVJHDiMfWiiZV+QuPagW
SFh3N5U74E8V1tV/UraxohJP6oOCmrU2VDh9tnoEdWmh9DRENz3Gat12npWGjM+x
bJpzwK7IwMaVHzWJmhwPkDMZKwIgKad/N3hndJoSk7Eqq4FGxAyNCvjMJSx+kLQY
HT0LfWtr0RQ8EGeKK0twauYmVJN6j3yhqb14QgAIMmFQrDe7nS9vrie+9P/irGuY
bjCa377jgbAhdtShT2TI62WBhQH8V3vWBxnX8lrR32ffDRBO4RZTPCyFVBYmQIN8
HwtPwy9FZdOnm6A4NrGF1kzpO3lV21bZBPFOc+31pcL+Gn/z0K/zHqqjpTgPw4q1
P7tWIeUpABs+viFZenA3JdEThjXO5xGf4Cmi/GBJlZJcL8cPcB3cxk5g6tcI4GK9
nCAGcWjUoob9a1C2aWYea5htuI+xggQAdre/p5ut70ii/Rpkdw7u8wkHMXqGorwp
HRMEhg0a0cjVpxIiS38iNnwvmSRTlw4aHB7O/GdXclQUw3cFkmqmDJbzotFBhSZc
qQr+TQVDxED1d8MBPpI8iiZt596psdW/VFviD4/IUvcTfeYdr5Yt66Qt5tSyi3ZW
OrGAiXs1xSxmmEr5T4WX0nAp2gOBc3Wn2NjEbBUd9LV4SX0/iNZuER9AgLqWo86w
p6aIQXcfWVBNDHbg4bkQt+dbVCYa0Rv5/5l4zSB6oYvB+TAvUDB64tQ9JsvS3QDP
wn9FwhiQZVU7lHGjs0BmTbwt7z2NZK2NC+GL/RwFAidhgJ2kJ8JtpC5KDgam8/yj
UfJfnlaIWUWQaa8mEkYWblEMFy/0cozW+iyU4KuZictJTtlUlU3JK3nVHURb21to
IZI4L6q110BmK3PDut5jp3o//fQ3i2TxsfE8onYCNeb6UskuLjY8Xecd+ioYZzur
R8Gd7/ix5KyDJncc/ACDxsbhOvaBgjNf2kuWM2R+dtAwrhhlq6us09isNeHs4+/0
wRI8ML4VcTX3AkzUgjBSJAA+dx37tv/q/TZ5ieeoRrzqHACBV04+iNT4cLMmIple
8sHDCaQ1A3RRhoRyuhhAKZGHE1AxTbz0Q8SyO66lOf6aEsUlooEXfvy2wQG1xjhl
f7XM4ZgbQGq9m3TgqtfbehGzI+oZvXT8yomKQUTmpWmpD3+JXXxuJa5sn20AfzYb
s8cBAH+hUO8S8k7yfDVrBfgUDuMGnLzu/0nutICfsGbHBTBjqxfEvhCvHxu7FvKz
kXbKDtEKLz1hdNhWX61BH6VBVWlAkDKRoOrpCPeUk7u8LmNXJOT7R5ENYLRDCB8s
CiPGlpsQY+XPbRZZLe3ylfs/ImlHXh2oWbyYAFAKPObGWF9iaBv1ym9zQw3Odo1l
ehCtf9XNMjqf+J0/3Q8OcZs771TLPWb/+evZ1hnwdZZm1dHhTLVudW9ClE7VoJ0k
bY+aoZdp7Sgd6ik/S6kAR5fsm5r3M04fLIjilUN+DpN22da9jJJndRjtgL9lzR7s
XftHg88rBkHT5Cj0EvAB4CO9J43fm3crmDoPJ6Y7tOjWu+VNLYcVsiICEUTLBizd
f6quQR4X5UJH2DmdGWR9VukLV9t6yD08BB5fbDQIkhOrobeY+v7V4ujdmvYaeMA1
BJqLCrg4gIMG1cKzMCUJbW7cE+Rf3HVRljUBzoA2q4NWrTsIzPy0NcxjOIU/kYTM
iFIxAkCdFb3XUFj8dOqrLEOBvkTiyEgh8CJxHb54ZmyCHBQBJawKlG2AOWfml1iS
BNsp8f5BgZU8fdm9SSne7Z14AmEFVc+fZoMBkNhcZCbqjRp76IOrXU+wFPdzULXp
PLvFZ5NyiA9NBwdHw4do+yPhZk/zfNqSO6N9T9fRQlbtIVFCwh+cRxSuxFitSVpi
+Qsion9WLW13/6G1I60n9874M9DdJQNKc4zsa+ApmXryQJAWhxotC1gWkROANW9L
azsw89CNzegAnnWi4pvGBt6DonKIYU71mx7m2m1hn5AdkaFqzGBnpc+9BQzmEKul
M55KJRrDdUrHXiGM4kmAHPnPHL/SfjSaTNWieiOcVxJlR7SocoHTBCDOQETgSzWf
jnjhAd6dJsWdlvWLOFDmhAPgjLyzGdGofPTa7GBhjT/2Oy+O2kRlwhKFx8miapkb
NVibLIkh03nKLZinL5AU6QfZcLv87qMYuw+9FtBWRVHQbcBBbUKn0uin2aDPCZ/4
oDk36hJaVoqNq+obdiSqEvK1u3vSoiRyws6696tpZ2jFteb2U+mF8yY55s0r8tAK
rhV9Nbv0RqKRtcSZMR+XgQxLPlF/shfBYGhRUrQD+vqHHCOy8rZxejV4Q0vTzqAu
osOEXeMk9nCq98biWuWDITMp4pLIJKc4f8qNaDrkwD5TEBzJR5qabo9q9tj520QS
MWjRy8buGXr4tc+feVvmuNSrOKbQ3QQ0qUVmWqxduh0vJKh0tHusMqnk4d5nQpPa
WMtC1YxtmZ0/nDHvnhzwECY70xf6reQTiWnlIj0M8Iav7DxyypfytfVvW3YQlAZW
EvNN6v6clFAIH7g4T9MYsSuk4SfuNZW/o5xzzhbzIA1nWI7doK0mT7F0smBfoJlI
vabxIblXnSUViGkZ7tky0M+pSd4MyzFKmgK6rP8yb2y0oMS51LLy+5gkgMaqLo4z
p4NMNgASZY9ggTh0ztitIZ9IumylxFTZNx/Rv9B4A7FaRU5XbVRa5GYCQRf8fSyu
8G9O0TRcRO2QfNfT+tiZVKwJLDRuvGjwtfc73itC7uHGrEMTKbT6sqtSzYqv/eBa
BRQ08IvFmqkqqGYqO5OTtq19FpT05uEH6AhD9wSMffXyV9rWOWmmALuY3BgEJDEc
dvO+hdDOqKaymPn5FAqXd1/CL/n7uKAquB7/gFoNEvDopyloKTD+sNBEPNE9BC+Y
cURHz5q4pxz2rd/2FslHTWcFBJy9xpAjdxocf/DDAkfgrFSz8vfY1xNlyFjX9G9m
UeSPP/0b+ymY4SvW1OGigZJNzk9f6dEJ2zfHDA1jW4xElrm93DWyhK03kMZX6tdv
jpNKmKnozgseoHSRMPX3X+ZDRYlVI37QRdKzdLNovMJnuraIU2o3guvoAsxxNUzw
doXyum7/lTWkl78Z10Kwupt48c1h+5J1ammPFg9L7StSHJxy+WA1PHJgGGy5opOZ
Fp3eINBybRb3WXud+AhWxXABc0tnY3PitxWlViXf1mIYPtlikLWDHnDxgZrrOw7m
jJVzG6MbdQZQnco1AgUAxiLAbfQ/kSPtZ3Gb1owxa/oW4IX+noYz3qWA6fbdu/ds
5ZcCZvkdtLGtOvfARzPbCL2b9jFOcXHdLj7BcI7xRr2Qrbhx1vn8Khql1yxzrClf
siDE/ezA8qu3JyBoB91IJdAV3FmwYl88VS93rgbJ0eIHM9mxkveOjCfoVBuHPS1g
BxelSvMnhGiCgRaXiz/w4+iiGw9dMWuk0fyEyNWFB2rtr9orKryLTrVe2c6zkCmS
yYGlXJ0sL+YwRfcAVpaJ8PV9Xdm7FcB0/BCWNMjFFg2970fQ8Bhsd7kxJf9Z+AlC
pdvr5+MeOSHSbk28SY9W8+mPqNdMU4nsDRRL1MvpX6aB4OsxSxPbODW5a7IWoZCm
nT6TwhMqwQWTxfBcboi5WyCb1PYJpvwZv9OH/VE7X6KF3dHfIycz9SyVhtEVAkXU
4I8kFOTWgQFisVwnh/JMR+aECjJ3O6BU7B7pajRcickSjE3AWAN7HS/gEKHMohQe
3XwWwKEAFwHJzHh/423xldXD25+mZw18PshIlI9FBJQOidUPyaDZmijF/ENvQCbN
GDgc6nNF+KSqcIXKW+nxTEaanHhlxLfduobxy3AKsShgRBaUQuZl+NblfJ59pjAr
trxnNfpu9RQvbDu/R+3cJdDT5jlAfUxSpbHjKmDKNlQMxZf1CCtjgykBJzS3LBtO
WIX+Qsu2sN5fXBFMj4QV8crWn9q+GlpwTXAOFHSYIPQxnGARGoEuSW0mdJ4pZiPu
Ndipaj+iAj6CzFH2sAxvVpcLXNWm+iZNI10JPWxEyXbxkCtSVEceOoAmxAzHdo3G
UpB6A4oywj/q4zsTucwwWqtRWG4L78e6HbJHt1lTWkv3/IDXr1YUyX5hHx/8VCEA
UoE3ekJviPFUV8HUEIXtoFDm/x4awjzAs6AByiIFHxi8wOk8BQWxbWI1XcxvZhPG
oATvQM52RmoMniddgreshV3vkwh/0QwuR2Bq/Dd3aLSF6ZcBlampy0tHPvA88qtC
PnIXk9a2MQkPdbtJDenGZE+c2HKM9HKxHaiIcuMLZXYjCELNzzAp9H64uvKu1yXw
b7a0x3Sw5/8gofcT4INwGy8pavRJaNLZ5WiYkaNoy/owU/pH4LMdreQqVDQkD4aT
98aiP1mKgaeKnXpqwL3HX6uBfWjPme22J0rYXJVrOqNOIza7PSTD2VvtWO5aizNs
HoYxw13l1K0A+Wkr+YrRfh5bl0tMwdM8Pun4DQO+Ryb2Y2NjP1lBUVJl3QcQ7nYk
EFwOMWBDK0RQK7waemaBXPKjdP52ZVoIcjgaxo09LIEZ8bfac2cO7asoXFG56WnH
iX9tTXoxcISkxboG2lOxSYAe6lklHnaqIRmXxV1a/L3RfeKcrIR5EY3a9Y+Yq2C2
p8g1YRootKE8zF3vSOHRAwLHAkHQtu1dspUISU1N0o+e5spvlpBJFXKqbWKmiO1u
sj75FPIzB/ExbN8bZS7DeBQUoB0p5nAA2QTOus7C5xIk4KnmgusfQq7gxTYOR2a9
PgRD08SZ5p0xlZKHoyzh3j7CP6HqPXcNnMHBy6ppaWxXZE+3N8g5B+wS56/9yfNg
OiVaqB7EjuXxwuA4VIHfL0MffrgEYPN4hxeqlfA7kYA/OAQFEL5WZUtK1wk17NEq
JmJKq8xsMFjjwVdfzOK4crZ8W1wPgqJJmygnpUFNPC6N8GkT/S/tsTNV4HZmM5fK
HrnZ29U0efbjCSc3cqXcbBE3RijgA9GnZwVSwhyfq19eU9j8pDKRJB4MCy1UudDX
v5NXArI8NZmoEcWUyzIszFK4Hhj+sPF6rSymOzFrn39anVcFTTc06zUkvHDvekYT
gce2zNEOH9MvlUV80jGzOU2A9xcoEMAP3US7+lVbvmehtk6faGw4dWDHyfTuCKWo
rkxou7Lm6Sqy4MgCrEsR6fMM/FUZByKVSehAL6aqsM4es4BMX2c06a9gEuD51F9X
k80/uSmkdM0qmTO9YsqTDzbkqLo/IhBSkVoimDrfryjb4PpmkPubSo81rqaDiCl3
uYruPWvD5HRy1K8feUat3OShmbsxj6CgB1sD7o2kgA4PrVsln5CJTO6LtUvXoPsJ
5+MYWdsnKC9ztiI8eu7Bu3oYbGDAXzKExiIPuKQbZZe0QvgM59/4pSfFZqFrQCOc
QXL+QOepI50cxwKBqdQpuQ+2c9fxWsym8C1NkOjAUAqduQsZ1LPLHTU3TkeNvgHH
a1WjHzxucgyvxGaPvvS/9qulbyfeL4ehgF9XmElBy5Pr4WFkmTkjaRk519gtYklP
SW77fYflB1pAXFFg6NFMyvhpPBKvwNb+vVa4YZeGQSW8zHhZ+HLhTGkMV7Ua3Fp/
e1NZH7gSE+8udWRvGhKV473ek+sbxSoKSSrIA/QT69wB2Kt94sylCIGEKw6szHFO
yYLdbpHp60zup/evOna2ENkatxvHiG24eggqImX18Nh4ZDu7F937ffBwbOucNbsH
04sNDPKcxd/fxfxYNNmTLtpW61WIkyeJuMB0G+OzaZPifyHUSHYmgS5YFf+IxtF5
R4/wDhgd3fCa5O9ZzKk0K0DsjMgvEXuESErwZT6yGWTozQleDGclUyfssVqpi6M5
XR4WjU/t5a4jBWZUt9foE/4bRiwsxFo2jQeNXAn+dn4CVOVYBv3wxkO9erktdfLJ
lIib1o5/NY9g5hJkmS40nd0dC5s9EnL4QMwrxijErJkmCI6+to/FYbSbnqHLXi0v
Ln3ek+M7EqONZJTbhY8T3PmgwYbfs7oBUrSv28mWSzJkZp7vVLn7cZ+2VWcKqXsi
NOe4Nxe9J09RKEln1O5HXHJOP92ty/xud96ViqDSSOxWhj4ROEHmumrFkaozsm7F
TSw8H/+0tZM1oC/HCTj6p0QzIVT4hVONtUS+CQFhmuwmBg0x1wu+DCJVY76+/bz3
zvrn/ScLgn2QAE7Wq2PUaZ6Y0PJX9YJVfv6VW3LAD8zHsRRcFET1wt+JxMM3MTUl
JoOG885eSnOHQmogu6sLf1aKQDjgvggBV1t0XFtWIMbCzIG0X18Xg7OyFBz3THRg
x5JPC2FCwL2IYRtKd/y2RACkP8PrqJqyKSmR9t43tsp/LVsz+aM6bNKNnRUoYGNL
UmYFNKREjKtqjrFbhnp6MuegvlK6duaM5hT5txqWqsGRrx03RU+VsfRDcyDxouFU
qCWzdwsRYZ/n7CD2pc69odPcBdmBpnorTkW00fHwsuV7Gn2RbMca1m7hCqs/XOKE
UjDt2R4RJ4uITupMJ2u3Bon/qdtsW2O3KptLO5YKe8D87L2+Oegy28oCsgWNuTP/
kQ+jFBLeVbqzHRXDZ0w7LCBFq4PLfBGjtjx1MQhvaw3hjvysl+ytLTz5BraHfgJX
Jx5Qjas1ssmeHSspEOtuwfz6VsRiaH0C9GPmJEssXk2Mu3LxWNu+N9+EJCa4Jbii
OJfORm6AEVL/tc7zBGqXiY+vK5U6HEjwQ+UZOduanABa/DjIZU8F0mZeCGBMXnzT
E7NRTlk37+hsFb491oNjIeMJvwmpzQKghz3EYJlRZIvyXlgX+gLBj0pHqM+hrjBS
d72nSWYjNLcaoq/+9e9f0zZfpHSsuDC+cRqAe/sVF37hUKe5IdxM3iu/mXMJvYnD
Rc4IjbdI0TJza99ovRn1g45SpGv5zHdNbRPo/GpZjrfDyptZOpucLIvFNMGH8iiL
Niys5/eU4ilyqIx2rgrSQWweDEV7Hb+1JL6Efr+L90gKbVqJ6Hfedj30j6qUYnqb
Xs8osXGVy9Jw1OoX/AhnQoUUXCXcxX4i5Zkg4TJyqwEZhaXjmY4Yl2WTveCh6B/Y
n/od4DeOUvRkH6o7U0oKVPQERwkIn6Zfme/US7IeYyiyfbuSJQa+8d83TBDejnK/
djYNvgYf5jgvIdAcufKM6n7wJWe+EL3d7G3034tSCPsNN8PBS0qWl1e87iHjlQeM
ouQ+JCYb1D773owZG9cPkxSVoCrpt3MHFx0LVf2j8S87uubwYk/I0QcuFL7G2D9Z
8cqfwIN7avUlPeXwLGcVAi3W+CW+iJC/FZ9cr4e8IabgnBSYGgWYnIk+6IAv3aSd
6xkohbReuTNEtwS2Dp+/OxEtx2FUO0gypUBiwcpQraQUj/aHpOjMngG8X38y0Iyb
CloZbN6Ihzw5SzXYHd6ft6KOzPzmVtweXKAyIRmXfStE4oTAEGY3VB545U0GXeIz
DcEnBnUIHBm2ipaIowk2qA9DHdZklRyw8LCLE8UbHLDWmlJ1Ftk2jXHHj3nY8itn
zp0F879RNvxwl7bS4lohUyTWdRBQaoAbKSDLLbyWVkioX3wK9eGVp3cGV/OUibck
SGcbbwkbMp9vtslEnzLV9MgMf6A6ZnucE1djg9yWorUlM+Cxe8EXOv0CaQoIptrS
Bv6KBJRpT7oQUGPhUPVNcJEXnWWGjyOtk+ia7BAQ6jLIKKLU5lKHAGaGMJOrg2zF
KKnthQGgNCT/NswbjSZmOtZpdCE19cpyuPLiDOX4ZWUFhcjFI+9IDbjaMuYEkurA
1eUgdUXarqkmPI+n7qjpfS9nP/eiXtLhuyvFeOlI/MxTSabQ+w6OmYjQD9S6Ym5m
K+5yjJ9uDFY9HvkzEGq2VdIggq4XptnCjh0UZwARKpXZoov8WDbjxb5baVJN2hzz
ORnpvVCXj67wrOx8RzU04L6OqCf1GWdbJVVKPaO6zOMhhcvbQ5LkUi3Jh/Wu2z1S
WTBpp8rmVmQSviAAZigQ/S+76dDTLluoDWPFb/8m8wG6+Gf63SnkNQSrODEhsOs6
fE/OO/AzHqXkiyHX0fA6lKkF6Js1WLcOBf9cUrA30XQSLmpwZDB6Cp2Q/Iv6fiS2
cZs/NhvkxxvbrYtr3Nx94z4FSNPFQ24sWrKgbvxABHpEZ1/MFAbCv47im0zDnZdG
4O/LzrD/2PWtdafbsNWfEPAm1krYtB6glrE2PpjfU1juQUYjrZacL9vJ1SSyJxXA
1TIaqkr86ciqQzLGVF2i/wmDZHeArIrILseSGpJUQ0/D2LuOq/x5YtCvKF5/ZkkO
8MZEwsj0aqbdj3vuLZhwQh649jYafz5XAo6HgVcWAT8/YY5ef9a+QftPq2OkcMOy
oi8/s6FmU0pnGJexyixb6KL2ow6e4Vn3+7kewm+Hb5HIJJ8rbRhyEaLJFTtl2xP4
s4GjRwu4R17+QfUhdtzQNvX0/tJ86CXen6smXl55D/GERCnlWSgOSHdHQvKNOyjY
MKtU6dg1G0IA2lOMyv5Xe0AS7DcaEZ5zJwV3mViPrCFIpJ8KLmpqOVb0sU6+7MxW
dFG6EUBlb0nLd5ARsbxL5SfnSjxCjcS4i0YqM3Tn7mPqAK/hJFkPf28jS3ypJa+A
SM4McT+LsDvAt3nM0bTdTHiDnhqQI11hztGZXZTT4RvK+j6twrBCDt0rmeBxmeV2
v0pbEMcHHAs+gM33zXCVp0Y8IB9nWAzat/9YHHjMkckAhkoTX+jgWhEHda2BsO8e
VJ42Cm2guDbZjhyqKM7rJBc9trb47ah8/95pIx/A3afvURCLQPhMV8CJTFXopLFH
dELx6FZIEe8jfxlNvPC9N2FcK5nXfltsaGMq6GKl1j8Q+JgUIqVLEo2AbXU5BPmA
Zt/UbAhlPjXoJg1TvqULtb06KQC1cRnBHeRlmFJKvldPJLBCdWhZwgNIryQkcNwJ
t12SygjztQyHWOuwhY8oWcRzLpPYlaSqndi3FlI9YqpWTzQMYzybb52YQsbyA1p6
aVAkOJSzsw1VZPn2A7ZC8hUQn+ol1Eki2eW2XVk9WHdMLFWPPwYsxzJEjgHQnFmQ
xRofReca0GAwm5AN4p72kETSCdo71RrGTbsjOwQ1lxdBcJ/v9Sbb8pQiDA6roCCf
h1WxUADARGqCM64bHlB8c4YCg1AzbCHX2W5CoDy5LoNviI/RHr4e0ONeMb9XnXhP
aO/jw5ZcstQ3q4weRHVz5DuBW813kOiQ1fAKbdNUFESj5Chz7XGAMQtYBkAibahK
UifKRYutu63nhv3DbRqitzPu9houEWQU13FJk0EDZiPkweVRBqleCtwORQRexY5H
T3mKJ++J5uIRgxSuz9RTqeHbHiSprcrR/C1AO7eKO0Ox/KHk77kVk4eGN2/g+frd
PqUHEI7Vxw41zWJuyxd02Qmvc0cbUXWsch31bboSGbuoWjYj386Fm2opqfx/PAK6
4Xjv5mg3NRCyNh2tda+QRGmRh8SU983hVS2BUpWfnwqp9afIlad/vmmrK7BAhxIz
XqVH3yUqt1O4+A5qeiJtyGGRvuolNQXXRvu4pubKATXVMiS3m1qjtAPIeXfrsHI5
QrNA44Bs7V2t9Co8Qqz86HmnUA6E7EvI3SOoNozASvocEKBhgZGgDHKE/KoJjnNL
46YfuqRkXyTUxspRNs4IsAwFo+MkBfzXyUrjUsaWWxI6drdR7eQI95NkhYC6oa3e
s8jdci+hjcd+uyU1xqN2bI325Rl07LLKinAX53S5R8K/NfybOomZz/nbo7jQPYcm
8tIdyIJ+hwgrexa5CJyXMCn/YSPNfL9IrpfMffNwzVXEFyBgFAD8JrzxjrzL3W8b
xOGJftq6n0uAl/Z4ouO6p93qQE5AKGt6VJd2qzOehtJ9/8iEU46NxZZZ+m8ZFE3T
Q1oS/8PWZl5Q8XdEWcNqq1Mce0NsdouCqT35onVwMdZNtoNkeBITtbLRw3un/wnl
trdyuUhjM9LAQSUd6JhmwPkM2j9GkOQFrhN+dr0AIuPjq74RC+B4wff/5XdS8Iu7
M2bESuz2m4xvI+58XmO7HEeIckkcWOuyCMBi3iuAD+V/x3m3pbeYSFAUBBr7sYfS
5sW9YSzMHIjoZVkjOBbXz786xYaJj3fT7KtR4fW6ns+vYkPIq3S7EE3Tdk1EkhhF
AMQbOIjH6nEeqa6gsTBqlfmqJeb2SWKl43Y1RYB95rtIyczpt2kpMH9GwpbTjbIj
2ohrgW0iwZ9/24XrUp8tzUokDrSIjOSK0RJSs5ix1ywMpJ8pBtS68pXiK7mXCW41
G8ahvhpXro3eIUb5jUlP6RnR16wIDg2a7RpD3Md4FeWDQkvAn35Q2MQ70rY/8FKm
pJkHqtn/LiTcuUboaJuZX5St3Qr7YkuATc3y05F0Ig7fJgDoEAcrHJXqyoPNK95l
CjSbcapb57gjOujCL/PEjSy5QE8S48tc2mRjGCIGv8/FHurbK6e+zpRYxnXzMyuV
SyPU1NqAxZQjJ6e7fkyimDaHfBXNqVjM5SaiVV9jp7Kgb58yNf009KTkCE8A5+mK
qD6g/ZDV20JVHzbPKRSMsO0rBLI0xZORfNyZosTOv9BJoEUpmqH9kGvLxoLM02/w
kVWAKhY7dADp2mNdG8WmQUX4jGYt3F0sc0+xHDZp17NvL1K3vCtFV61bWARbFIt9
QTh1buI4BOHn6cCVzLXrAvgJ4ROGvzlAiDgp3hAnpauGIuKpwx4wHoTxVOfnO9XV
//JerHGHswjgzK69Tq+suRzYOWcDujaQr17laVjnjOmzDR9k6nv7QpXPhehlr3FJ
HzzR9XxOR81VAM18HhHr18F0TKAokaHWXlxXeiCYPMNBGmEhbqFF5WIAYBoZCDY8
jP9RhaedlQqMWE/TClQXU7vV9qE0VEQu/ZBEN3YP6RuB4xdOr0kkrnKHdBr3l009
AY77GbmTEbdaGbdwP7fLHw57cWhhkPT/jqN9SQ428dft1QSlICo5pGUWeVpasZ6R
rW508SxPMbnaS7IbvwpRlTwJZPjhYqW6dOe8HIEoNmZOakqvuOXTJLT3D5Dr2CaN
DUoVISaVtvNdgaiYngJuxqN0JQEjYM5RVHdIVAqV/LXqIqtnvuCLphDiEHsEgt8x
EvBcktPP2Js3+5cbpPn0yEg4lVvB5bylDwi2r9bk1azymu61USV7o5ECyBxCcKsG
VvbWJHnNPv5zT29EdRwM2U3WfAHqeR+YEXxkKCsvMniWa+6PUrOnlqovJOrFCR5H
LipBE1gKKojNPAd4Zxfd4KmByVHYF+a4ZNuB+yCuxnf89lx4fsEPBinYS8bMT5xa
7E+U6hCNk9FYx1/Vsc2nAcFCt2918MUeP2mAfj03tQwC56j2e+z9cA3xanF5E8eG
WP5OCKrKtZ2SDQrwQIi966lI+z/g5ZBmBAzNF1qmXneKMuY+ur3YXyxaicen5gvG
mGhVY2vuSUy+XYA0x51jpsq7QUxuVB5qvqvoIBWWoV5saOZOmZN1oZAwqa/x68H8
nnYvk8g/y/1y2jUIUejYU+i6RANgnNzL+/O1aP3/mOptem4i37iK3G3Y6LrAV2XY
BufQ6AW0/kYwkuCuuNkNwGgD3HglMMjRGprpwFB0+jRESEpBHhMQnXoK3uAR09iw
ZfICwbVTgKdme1KOMKlNM6wFWtp0DuoL4dGIA4ZwqyUcTLrEn10H4yp2yp+z67Sg
xAfe7gjX812t3EHHWKpVSEP05YbHRKVtIfJUwIaqWiFjp6g1GMRzBryhoO6xsQD7
m/LbRfHIokZYRvzR5rGPEIS9CfNeuZgllO0IlGmPON6JwNyFLKlqtB2Kqs0pj2tV
aoTLu6m8aqPpMxXSZxb8Sw9CwWmI8bouVhYGnSDypVgMyMAOPm64hEkz5IN31+fF
O9RUg9qViNPexIqLvD/d33lvE+1GskanCP9MxRClULcRIENMiybF8C10RPY37miv
6FEq5MIBMvig5wxsXLTdJ7Xzx1SHMHlWIh7Aw0tMNik9zPLAr1uPA5oxqUL5y+1Y
dbc1ThuGTgB590uZpen84q6fiZuiigbYEQJa/WH3S4Xnqwv/JYbzJ0C8prLfPlpI
DgEdUm07jUXsVAZvS494xV5kvN0/sQcu9FQSsMBhsEV3uxaghcfjUwJyppU9jD+T
TWPH77OBxVf0ZAOp8An++SAD2N+2LX05hoj5skSNuYyknoWczmHgrZ2IQAo8mbex
OckLve2na5JoKmThX+buQi8jF2wQQ83FaL+SsmI6vAprAKPo1K+9BvvyO6S8+FI2
/gnE0Vlp2XE0/Mey+xKG57j6NQ3fgL1MDwT9OP6uREkoMiLdTlFTnqdeKGXCa+vT
o/Ut4CaW2lYeMnEmCKlkKNi8HBWBT1doOSG6j4By0Fa/ohRX1saUOWw61EbyKpn0
ZN88W/6iPcaGVlAooBLtzhMktTnjzFP9mE3vk6pokOQAXiKQg0kVSEwPnx2Avz/X
vCf6ejymjsTjdr1xUJn5RXbLTJxPI4Jg7GYRoyNt86UZzSpBmIZcepUxzd8aHPul
zhT3c3j4xWQvMpPHLo4yLwqh85vKq7UX6ux/Wjl7pHxcH+h5oHfIE7JdPrNllyvy
b2ViDBtdcgug7scFt6ZLJET6RVFb7FJyaBy7yBIH2hrA0fPaRj+3SvzC3NSe67+i
WWW3qRJc5orENyCAEhMBsOV05l3D3Y1IM2ZvaLX+gz7LO/3Ne7yHGKChWQs0xYvA
dRXVWkmcwMdOvhGgao6dir2Qq4O5Xionz+VOgCK3iquqsBveX6557OEYv3Fe4xQ4
f47RTQALmr58dvAV5907G5eH5NJY5/KwMj1+nRgvizVUeDcXbeOawgW46Po2Uo0Q
rxvBkeyie1WsV7k2VKEev1Mgtl5jiN+ZeXO9+bBoimWduDCbhr+L1CWe8MR7XmvV
pCxxbEFwJ/j6HK2uNLhO3XacJ+lCRk5ZmtlECpphzHKFckvewzdSIgkGR4rUiRV7
XjURScZZ0AwrvZJN8k8sXfNmnIcnHPIiuwIcfqWmvnnlTNWpDFHmjVeypvjB00kn
w0SW5TEM+Oe41ViDXYAKp7RT50pJsd0bOrbwoAXvukbffQxWzbj/xE97/IBKa7Vf
tNH8D/r5uGYUEQ0YLlhQOexkj0DpDbATpXZLXhyXvOfUwMsR2NwEJ+O+hpRnlvDM
VcSjzPe78j98AMdaEkDij87H9h3JPi1q0/Nec6Db6oRUotgk/HAU5Kz4qTEzRV/q
HyOJrzb9Ty4chIo9OBwwvVnfF+H6w4x0oVr8eDsIXsBoNJ8S9Z6DZJeQ10zlKvlH
hYA5CLqOwRKnkRtQbVrKObFtygkieOINrMBxPxbiyvImXzW320wXUbTuhqzEUw9p
NC4nnj33GjlFX1HlaVFS1N3/CurnrpvHNd5rJSTuxWq4lw+U5QElM6cuIrlfnoSV
5orbUb6BPbSrC/XFsPNQeEf7njLnRpRO6sjGSc17RUKhixAbRhhQ+kqwbRRrjUP9
TiL/Iaxs4PSYpc8k2szAbe9AzTrua0g21Owoww8UvEwVIa4PoBNbIesI815rU5kA
aLPd3bjU3M7bHuULQu9IupSWo8myZtlkALga3FTSq9YhROxQ9x6imyackdLawlCp
nhOiEohk+B6gp9zbsNamz6F33WmUWBO2vpMRm/8ay7e5whVVy7I2xtch+SdJReLJ
fH7o8yOdA0Z8cNkCuSY2RGbShFKl2b1D5OVwYKrw/Ibyu3wKcarBzx4cTAUjB74b
n5P7hof6Lf9gwf0ZdmjSmLTuerhH3fHLS1pIsR8u8wmYuuOO1weItvgoeRd8W9Kl
dAuxqHGv+4UjkSxKOEW8n7hzXDheg7kH5aEWsUzcdykS2CkejL8DKv4yv1ab26aE
Ld5nEK+xRy9q7wbRXQvfpwPaCPy5VTZC3kPJKAJ5xI/Lydhoikyf7HRypcSXKJeH
9ZWbjRgpfW2whnK6laDfmmVzO6y/lfu0UwOIQ77PbUeKY1Y+Ax0MnDsW9u24WWRC
bXrMrU9CpdOXKoFkSd7Ig82FwBsHbWZO5tWkODSruI/mqkyk2or1KA0PFML1SaOl
Ru2vTd32gQTcdPGcHOpERQ+5RFKEsNfXkbwtTV+aEgLZkdOG+1pTCVfgz1P/9oZx
tQ366dUeyicK/10eeilAV6txfANpdtXeKODOZRtoIjLXknt93pMbVefOE0jGXT0Z
g/WQCG+OKmO/STYRK3YzcWUs5Th8UPhXDD0aBK99QNoeajxzkB3l46qHkqNC84Cm
qGibsGkVuqdawNNq9dhKPbmAgNo3VjNWrRXNDFT0KG/yI7z7AEGSGjsxu0EAb/lp
rwavfYwnVSMnt5925psv6Jx0I3O9TsKB17xEzn3kOkCdiAQWz/beqqMILNujIpaG
h6YxzeYohCsGzFJMxQFzB3Er4yxqRfkA5iRMiuCk7Jr68tjcHzjRtLh8qaFoh3ns
hqoTDiJpAJuZWUhn+7bwPd0yETxzH4Gzr584icOVtpoROLyLxpZvfPFA6S7yejN5
sGmd++0ej2lnwUkAfFY06JiN8Ec5R3ZW3IWrXeDg0aLqQRd2iOwYqfJ5SCgvH+fa
rAyi3Yo6BjZDVf1Xx32uLVwxNWdLxUp6bS9keGi3IAl1Loyx00IQd8dB9j+cpYZ1
5tk+Q6LMxZZHN009dsWp39s2pjcpfAOIVs05XiKNi96HiryHujzy7/NL64D7r6rp
8uK+68oytTcvwQ6tluKa1o7jcxJuyWtIbOn4QiFBkxGJdXVAfVZpitl5Jaxo3Z3M
kQK03gwhkZ9bcH7dHFEeHbpPXQJcAkqtTAc+7AHS05HttVOcaYhttFZGGLxv3Os6
Bk97UrWOZZ9bs/HUQrpU+x8qOAUK/pgQnN9HDd+Dqbve7CL5OS+gTXRGRT6FDbhK
z5EenQylemLixTSrSPNWqqsb1IkMsqf/gaz+LzHwjX5CigjrsTcXh8dQJ9isgbx2
1AOsqvJka9bvaE98cOn06UipEbLEz+Ylj/ypcQllIarytgB81Pf1dkV07z9rsqL5
8oOoPXoZXje9aRJ8x66OB9k/S1Bu+dkQYRn2ZesOe0WQ0CU9GAu14ABRq+1iXEbd
NkcnW9XXoazaK9JL8KGjD8epQVFrEAZ5AVxWZVTFD4pANhUDR6RsIT/f7A/v1cMJ
hgPPw/mDGsoD2icGA+Osiat9GXcySOSqI3+m3PX8lrLwVPzK+R5qbbuMel2sMye+
Iy3dV5qPXft4jJ4uIGlXUf6TSUcCdDyKWLxx3EN5FWPvoqjBcjAmM+iTYaEiDBUn
NydM6E95k1j4aK/X/Ex+ZFa2wSsDYYReTgVcbSVoCQAfAZR7A4EDzKVZ8L18ZI2U
Z77By9uAFlKx8n7rRsGGx82ORc6LqIB8CCaYpmS1SNqb72vVXZEZwMYlTvyEUMyF
2FBrf7XQr+S61y++5BPnmCN/CVJxobuyledrnV6TAa3FSS812AoXXnrlwbJQnloF
I7Fuk2VCeKiTD6EDrAODFik65dz6guLy2lDc6C+t8mfsypNNJ6w8pvrNw9YGcvqz
ogZ+UwWqCccuMpVN2A7J0eEOZjuuwP1bwfwNOommBiuNxGvbm76uZr3xhWCHkLIH
oj/P//Uhnmx3Py5eFkfDo+th86aIAwKlpi4TbWPyLmRU/TSm7wU5prFWscY/Zn2m
r3JwrdqwGUv2R/F3ZNDEvC4oFZTGsQ6Z2eFAtDGMWHxgw9OYY4EgKkQGxZpoPloY
jykiZOOl1RIkNY1cKr1kiWsq1jqaNj2M0ETFaOg0buoyrFy8O6wFOB/IZFfeml9L
EOWnnc+caXb3/4Skb7hA41ubtedsbLkv9ES4cimZO2e4ySV9NGXK8TM2IWbwDF0T
iJ/JRZLr184hB4bLECyrVshwu4pzjOMUTVYDBMBuZi2KFGfGXiHz8k8Vl6N/yLCv
Nxb02K62FGwwox6MDWDMr3bLl3iaHbgmf4+bCfM+KQd1Emz2ZeEVq6Os14g8UWOQ
IDaVy0L8cS9+pXwlVeQnicM6AwKfu8woNr/wcFhsK2Kpn0XhijhpXC/RvdjqGWNO
pMeTQHaAmOjLkEjNwOB+ejGxSBdyiu5YuVAGVw7kl+nE6GlWLt/JKmnS6TjRRMZ0
wQrQjvf0dwXtgnbOD3PKtAxDxNGJ3CJx02XO7NrVHh37WjNHvxpRK+KJi7UAbSfZ
7Ynx7445LM2JDGDYgBLRhKgOsEdvH2NhOmlNJXDm8c42IrWGRTbZr0m8yMUXoOmY
KYN9unbbNdlXmDzaxrqvKtewcpbusJYiLVxcexRQKKJKHCR9q2XpoJ77jW++33hv
R3W/o7IO4R9ZHIoAJGkT6DlCKorJZ2wjAwqyLJ7npcpp6d8x+6U/RPqpYjvkN/w7
EXRx92Zu9Kdk+euLMiz44qnwOY2O9b62GlfrLIxL3EMhzzLJT7eM8HYm3apitz4N
Y5lxiXxEi5ZmWwr+4a+j/g8VsMR3V60Np/arjkJqEW7uNNQc4BpZo62Kq+6l8Soq
uCWrRUiOIX9Yjvpx2EzcRLUkWeDJhR9qx20PNxOOw3IEm/2zBo1cYhIrZX0wgoA3
gMX5yRTpq87rlXpUtljRCnb/Qg2OQrI+DnVSdCbyA9uFchp0d7mUp2BLIKiwOlZ0
AAo3f5ogq1496kKb6W3yW0uP9WD2t3giiTcg3S78eBACrgKx6wumcdqvEji2hdgU
E7rmun5D2rBfbZewFEqKTh1Zab/FYSy5iVLYYDb3aQ8wd2ZDXkVuJOkw6VFUq5xx
Woxe/YVj1Zp6tlr0A8rB7WMTWYtk6WzrePA1rhOt+9/MqtQNQOhooxF/CduV7y4M
qLjoCPJ6fMoaH7MiB3zvq8vgbxrfnJFq2pigA/KzOrIDWZaL8Swtcz4uOQYLd44+
7IHYkYTPgibje0jqNQRdGy6hoPymX7tyAXRARD58iv57jkz1zEx+tAgniEJnpOnJ
2BPOJJBnKct0jYcnmMxiII6kxfukBL66OvycwJIOCiOyNUNNGWZOemhm6nEKyopn
Ic+UGtwxgAt6OMu61tHD3cBSt9T072Ol+lct21WddMHlCTY1viLfA0IxDRVcCsMl
TRaaZkLex74UaaS81aNV4Urgx/LRdnzBoek1IvP8RSN7S/DsSDzEQBTmlaTlMJ9d
LxYb5JAMc6Xsslh7SkwX0kk2Ltgq2ENvE8Yl6+QWuLd0Bkl/A+ovFyfEOWILh8vV
BG97mbZ5B3ZzkZhPkYSGv7WAVDVLIgJqWXhMz+MnA9W23YFXMcjv4sNv0Slj48UD
kWZAyUm2S17ABcdWrPwkcqARrMdwzUVJyaMGV4HzSpHXf0SBySO9TpYuKnjKGEqA
nCkkjALhy7TYmaPpdSURpEMrOSucii6qDZ6I95juh7lU3rRrD5sBOJLu3wnIIJI0
09JACJstBOMuLtLptgUtKfwcPbOf98ZSm7lhGB2h0M51cpmle9TePigBYzfbMJD5
E4dBG/yHBUhbkI+SjxIyxkBQ5aApCuJyBZpNQ5K1rnj20bLqvgkeBdYGkS7Wd42G
7tTR81yLGDPxlonb0Rd4ItA3DiCcjE1aqzBJkE2ujym1sl6qz8ZF7LDrRKz5Om3J
Fxfs1xsXSEZ71eYEU+mTAp6ouiDA1Il/SHaxKrcFKsRYmltRlC2Z6/AOfsLXbinZ
aEVdEbBSAAMmC+YWDNeOR8C0CzAMRTWKXorziAbEjI0R2IpY3aPERrIqcSBuOg02
Ge2CBlhmJxEt589QYYzBX7kY86HNLTbfSMbJ4Z/UfSKbCzVhySdUoaY5lkohavFV
5Bra6XbzkKn/R14+Q7rAItsvrOkKx9INE+cQ6SAedzcP1a4/xSOe9XGhmFsaZYAg
fT1yZMXLcABKxidGZPlhMhklB47fcyIvQ/isMJaKsfZcaV3IwiE9HLZrk7vyxNEY
cyko0uVL74Nr13XbxhxJtGovhcY/RrwXWuvMV0xd+oSMnr5HGhEuGFmw/HZzDpPT
9R6QfuFYPkdfNZ4KatqYQHhj6pZf0bcPmR72gG4zBrnWptY3sgi2+P4e04ewz/mo
SAuZfAT+l97CkHQS+GpSt2MXNst96FA2YGq8f316AC+50fJ+Yw388f4mVtPaZ0HL
G0U1kVDw10t+t0CFbXZzCMH8HZCWbsVtpIRZcvizT2epqsdfgyl/bcKykDXseaBv
yG835ipGsyZsDlmJRMYilWmShlSBmRLwet7yiZNreOtObpq5aFZhlfFbZu5Q/8ex
nbxHdm7SdUqwdrizDYJSzq51CVph8PbLHwgkCJfkbUWn7y86Mj6YHaZ4fcO9KlNI
Hsrmub1qoflpOa4ZsgQnuctxkJ7rVVmAbJaVaC0PLZiTZ1/SFlsZEqfhT2AUVhjT
rmRqKEug2IqRif7XYWlI3sRSCmM+vQNFiNXbOatGbK84LYJSfoQIxtYxMsGhR3nY
Jb8GPt8Q52iv9qCswfQG6MV0XFmvIyZKkonvLY6BuP9gqEQJzAXXSC99f2DlVAjm
IXO2PcFNkd8OprzZq1b0VU31r2wmVZ9NdxoAj60BE8lAdvdzRZ3Xuvxs3E53XVKH
Rcg2xp+gTGqFKTN/EcuzNsjq7fVR/CoWRnZXxnjxKVxuflO2RbVXzRke7iaKBOJX
SUJB4Mt++Rm2qhuuZC0cqSewKzO2yDIRNGoOLKYvQEa46HP1wIn7IvYcTH4WbqGC
f01JgWLQLPynboNxMvYx0KNR9BGHKKlv30734VnqTkGpU0N7gfuGhED7CiIcA+27
+/+B8L0Mr7Cl9geFDYcFmuYY8XHXAVPEPalWJD/Ldo8Zc/McXPI2jfgObichbEQN
XwGJXCkW8BM5MZKhuBNTEOdKhZ5fnr4KLK7JU88JAnLpOJ6cJD28uJsIuMkYJXSD
zzutwJ2DpRFcMv7SLCfFLlXbpj8qkrld6qiViwWUOdSVLZSjX0097cjJsx4SBPqv
2q463cb9eci7M87ysLlYfUPn7Q7VpAddl96uwo/htZlbtVwSQjU3Il7ejSaZCTcQ
A9QGJpf54SmsHvxp65OISiIL1bLGoO53t9ITCA8+msiqPjAN59S2NHx0mcU/G3M+
Qyx6F30ea9r9Vcj+ZsCq3q+atpopiK7YJ5CV5CPPhGWjmxxxiWJUSGFugy/ic6T0
+C9W5aPb+6VrPVjO/eh7aHkd6kajhCqsnh6sCcSN/cNqG7GAmJw5wGFKg4vAIFyB
Bsc8Uk6RHwWL2AXQ4KcozHs90ahfjlf8uRHkTIfHxbKHkoUqJmLKYYzEUcaGRYyr
tLkd+f7k13mvdIwzhxrJneccebNukNQz0Fs1esb80zysLDOc3SLPUA+7gwGntORP
CTBz/4vFVfVuW3f/7Ca/UAM9uuK/k/r3eUuZ7aBrTyE/cNo2gUrv6f+nJA5vlt9M
vzCZYRRFG5Hz9YTlRRVZ7HbH0vysHmw/jAdlzBF2y9OZeI4xouE1QgQRqwa08Hyj
E59YBZyTpcvHMa7zpG+9WSDvb8p/U2ORDHWOsDP9DCCzaT8iFjjD5OKmxWkqcd58
rQMBKMWvyeu/U5rlmFTceOOjCcR68C/1VBavH8CQjvTRwBRlp1C28Curb6FkkJDI
wo3rkkaaq5IPLdLf4d9+NqDKPn1XGfL+0/dF/aAGS00henDlpUQIo6gLwxcKykPR
m2UtIY6cBHCsYt/mI7UIgR+x+nNBBcqjllx44112dJEnuBEmJ4N6XCVIh7GM7b4h
DFAW0J53YMZSYmbYZLAz5SWc9rBtFV2GCRZSHhK6FuGzfK5U6Dcaq6GpfNoygPgQ
DQ5YY085sn4D5CvZ9gFvJdih0+guPBUO68GJ71zfdHBGp7iS9TNL6vEQB3o1zNWr
kVSdJ9yE7TGXNmXeYbzKify1KQFkUO6c20CbxswD7RjjsmLL3nNHTpJMjsKthrOM
ae+E9gdqBKhCSovxXYb5v2I5IZj5hmq8wOxzR6bH1kssL6VbMImXAMnFltBg1qAn
XKx8CPZSCluPGU3uxcVkmoSKqswzTXRwgJPpqp+pq0gW3OE3rk2QfLAlhRwe8s7L
Tq54sx/F+xJM9OEl3Zxs6rvHIsDFUKz+OmsweFhB5S20ZT9KRKHBmaNB1gkLbP9F
Mm6Rcu1ftmBOkbgUkhoS56JCEfdGRDwJOmND4wJJRXl9Ahry7Yg/lYbETlONEXLc
uDuHGkgzKpYT28UENlI7hYr9a2bwvHqzwCXjO0e4RZ8nKOAVoNBeXEuiSwXfrnvW
IicdRuiEMdBlxhI5BD+MLy9SHqN8IleLZ4KfoUUduks86jgFr1kZn+kCqVghmxd1
ZiEen1tTpZX4W9mxZgAjBCFPu55B1LcJ/cNEj9D3NAEGjZ8zDK2SaLEyMimCkaIU
JczQ7WWsUT2v+LxZXo7iEauBrQ52v/4ajszEe8x/JRk6dUWo/Lv9tf9gpmNZLl+y
MuBMssbbPRLC6UdpLikOfN6bMYmWj1oQzA7oHvENePe+IR+LF27Vb7xc/i5lTDiI
vkkqsYao3cr1FgPR9YI3nvbBdHjWlW/fkAI2Z4Pg1h/0vcSzpKCTYlx7q+dtc3By
pteAixP6CLqsIwOGKRADklRyuclpUwzEOzElw1uGjg8u0XlJH4iSepPK8BEy21/Y
mHDbpLo+W/ohV6/LWnG0KCaCPeTla0luboa6yiYuKLvTwsLjonekuYyaEgJ/zvDL
qLK/pUuwmpev6pqi+0jL6zIGMSeQR4lS72eUrzx85mQ3UKJIyy8Q0aYmXlE+ODIf
ci/tt7eStwim9cjeT9OO2U3fDNXH3GKL4rzXcUyVcVJYDOtqkzFuZqXS7B0ftmrK
AsXJbAITiYNzJmgl5ywRJeSSf3xp7LLwOFKlt85SbP3ATkWvMoytEYTIIszE1TXw
NSmtxvAYPBa/FeufieXor7n1osdDG9vbiKOJB+x0pBh5AWk6ey0Az3v/bj0xUJ/g
kRCqa1gCmBcKeH8NlFcC3JCcNTUYBiiWkaXm1JHiGlgHpFvatVgtmYmk8zeCi5tH
ycOJvp62n1ycwafNLjyzm/9sfCdQa2sIVI/v7ucqN7Yn+MNPv7rEW51tjzxrRYxj
wfvQoOuJL2HlJOgvUtwQI1rg4UxBfhoPxxSGXDBa335THV5QXx27w1+7riV0hhCB
EACxC8M5t0p9wNyJ33RpWQ9+gmU5OMTdSh4oMgOiKB8RYoR7CQvFAy3RE8zhOKzk
8KbFANX5QuwrO8IAuGz3A3eBFX6b/bPiB2liNOxF/kp8vjQQaCTUkF9VFGDPfuuL
bg/jIH1b3hzvvMAhw2PAp9Kk6SjBwSaPOQFO1x4ldVv52D4oDSsz8ZSknwHHB5Tm
+YFmKmmqF8Cf3ImTAn2YVphPR8zwpgV1TfSYHbJpi07oA074tBMcnRsk8uNiQmJ0
lmOqyHtgQd+r+8SMzmjjdBDXjnKjIoERhpLGI6sIKYXHAX4S0Zj8Plk7GdxGh5tp
JQ3A4a0VBTlglz3G2Mgw8sm2FcX/bb2MRcaz5lnHseCCSuy/ZlQ3fHRtiPeSxtQS
ro52TV32MumesY9vntzp94ziSLsXneAQOLTVK3tp3mgGz2pvYqR7QMMeBJYSxLM/
uMdlk5DzilZa1rsrKNOZLPpd7FCwuu9qjt3HDBuBOiDTfM4vlMUWpKebu19O1k3S
h8rRoeNn2N7uLiZR7VrE8eeO0Oec+4sL2KcitrMidnoAACB70ZNPTdugq/EAouTS
A46wDIRR29nl+LCvsa7BJHcOvil9I+rJOVSWm5JGDKRpB42WFsTkzJ8+RZEehZWi
2hnzEOX/kCuNHmntP+kW0MQsVAU6u7ntgPi4W+A4bYSCV/sGLDswdLsR43JLb4wE
S+oLIYBtFozGt/VBztsq7Qfspa/XPyfEW7NrtaDmwuqb9f3ii/FMGa8U4ni9Gi66
BWvc9BUm6iHubDOH/xMH/KY0IDS2t16+guq8eFxmGDloFiEX1YwUirsWfX/rFlOM
RMEDEGk0Na9/UgJTvQcWowcp5aBqg6j3TKwtCr8xA5v1aGwfsNL7lfdyDbQXXlSF
os+Ch0KO/t/lG9BZQOYhSJqlUUSMrF2ekKtv8xhRc/rQA6a/A7WfeKaaBdnbD5Ss
7klH+Pt9LrAqVrGU0+y2rK2P1h5qLZeOxUHJS0sQpkPCup2tb55VUOQbQwhTsu+W
UgGlFM9jNgNh4lY0/dy9yU21icD/DjL5ktg2Tnoye9pOLszpxiPNlueKcyq/FoXr
6yMQIEzYyyxy5wNOjvPEJLijZboKijWZ0o93ef8eAG2vi9PQ3ucdcbtFZCOwevSQ
S22+6TdaqUAruo4y03uAASMwYKX+m/9UCJBk4JCzXJuCAc1vGQCWsu5B+lD0r0mK
xaST9OqRDtHjrovWKjciHPqByOo1atCrSzQ8/2La3EkU3C++NlnAFfOPicKIPgSG
iDDVPnerqcr1tuyq8+GlYP4VI+l9vclMxgaOQSTisZUDktyk06NPzaWBsemX1wWI
nYV79PZ+aAZkIALrsuv4G4M6imiesWiSNz6R99W0jayeHLm6yhcCz36+LucFEoOX
bul2eHWzh5O57F2y4wsxZoGwXlrJgNT2FOVXrkRifLaT4q9OBRkm1wVONBiwh1fG
FiXjy+ljqgKi3OR+qfoY5rbjrqvOVva87WFYOnEM/9yJY+yWUKzioTTXLclv3l9J
DUaEZdfRZUt6ZswmuVTT5Yoo6umujjdUYEeYegX2K9enGsNYLd2LX58aN2rxgXUB
gmPUS0DkBQdpMHmpH+JD8Z8cfAYkI7Mxd+5pKwQ8aPIJMO06HlNThwVdN+sdbHE0
7d9AeDwwwvudf273nM5VTFiv6Tt4qRAQSsuSgUKj1CZxgvImHzHiU0eJWYy7daxD
U/2o0RQNWFukTDJ1ZY9aEf2EiM7qNKws0GW9WA7H/sY/qsVPkg1r0j2dCRihZlOf
qyh9OUhBJRrJAdPuxLeiKFO9+R79VS3zFY/R4aYzjCqwLscW+11gFZtzMYGKRGy6
mnzwgA1rpvty65XynUsr4UroJFDDwNuzb7HEkh6jVAciX+f8Aegh3AnowwTLHaZd
hbLJ4z4QBOfjX1TdrsrDRm7hmzDk2KczdYPprd/VCtqor5zhDH8m5ttnYQBc5Nab
Iv1rLvLjDRKu+sRsE42h8xY8HBOXAHsXoLeHH5Sdgm16ss0Xa1P87lsZxgemizCR
EB3cUasMhdfxmeKeZ753HIv0+jxLfxHp+bK9uuSapFSx6kCzp5bgKz4RwyEeOYrn
CgST+ZH0pkPDw4ta8iNKDenr2fz020Wrg4AGfznt1fEL9Y3WV+kBZ4J6CcEwQNDF
nUBKcgd5tb1BMSlYwolgMVaD2xPM4M2yo3BF4Gv+FeeRnkiH+qL3NKAT5/Raaz/+
DvXTgwKqffyYGdDPrlBN4De8B2GQVlTWdy+8Q4NgigBVE54vUyFmKxphycWSKxAh
Vlsst4helIILFTsi1G8gLaOurLUpyfY4B/F4OvEVii6En7quhAHQsmr/z3ZtenoW
08ayLpJHxv91cEr4jYhLM1D0VCpekPTcUt1k9EEoQ8DM4qV7F5tKXXZz8Ao0ktkT
KT4qsxh1+IpnK2LaMwPshM9+vi1bT1UedsBY/gTCREDzqZuUuhQTZWEha4nfGJp3
bS+mqAEKssoSlDZewEIBRcWZGxZJ7TUOa2Ys0WcCtruk//H4PFXi0LHu6IEV6H4W
EqlLLOcg6oPhyCvV2sntY5EzXEuHrA12PGkQSv6w0vjmDqVGQuF5dP+I1fGWqTSb
aslhap5ys1zwTqo29AWeB5AVteNaAJNk+xXiWKFF1yYFkLl+qbXlTZXOFMhq45UL
FhrWN/FNAE61socRDxSi7DiZmLwWWmHgwGjb5YS3YjVqBQajAIu7ejkQSF+Tv3fK
cgTZsDuG81PjkIsVum5l5Id2M/GeXtsNggC+rkWVOFQkUJHihz0wPfVyOIElquiF
W+kxA6chQe+zNzPy1KURxtDVoB2L+dSZLOiN6GxUa9m41R+jM2uexVLNDrFpw+qA
gaUgiKqQuskEFkIN0TjgbJbbFGErPFWfrznZpCmw9TiHSlAYs1FWOMon6P8Zr1EE
ZwsKZnc0Px+D29joijAyq1MZEHD88aMqe/XM+5YatRDXHRgxIdyG5eEJjU4H1kuY
L/736cvboG0JHDcLwGDWwwxFJzlj1YzvaY0LxwziP+oP1hVTvZSPx8/U6S7a4qoM
Lw2+f8TeMwdgpmSqKZMTTK6gSYwXsvTKP8frqKoOQYPvPQKffYbsesBIV266AhJY
3FrlfI+iMTZyLXzjVyMT8P0YQcbnhCJStZKdPPAVEvZhNhUivG8ivWuXFFzM4owM
+ClmmcPa5YG5gRaD4DWYFPH8UpaYvw3eUolgK8bg5l7qfi7AqKJ57rIAAQK9T53N
KeFrS4wPrX4Gr47atrDtJ5rjLsu2xQoSl7bkispii+dvgqcYUc2SHaFaU6J05oqp
OXwLfg/DYxWUTsXuqJ5qXron6/YrOi2/FOQDJhlKbyXYRyariZME/K4xbncA8Owf
jb2AfyxnTBnu8BF3KusUyLJsf2huKjTdRlHbzYGyn6apgcM0CQjB0WzYpre52/Kw
5Sivg89qL26bdxm1aOFxSTbhcjO/llH90aUlfrIIlBSzIzuF7D9FRagwLXb6k8tj
EkKsNNtrjoCMAlD5hBSNolS4b7ogwkueRUMvEfDZBG3mR0hKdU2OIOFmcJbs96+L
MCs53t3pf2cEVt0VPG3vqXsAiEPGezM+1KHB6+IJN5r2IMCGxIoynxgrI2AK2rMz
O8d8TIAvF09t6XhxLZ7EX6yes6fmo+3h2x/KUdcZn2qfX0vgT14CSQ8RI4e5uVtp
0xwksYBAczUs+eK8RS7C2too9xNFZ9HjwU2iw7zPDfP0NDI4JfU9GjGXRYDIwRMA
Yf42An3XSDGuRkoIfjJhxfUZr6ObWdVvRhCN/yqUBH26qTMXsST1ExM0iD/FLv9Y
tEUmWAT0WtJbtSjXgU7tb1AfJspMmFDv5//wyFlrcPge2O1NdOF0I1xjgszzwUDH
XFfwB3NvitDx54QJ3qLUgbMZqKRdORqsYgci3YS8Yl1Plx7ig/7p2HRZ/ALUx84U
LvW/AVCK002229DU72fzNpAZLqGqLfT5J6tRMdIKo0Abg3Cl+6uAO6zKoE03i4Yy
slxskYay7qhV1FUbN1mDmdsbREBZbiEX74rlr5qEQVQslzAmHgey4fU4nlV6ms5V
RS+t9EDCTCOyEEC+7M5DF+zbsYOk3Lv8STrHQKG0BR7GNvGW3QyPe1iXYMogK0pz
ByW0Hxc2MMcIya0eaZOJ4StZgdcgBQ3yH0zgxoAYU0aaj2OgGx1LI0D4ES0WqWsG
eKm1Em8w02NDLOnUs/e2EuZ7wjpp6lNSq+VzIk/QxqL2DYgHaoJkQnfrrmTB0qut
O/F654VabiffYD4M1Dndw7OTS1ZRdgDlLvSOKY/4EWeGWnQGHtU0Yz1aPHcElF1h
18igCuGoD11Be4s7ALdNQwRuLKXbjwiRqH7Cn1nrgrO4qgSyy4KOzR3a+avVffai
15k5DEc2LdpxjL9Z+TGPi8OMk9oASkMjyeuUW/VKpWTGu7ctInwQ52ptWdnx14R9
ciYIyiHZbkONEotV1Rp+EFlUHk1n0nTEL0Yyk79wHsSBrcTRaDBMp4RqXga5FJjM
rzLByGBsevrePeUWyOTtWnPY3jyYX4kA8aVr6sIlLMSuLSjvKfl0YBvvfiOOCUFv
mJuezZZF3iuM+1cJ6BnnQoYP3qavMH7Y77sFPUDJY5ZFsgmEICkctHyQBSm+HMcZ
KZztByyHFUmsnpL3BTrGwPvE/ng6HVnoGMwmeE898b8UoM7TN4XCvcx4UwoWlI/Y
XjpShzMd51AQuygcy0xd5R42Z7yHBtkAzTc/EqJY/LnA/L5nCK9IaHLxtNMppJ2U
2+4jZeASshB+TGYQ8PzpVGP7bXjvUaF3b07y+By21AEjSWoPGu95YdZ5bFtD8dHA
vcprGb7DVkD+ATmno+TYZ9ZylYiD/VlhJjVBIt3IFdnE2BUOPOk0rOkTRInG+Mu0
yHTCshByfcw0cg8Vxwq2x1yBt0DVJcewM/7tDeVEiTKxlgnmLWL5iagGqIObUJ/h
2bBHpVwN0Ry+/8BDZHluNfLuODR1ldAwbkJC0rsPTCc2GBngSoEClN6OdbkGoGM9
nRjpSfohqFAhH6EVek+3zXnfpSgk/ljr3TZWFejCuKdIg6OnRhCe9rhwU1B63Nyk
D4gFi+XPVBqleemWZI4hA4TwacraPVB+0/XVx5fSuStZVll9Z9FSpbgl1FIqNE3P
Bb8t2yx7FF18lOPOcYOf9Tq5Opf4JZXJzdqceRLQ7xI+K1PPYvDyQnwGYscq9QUX
uY4TKplqTo7NVC8I0Blex4CPiX1bx9dWfKV7QCT/1ukSkIMr0UvHrzqzNAGGLual
VHW/X4+H/r88Imtrrob4MwJ/kwYKAHM+NVfkN8TyJepFHMk2drz1ORJqicHVUzXW
xrcMABSfMVqLAUKI6YToWV6lnlCE5bbAHlPsnpu91mSf6y5FNwc4uOVyjZIksHdW
RZNWmxEmnEZti0S5A16umVuAzj0bZaRQtyH6pM1GE7GZ39U5j3HL2uazvTnj7ndv
B6Ij8nMMUIPisNB+KhSlu95geM4HV+SA3deuGPazBhsAQv5JFC7wSl2ivAPS0Fz5
uEtdTsuGTLN4mA+1fUQaDcLNjVqu/2WUhCnvPJJzOQCP+c2duIAxsAKSBe/iiIdC
/mIaBC51dx4jJBx9FYMAYHeaIaCJ3x8PjcERnbTi7CcyhwRMLQkahamZ3oIQ0NPu
5ngat09fZqOR28mnWlQbG2ZwxyYWmG9A3bltm95PilkmwdgRE62sJ24kuGoMYiSi
u57VqAMOJZhRxnF0jOcDqQQwaNKeTJz9Q6/VbtsWC9ZF3HCdAyznqA7BomQG7bE8
AMVQ5DctWbwPvCEDujEcrx4qngfSHTbgRPTOv2ctC8s1jQDy3R7lvE1gADsNCHSi
sXugHzd5DvEGGVTBhZEOoZsYQwQslpud4xBddt5Gwe+VRpjby2a8L4A7G8Eh2f5S
NXkvBQWQmQVW2wIPOPw9el24dsnNKD63hJqSVlsHueFqjcq4qZCPCXAnqWVVC7Rd
W+hSutnseZeAaIXiGmRL31tM4enyiT+jrnZuOXQWZFurko+YZvwtvN4CxdmucCaw
e8YQqG5qF7otiEBERpiCLGn03kV5jPUzscz9nPNk+HpEFF/Ab+CdZxTbiRr5xJWJ
kPyc0+A5yyFz5+D8aeP/nv4oBb5rvmME/0WVobIMijp/nF602/d+mbi9dK4mR801
v+DJlWlm5wKZM2rc9nD1F9X10jL01vY9nGqBxkXHLBeIX2xCpXO3f5Gamuoatqt4
vuSFMbWNqhJPBJI/jlzx1vDlgQYcsFIvpNsY1PGI9Asd3MCu4VTLbbuiJGeQeYfV
FpFFImoeEORLUlxLjqbO18EmohAqRLOKNyQ1MIhyOq5zwQxuirixdiAplRtTIYAO
OxHdh73aVIxqURbz2MppTYacfW/qALEfNZWUUEUEyRv0m/+suuJS1A0pm4gV7tUV
Z3YI6oVvIMy8PgTZ/9Sl28SAMUx9zSgigu6iw+a5ALfxFtiOpWz6HhecHDXpICrm
cdGu0WphCkfHzqRZnYxD5MRW6/O4YfT+V9o2axWrKx2HZceWib0H4/ZsIzIU+HJp
k69IGdJP05+Hd2E5lU1LPpA/6HXXOzkqtFiniXJWB0Kbso9qjw0jr4SaZpwR8l3j
yMrp7G4sbBk6bwvrZwgHvI4bV68c3RsfEQhgtKQRjbOJXr5EKpgbSFekahI3WIwh
DgfFup4yghmHXem+T2pwpiNeaH1h3eCH5bZ/EW0ahv82D+dXug97RSCbd7W2LN4D
HexYxsVjKI8tQ4txdR7voA69X/Hmvq9f+f75MDPa/xSYo5+yMej6EA5dKREiw1pg
xbLv3dS85Fn1/JbWVkOopmajT2bbYpqfvAbegq96vzvlPVoUS+2HzvMcCdGfluj5
Nc89y9uepmKvYJsSOKWQK4y7tQbhyS8MXKOlJ3F34WlH01nzoc1wmvulba5Ds0sP
RN074oWBs6WkxteSHCs/DR30nv9zBc3C0iYOoTxDwGpOLIVfk+KbABhWjzDAoNKw
upAsBUYPOkyTuxuKRXDWtmR+OnuwCUB71nVLl/JjAnZOyStmOqsSh6BjwGF05mtz
gc8XCtXcm/C/7Alx3qmxIFr8S0r+x5i/CJzOvS6O+jBnnFBQ4uIePAG7RZEBWCq9
vYP6OohE1R23ov51CTcY04EpHJ8gb5Bz1gF8T3A3fhJJBeJpnAwlfq6xOz/FzV3Z
Ka1I/1pUITHoT8YBhzCxEe0iPZXug8iNhoeQNC6NAuBpASWgD4ds8db2Q9OOPUrk
NuoIA33lvPoso7C94xz3mDspGqRBH9j4EyO0Z6JgYzn4ZI5rqyd2g6RZbjky7NQT
X1dsyFtLF9fBWu52LBIS+YehgtqEKFn+KiUQC+5U1tlYdJ9FtdgWvdHz+mojeQFb
/7EBYzFu13wkkrqXgS9/INVFXNOL6Ntjpgpm1mgdS45cJZxrb7xfm/9Lyi8N4oKr
YkCBUUAWoWBJzcndOE+LZImHVmcc+CbcgvtD9o+r6RkGVHcBl/e2HOc966BOHyD7
zhQ6028Yx6Vj/1MqJeI/Hc1mBbMaALIc/8ljCmocRIMe8e96pTIJ6KdkUaFmYQTQ
0ambM3bBuXcocRcklmrodKZStVu/OzbegKihcd+cvnLcZ45BFajOUJRNdY4kjL9V
Ac3OTa+SCeSt+UZiH68YviXPaoKoSkfX0Mym+Ze9AdX8/CLwHpEI4iQj4vPK2g1H
dYi8HqEdzOsJWa7/Nubc0vWrfYHPENxwmujC5yw+5lJIhMg9JEkz3jade1wSvwDB
wwwFoDWk02NiNa8CtKVO0J//4eXIkfPxSZIWJ8ME+IB6qA9l++QN3HAtKFjeMAk6
NVLlMsEZRsmv1RCkmV4OsXngpjFEYu757JWzvx6UuUM2PZF9jSmosI/laC8d/MzR
5RdVUD2aLectObTS0dJhD/S+uWbOpLAISRCTUKVxmZ8D0mMXRb2vYVhAe9//xbPI
x1vkJJIJhuorDqYK4GhoNo+LbxS+TGQsgqUTT3R+JxFjxCudBULGI6VxAfvBa1E+
8i2ub30TvCS0xaxyI5JQuq+LC6IW8HRMPxScBarEqMZE2VCF67tCfvLRtLpxdECC
oWhtxm2Kesx75lgq43N3zKpJE8HImK2JQ4oTif2QaaWMouiwZR7iqaShc5eGoXd0
akopp2k4dX97lrbHFs8Q51Vgo5qNdlhMVrnnVRi048zKIlV6hjt26L/Nsf0klx7g
u02nFC7ZN+mRBxvZd2AK5w6FIGoxOm0p5wccWAwGc/V+zIlAyDqUozxacLytwMXE
mij8EtuIB0JPX79UTkM8v1LEfIz2ZDsrjxnwYQrvDUJlNw8s+08zSWqG5+UYzz5E
OkAHtmuPk98IU7uRsfzMV9HRCV2cd6f11AnwixuJCgnYs0jKpAoVJ/uQ/9i+mWVF
tK8E6XnK1tPCcRmEgbgpxMqvKCHEgfZQcWbRcLMe9+IIFYOVX7k+sLR+iAxrnvY3
oFb5jdeq7jCkeDPmGF0UCbdOIWVVbnlf+oLsjLcO0VBzjrHh4hUsGpjx3dBL06XA
8KOVAj1d/cynoD1lgMXbVrOL8cJjq2rhbGxra58RsqlpQCax7kw196qU5U0Hy+jg
Ctq9WxiTXRez6i157oNEVhkfZ9iXwEwu9KHXOqEXywxYzZdGzU7ZrqZt3Kj9C4C5
HQ9ZR5VX80Hs1MQpFweczqeQMHksWcj3pxQo/bfw34OIVp5WEtpEGlZQuKA/9jD8
6OCNa9QtzBJedK2rgLQ1+VwzoIOLIph/E4pdqkiQEv7FiOI98XdA02LEpEEeykxu
2loyU6Jr37TlN1a+OO5maVmAiwvKrqu7+eikmcUYTonkO95yGBV4qfk+EdXT9Xks
P2sHL2BdK7RB3vDzZosXU0BDprk0xaS1fQ/PdMqsGwRQuTnt4toBf2P3TchjyrmS
sINn3hHHullHERPiK+RAssVRTd21qvbw3/nf6lpyqWXEbbTqln+zVYWhOFdQ4Vj2
4k4i/k7ycZ+V3cc/Fdk81/3sto2p9C/1LyGn+4Y1HrjwiCiCsR5piJAFqbHNoYus
Olen9fzV+cm3WsCLOdIo7oV4KmPcPAtO90UqdVzyEldIIXKF7ycenis5FepBvS8g
qcQ8hmAHvlaRc+HsF5FIvVpQDPlS8242edRkMPxqvGU7d7CClJxYxOYR4iHxRjwn
W5fBmgAN03wDp4PCMSd2/aa6Sv462g0KDG8i2mT7ltDj8O+kMZRdgi4hvVocL//w
tbvAL5Gw0BNm/qjvsL+iOVX/wBqG1UB6F68Ij+89uBzQy1b04bPoU32kLWuDHGUC
HHzyDoTEGrpZqSw/JHvTnMFaiFOtDxmI1HexComL+VoX1YB0KxGjwt5icOAvbqxo
NpApxBaJS0ejVR1E8XT6UVt8kLE7NrpZznGvLpHPAZplCho/EXrM+JwiBs/Ejjne
SvpfXONwuWLflpmCdCcXwrFzK5HwnL5WwRcivj36n3a8tDl1nqvt+1pLmmf9XeYK
FM5sh5MY04TEqpsHYKbrEr+8B52jYSXWpnefw2i8JvGYdMfH3k4Q3OYKQS0GpAnu
uS5Z8sJwFB90RGG/6CVSzj0wf+InkFdWU8B8pit5DwUgpN/NidVTbifMWporbnYM
K/rEi4oQF4aKdVP+laxAqaoN0sgFlO1h1GJ9xxsTgKr71KAdc4wDxiR6rEl67hU5
JDskj3fy4xe6rHrRSeZUmoL1znqnFAYtsTfp0gFf8HiAzNCHMZj64eM9iz7sbH70
+OBckXzEWaT0S4ORWTw4gD5L9rQc81k8EqV5ikpIoo2U4c4J4bzatnofCEqod0wY
NrWYEtQHOhb6/oxMiZBy+tgmrqhkiJA0uT29bl0BHm9SGMqM208G8OigJpSfRBJE
grEFrIEyWDcDZNn4i8LgGN28020EG32i4c2v5+iqDpbXBn6WF2NjV9PinjW9J8s7
Bfec0pyKLgIWUxsRjR8/5BQ4kLUZdrfRwfq7TziJXinKO6AqcVf5wQllR9n8PIc9
YKCVJtdUS3Sjrv8sM1+CbQijPIqXYQlX0PmckQUzExMRfBu1D9RZui8rlzJIGQPA
FWH6scS3VdmrEbDT6pX8ZohrKSTMj75xXIj889PerjvDWzmacuZ3S+PJgT2AWqj6
uCasNJ06e5a8WTN5tMkBZTJSbYdvT5amWnG4lsS1L5X1+9ML5M/ahqdEi/fmqR4L
5EUBJMa7aolyEU2qmOUlRT+vJb7aLkdWtsJFRfhAQcHvxqk0WWcFSD81suSzzM9T
vIiYn5Mjz1JxKoAWiz5jpn6qxSow+WBNTaOPRAvi/sXTx4AHHS1WeqEAxa8OlsdK
rAroAMP01J5bylg7kPFFCnSdTKs5vq6QsXHF8gpTyMD+siibdjzrbYkiDdVktilK
AZczhqXvXp3ko1eXeG0Akg9oBg4IhcxK+ya0ic6V9nr3rGJU8D7PZbIAWc+2Go5g
53VyP2XmKukZW6Zd6Sk7TbW6TgukgbHCS3JM6VeNKvYjdW4amxMjXMpy/QEsWRSz
gYcAWvD9vCkJqt4KkEGXtOy8mOAmdxQK6qOgYV3P152kT/AqNFmevfF3FNGRRCoJ
j7SvzHwRihEIUPSigp2rf9PEPVdYy458v2y6hLXnfpdaqtLsbWzv4PCeG0O5VIOx
neCwHcKV4VKkrXcKrScdYS+JBt0uRzLceasYJsDUdZ/k2wjBeHM3whQN+T+I+uWx
ac3kVkjp9gevM74GmGjVQ/HRoWLsQy7wqHu1a0okDx/FJiVkTEhKLAW2cAXjRYLU
kTmwM4DOJTZWrnHbzTHKpMYtaO0AN2xcomeZSI2FI1eHwx/jzT+mLb3bjM559NQT
iAIiF8w2t8tXwpwCCwtSGYL93u0BU4JioOvIRBTksMusy0nFsXI4ScT2JuwTszuD
aC3w8yvmzeeTCGciwN30i1BNwKh8avVcm2LY5B6foUW1h93dOuJdVld8HRTQk0U/
Jr2xtwXOuKEzN31vIWy7ZbAOMeuM5Urmra87ebkh4c1QabDd40QIFxRMYjUH879n
GlhdVzh2HGGNeR27oO+ISiWYlLhvPIQwerbOn9+AvcQcu3nXVaOKz60OaBvB7n1a
LQRntyx+bS++hqbsO/pJle3xfT8Jfnt9WvPj/Gbg74zGfVxxlKs3fpoJrwRrQ5SH
UUvVCGny+R8CWWPB76vsipG4M7fne+Y5w+qchuX+uj13ZKd/y3dYJxAnMAeXakRv
BrDv90mGEvbaVr8yLZBwpZLnY1WWla/zGRS+3NKzd4zrNZyoL4gDdCIWlY3UH546
5YOm6i4AdvuvhH4Xlw5HNnGjsUFbwVgLxp0+ONaPBWPn3jRV6LORt8I83Nwm1Haq
Au66CZrxAOEbbigABkTrIkS4DhFw257AXHg6NmgDYx4tAGQ3TPVBQqsz5iVXoGoH
Q9kFHd6n/G/8vrcNhXKsU7SZPb/0fOBw5QmdZE8r9oliu/aZdbS2zfh0JM/hf3Zd
rxVVN2u5OHYT8Su4hnZQxut0uEJU1eW66nUwO44Fv+VjU+/BSG/bQmTuEAHp2HYW
+wczl0lq1q9eXYwDyl6QwpjEeVoCVbUmLwh9oY91sUtnUqLL0fxjMrGmGKtGbGt6
Ffwksk1rdq+aEr8BzyJZY0ZygWKm5soytlbFeh3d7IMzL4JiSVkaH/dxbvo4GCp9
Qil/Ph5fCyqb3K1qeCCBAE2YWhH5c5WLNx6X87ZbONq+fDv8Kgg33NEXyVBOllnY
IUGOWtqnGlGWZ6nTlRF2yHNARBsgQ5Kfmx++sLZsIO3Rn2+MU4ysGLnOY8PBVO/p
GQ7kRrsceFkm4qV0PeE50axl+7geIZquS3MtRtvx1CK7cuUlfBBgPAjQ8I7ittH2
CuYFVfd5x5Lu0oWroXEgBW0uSPHCIAhTTOQOjLHfHY8ZkJDuutffioKQXabO1Y8W
jobZO8T7QalgjcvH9aUygneOH8umMwSvL/35VVWrpvZOMIKTOYxM56XxFj1WNgjO
8D/tcepEUyiterfKMcBDXCS6qVBWBB1KONMlO224gHGMkHhdczaGpf0SePclvSQb
OW8xoMjDS8ZGr8hgvBopNWpYpKKMf+nh7a3Z7E+5aw5qKjJe+fdRt6dwCs57+yhp
lGctq9rr/6fVa1EZ3BUkIuiM7TVWBc7Qcz+bgHocjUuRbbB5NUmAB/Ffs3fbzGr7
AMIYuV9C/HLpjMSuhErW5SeC7pQYCs09YUcjaoCivrWbW6B+wAWALtuNFkdgxBpK
xmxHORZxrkbJRSeIqyFgqeqV+pX8Hm3j0IS1xKHp7Fy6jaBcEwf4WG/NZxat2TMT
ScyXmmBMgH+QsnzpCfbhQg3LDT0oh4e447dI4WoDv2SCAKtRVh/4OevFQddXjaZX
6tWsLxMg0uoXmnV0t2hqN3ISbFBVLrwNCKa343+NAW1iOBFNMG+Ydm8LFG40eqyn
4vNX4kRJbCxvMIUWDv3pAetc5ueiPWWxjh+4gm9oKX+OkYltt2Z1WKARreceXmmK
dqZpvsPN/W1ZTMcQvwUoIWRlJjQayujCKQ8fnM7fAU1+xoxdINOkH7VsuMSAzbJW
n1xB9FSh2Ae9FycWNFVv0sN86197VlTC5TqUruNFG0YpLL0TmwB2F2DmlEf8iAoY
bl6pJZV60yPfYJITIGY+uN7BdfqXmygJOfEN+d5Ze2UKSknD8YpFMwr6e9b9Aygg
ijtJubJtq/XN+FssMcM1t+qEROmTiQXGLGe9AWN29QF39GGnb8DjiOQgqBDdtpWP
OoQunyufB+Y1T5EIZbQGwzXm7q0am6l8i41l8qp2yub3MVNebjJqi45rQNXrLJBf
w5KCe7RwDuiQH4t4Xhwegk0h9azd2ACG77jTO91H8nyVIRuVpTl+jPd9kyi/TMLb
KskbJG1hM1DPKFi/zF7wDjdzh76sOTm7sL06+rH40j537xcxcwYNERGCF+c5EfQc
D5pq3VmU3DET2upjoO2J3pMi5Z76Bm6VdkOhBg8yCfi55v4JOXHAwkfxnNF+5Mq/
DZavzzy4YQ/n5vLm2n0SMOstCdPKnfGDYgEavX31QIG9liXiwk7X4eo1s+uXoXfw
1R8nfNIgZHr2nnwn3YPGvHNZGY4v7nsWSlJ+BJguLoo/H8Q8Qk2teCBzpjC29O8l
8NGDNNFaD7FfzvpJDaeSVrk7Ai3XJBE5Q1pV7h/6q9upPi72DqK0WZm30SQ+Ru85
S7g5z3XwnH43yyPdyMF4j4LLXkpQf5el3pTZp9sPEYAKWXUbmv8RF+dwoz6EiKKT
8qu8JaxHFkrAKdAnBp+1PSfpA1ddzhUvnELbJP8tgyJKMpHs5hh4ZyI7t8tFWhE6
ZFIyq5MrkpgZT7GQWjpVUvgTPzOhW7h62MWC0flI+maqwYG1T+Htv7/pBJD0uvQm
HSBnzBs1fbbSfLAHomFBkEbUIFXZduiuuYQn6ngG/5F6YOqP3HRFIgneORlCK4r6
jpstoeNagDtte3u6nthaITY3tyYfnYbL7HJRmm+kkQUIz6mdUTzfkIaLtC10Vfg+
2RxgdsklVWIhIAdAAvfl1L+eOq4URTjrjYatTHfad0vvlAAYI24MMOSu1bfqFgXW
A3E3rvfS6EFVsKZW4EzvtEE9Dq6R13jklc3oLFpahN6OrRP91L9jfCjz8sscgn9+
dIe3/AGAyPUMpG3h4dbxYYD3jrMO5vL0QhfT5eQvtiuNRRglb2RdzmyFUh8dWB6m
hMMOmduSuHx8zPd1HKTl0YBxcFQTjy0bwNxDRPChWWX42Xm2Qz4VPLfAdunNMuXO
UWru/TI7iDzdlDOgLsIsiMRHt4+I37B53Nv39TKredLbQj5SHs8I5Dn51SA7OW6g
RgbndCZVFPL4gy3dD95RL7bLNCv5C+Te4KT1WLiBar7r5/f5T9cKKOz0yP0K2dvp
Yscqza1ptnRe9IkgNDi1E/SayuiQ6dPI1gOsXaAmPohhKGdtL1FZWxjRiu4ApE+P
Vz1znTX5zIfvKzSxUonBLSUevHVrQiaVX7+ikNS0im7UsMsnTn00szqtWtL2S+cQ
5km20+FZzemT54ZkP2XL9mG48DMu1xmSlxQjueiPxYJknTzZTbieCN+gvf7wYpWw
fcmOtGJYxOV3Az4TN4QwvrBiZI7mYPDDJvZaPsh185lpOALCBYmfVnOEzMJTvMLk
VyESf9MoNNC095Y1qncyM7+Rwl6nRv1ygb+onp+g3hkmbS93YrSiL0NvGLXuUEHx
jpWGCQ4lX4gtrJ5RK/0mAEWAlXTetL8eGvoos4s5fOIk+EAatG1qkmv6rdamFU8T
ryeKDixWw6vpj1+uvIj0me7t94VVlhzfACojcKvhN/N683XbDS2BACqctcq8idns
HZNUo+jZqUxz4b2BOoWrmgUDQNPi7pFNCYVGoPyGuhfxK5dFLMqswqquHKc2sArW
+cvAWCa1nqA1pQSJO3mY6wx2uIKBDL0PWw0z5sQun1OGtoyHLche99s7MZRH2lF+
aY1Io1or7urBz9GIYgxypy7lGct5znEVBbWNLDpmE0aZ0/rLIDAPZzQz56T8LuOS
4eBmupdOt48rQeOnFVdKoShecxTfTgKqzyjzD1dMGbtpnOkxU1Ou8adzgPklffgi
U8IT+8iwmq/mZh4rNILQNySM8fHz6GD2/K4edPkK0KbNj6Cw/yB0rH4mYj7irhpN
2hDCMbWPOC8cwAfQ9egxqxLNgseuNF2QZOWqayLxx36jCdfViJKXh+uYoFZohV61
U4/hCMd72i4jH+fVe5LKEH/kdt9LJBzr2y5nR4pRaHv1v95+mAlJz4CyZc84YkTQ
1icxppCcj3r7GHT4ZFyEs9LScXtd4iYnp3p1NcbzBLVblyhBsW3zMb75+W5bwmyU
4GbtZ9O0c8ZLz6srXLMBle6ScI2Yx/vMxRFvPNucCVaNGovV8qTtvOluYzKQ4EI7
QFp6dEQhBygzJ8LJQJ1bQxWPXbSAeVoBIe6fRGdgWYzcz2vo84RVxPibsF6ypIbG
H69grb/LZi+sipa1o8PIormN/2YNjj0YZqi6GCotTE/UN8Te9325sRDJz0L1WUWA
IgxEIGSQluumJGG8moWlIzi/2a6eacPsVIvLOJPrG/5r3h2n8jBf4bOTgQln+YNF
ZVbfnd9ngoF8D4wxwudZloxA8BfHKsPj1LRv4/vdo63wjIdLIln7FYT8HED8ds4B
xbuPoc9RT+gJiZYRHNrUnzZnDesfxpivV5sicbbXmHnNxd3RKsRabrw8/w35jFw2
B2Y3nDzQzIKq+KNcWBTMBlDELEkNeYCOfZvD5HFhRYcNCYBiuOsvLnrPi9jeqc4C
aQFKPX6GBud/JCRtJgAvAh74/cZpNrjP0nl1Vva6SFtqek8cRixO0KEu/d+OaYBl
QRNEBEEJmNKmtWCmUJYxZ9Mp/MN2JVbelg3lrAcR6/SAgTfqISdFVuVt4SjZ/Fkr
sK3VKr/3vEu3zlKNiPlI44rSwZxjjaVXaDH0rrPsojQnkw7o6fbcGbGNEQT/7NwA
PAiT8zHRpHkFAiyLuvRh14CbVJC6zMbhqotwXGVbLfdLla6ylqUzt7d7lMBViNIW
o9WeR4n0YZm3Au2dUS4mGjT8hiAt85x1KOPdLKEqUSelG6CON5HRZF9jG/XFvIs4
nRc2xo41So+PHGx8GVQok97GJddHQRvED4bNhbd8kchXaF9k2AI6OpDnGzMLXl+Q
jhnO30VZBiP8WWcWsePb1sYmQI5DAB3OYs0RUuhK5mpRSfeTd6/vBJke+LFKlVcL
3KUZ48wgiiTRlDRX2erjM8R2Il47rD/Ml6cctc24UNxY3QuDoCjk2bT7C436Q5YE
Te8LOSE1EYCvii/75ZkBXqGqrZBkqxXp3fAATygNPJjy65cSPFF1ITkDVbqVAj8W
46XmPjw5JoKVy+HtV2yAfA==
`pragma protect end_protected
