`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
OO9eFpk8yc842zWfF2l6b66WwvCSpFPBiiCBba9DfHNE2FmHQdy0vMicw9Rtmj1Z
l4VyN+6HzBT58Tdi0Ua2W83KvXp0urY5YZoaKpyNg7t2kZot6QuEKGCWl5Zpr1lZ
iaVMu4WGc3DTKrPD9KZG2Ebb3Krq77A5OvaFv0HtN+M=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 3200), data_block
txMAM4xx9anlMxUGr8Q8peoFck7eKq1sGXkmSUKr0u7Td46SeoMl2gnjWH+Asbju
3UBb0hqf7ZJeqhsFbcgCiSg4KKHQkvk7sxJ4tqZp7Obhqfg3RSgCWa5f2sH6hStz
tijXBbaWNVa58GogiZQhe2V4HPXE+N7jwx0NdTfCQFnl+Us2Nu0MSbLxekhZDI97
tzaaKt0o451bdVUOGO2VTvTBY6q9xsMQhNqXbFBqsrM+OOJ2hho9GZI870TEyjpU
fIVQiUpT/qH+FkuunQiPlKehMDb8duSVoxoF+lkxJQkVYvN/+OscsLYjTmIIJ2ZS
wsakLeR6fZ8f1gG1lLE1gmNdoM2qNaND58BMD+HbCihMrQj+rHlH6ckD9y/ov2YM
QNLtCrpBZuBrUs4Dw/dNB1IBppSmPhA7keh7KM1gW3nYj8G+LavcOReBql5QqfzW
g8yA3gLOWWjgbtLMidd6GyIm/JZd7WkepKPdVdVTQ5zxer+t+gTWlF0E5B4KtVWk
B4kkJ5kkG4qFYow4oPaMjPBc5wDk1qhbzeldem+WEmv3i6HjRjcmvzk41cugcOY5
QlKDUTrfTP+67e857n6D50RpHFeMcv3aLygelyMcyor+MmzYBfqPZORow0JqJ1TG
dNYjj9PCohSmlYymhC5CXVy9h4Y88P0uRxLR8OfcZT8H7diGL/WSyjDGcyHTCng/
9WfDMmb0IfzMGyKnux/uAFIHSjWCrU2gpYQWp1GdABKlxx4iSM/SzV3B1/iKINNt
iTDaXfv+YOGu9JxhxTQbGu7nXKoqxUY2Ad2rC213g3ca5CTxig7FxBMGCj/WyMRQ
GHHgydK4Pd4GNniohj1fVkXVVwokRSaGd5Uhw+y119oNjDyF/GO3g9gtOGXheclc
zWfXWLLAscfWq7u1KEICAg/XgRFd1mEYA0blHZcf+PQT4rWApLuwIs7MIEupATf0
EGPgpYfygrO9e8bKoOGX0QTUkOFJ16y7PWsnkEbk8sgMvoYQr7QvqxR+2008dD9H
5J5CmoMQEFyyx5z06PkQgVEWCEHtemfogtPytYVlTrUgQ9pJeDcTRg4CgLqFKbkg
sWAo5PmtfWSlG+D5SQ/V4tlRj9j1+mPL6YmWbeCt8h72zNhm6+wcixPf6LBWEFU0
IxF0gwjfRuScWs+L8R2RqN9xWP2/I/LaYw9Cz4c78HkPJel7txC4J5L/3vHboxEZ
CgmPjZCk7l3WZe55ob42IfNwWCBqGWnLPv+/Uk2Z2knw5XxkcbCAMuFMQnHsTaEU
6KbSNhEKkqSnnsfKERjQ5dj54F4WOtNVAZGiq3uWUrmDIxQAIDj5XeoSufAV+MLf
arW1tkz3UHIVLYQM85pOC/C87/nY4HX8fqwZm+F3js7B0TbxYU/keP8daIQSAP+Y
LZ5g1aGCS7lrmZcDJVgf9/HIFQFRuXk+uq/TVxDgJrtr+8RLlJFX5S85858zcWS7
6ZvbKH54v6zxVZZEYG4vkncx5g0XaH44/LvtD+wO6piUAYmIQVN++6wlC7YwEirn
ZTq0Ei539h67/BqZzU6B1crIY5gBUjV+noPdeobUCuvDOG7CmNdcEgmDJT1OYE9m
CTOsUak5LahP1NhynzIC9NyPhlADJEKuoKSTNC/xHqLXHKvuReIPyc5FjT8KG6DM
rdwfhTw20nBq8IXJ95heEx60sZBxVr38YFDkTgcCd5evq+PO+V2hZ2QejeeArczD
wsuD1T8PeOBijMFvLliKX7kI+tdTx5PbmOP8g8RrUnSoZbYoOWHn9I6N6513cgxB
EHwlzhHkksyM4Qo9ZWbwiTzcroVoiNoS22VKHskFIlMTzA/j/oyIwTPC1K5f6X8H
mqwxJDhNMTss12YHu/EXvFjsL07cXCLerzf1K75cRtoaYHEvFif3Jldj9PFr7tiM
v3IWG/ni9KrzePdzzTYBceZ8mqDPrfC0nrFiFB/bk3nwk6tI+7StJ52Koqj3eCDE
Q3xzC23qshV8fZLzkl4/pt1tV6ZklrjyeU+OduKw/15B4+XTh7TIH1FpUtP9HRHp
cRF9/x93FUOhrcijusXMI2f//5bRdx2GhkQbYs1cAgvxKa9oNiZ3g6a/J5C2gOqX
YOYbyf49TQq6YhvrmC2/DWID2UobiGh2skLUKyKFFBgT0JTEVJ6TbsTFWMlo7VkG
Jv/FUnBRUbskoUEp5INAR0tnfTJpQkZSzLgFXvnAqZcaZ9kE/do5GbAZ1G9FM9Tc
HhHRz3a2eIeyqaLsgvwflQqyzjdoaT7c6dGqBmX7DMm1PHD+S0uHVBxyo9AMXWcP
h/1hBjwPiqgWtZaKPgProkMyXJTooR1MO0xYv35juq9cyZhwtmu99eknlSO4RMKx
JABi32tFICaIz9axgtK6EGptCM6RN5UUWuvRs51eQLa0K2DtYqA3Dqz61QywZVs3
KTjWjADPWeRsSDo/usN6hxRe2by1zB550sqTDnDkgPQhUW1epkhFnzNtx3yINC2s
S6IsMiJaLHGm+exq8IBafDIPuPt6XlfCqf5UVXlMyIvcgd0VAO2iree1qUi3cUDD
EaEmnDs4XNCw2+Iv5Sm9wQ2zorLViELbUYmj2hghtIgNnRDIdvr1I/viHtj8nJla
h7OnNhKGhbN7UhKnRknUdsAfgihvAS1klXoud19JwkcjL81Dvn3CVgX/GHcQWu3u
BIL84e+PxMdoSvNbF05ZjpZrXw5EYOyq+7j63eGYh7VE2XSHw98siAb9CUBv7t0R
dNXHvvmHoLMBiGl9X9ajES+LEf46ivUpiv21T2gPgBJVFIcFP00k6DwBI3R8MkFY
knEBO6bAL9fuF9CQUPvTR1nORyLWT3yBpKBnl8skypqOjRfALZCJB8Dpu2lHQE/6
cc35qdAAtqmBoPRA6j1gNQ7ikOZ1rc8qDzoU1I95s3AZgfDcnLtr5sHuez+5sLuM
PiOcI8QixhrOHz6RWft9hbl0qWUbDz5jKRMpGjbF4yMNse+gqQ6PFCrXRqwPldch
xClduvEcLVgtCsvmfgfJSV1QZEYoUVD2ZiWroKCTy8vZzA9+/kGZqeu4ZN/EZ0Ob
LfEcgv98p00vX1fj44jI/tYIwHEWQ8n9M89F30oAjm7jlwBZVYegfEm7nXV/DTzG
qxtLfm18sdrp7D/6/yd9G2YCGvNZBfZZkYtnnUC/n2Fnwi5fgpoRMHT++UEv3P7+
TcIFmPC9Lt/sW+SbSmqWN3I3rHTzRnzidTKllWwbyrIHXra8kFnm0pbxJhf67rl7
pO/a382xACuLe0/Li5sMBRdFiBpUJspk+Qps6B0d5ci5ihcsKPiqwl2l0TL6mW05
NifsPmyp194Hmet9sjQYkzFl3byoh7vBxxcCimM4BKMwBmH3B+Q1mvZKt5NjxDGe
FG2OEYW/VwdrJSQzwlxDL81dlHhWMTGCwN+i0OwhAqz/bBe6AlUOnrphwQbIAKOX
JvbBjtrUi+y2lTFIIEF8xXp03g2perVO//h02w37ncxPQQbncbzyGJYwi5ce41/1
qN8/VqDamqndUv69t0DSY0LqwjyKFf/+nkUr20sPeap1DQIR6BeORZbzWhJrQEXM
ffrQGcCSTI55GgcLTK9ZM1EC2WjaOCX2pYrrQVw9wIPkEFLgJej810cW5yyoOe+g
XyubkOsBbIHgQsfiA2CskdeiZg8/HbST8y+xs1DRntvjpMgrfK4sqfLyTTHe9zi4
HCPyy869IN9Zp+iT6FMNjXowRPoTfvOSd3Vp2DH0eXyD9yhd3+u4pgVb2nw7Z9xD
qvHTlGe/z1jIypK4+WwTSGOoNim4Yk8hiTBj9yM37ez55MKvji2HeM5jYP4eBw2Y
YoMt2bF4CsBkWQSOf6hESQMZ7PR+x2p9ceNU6X1/qRLEgxdKWDXislWJ3mavH5I+
xuzY7lEpR7XRKhEZqIO1Z/BeYRkR//uzgkqrxCTx0jX88pYdbuJadXsPQtSXAJR8
OyQJs8FYmaK8ToCIYLhdGhiHBY9OFKx9LcVrizPkH+OCVfnw6MbzKX4LZd/6LyE4
7gdkAthIW4cLRGT6EQtSVBQ990DLAG+/j3JNgiPeCaw7jQIr/5J1tECzdjka5FPy
8Z8WRYzJ20bfysaUji+FYwDX2zzT87xk0zbyG78ZJTrmBsxcuEtbQ9CbbvvDEAK0
CaoTF8nBgENH+wv1UUBHdCZohX/fW+EThlHbOT2RJplBbpJoI0Vb1eaTgvRYjPyR
jq+ch44t2eIhQpT4iHPHsc1Dq2bS2yiuyNXvo24kqi4=
`pragma protect end_protected
