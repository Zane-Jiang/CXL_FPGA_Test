// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1dsO1v/sng0atBhg2Vwz6yk3FBkAtaSoJpCI0aNME6sKcyO2ZxDsFXbUlJcbHcS2
Bb6xcm24GOsEgWbhe93yVORoeAsJh87GeJxCLEr/MG2efUSuxYEXKLMjKUgr60b5
/aKzHTUlTK4qFraadhzvo9dT+6TjlqT4BAuKKwfkyYY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8768 )
`pragma protect data_block
Vk6KvvEZin8hbCwpGr+7Ev4Hn+KD+X9Sm0Ija4IkWjfag9szr7YU4SVeXR1Gx86C
vM0ev36R2jDxtqx8wbN2IfutgbOBMKnWoX3rC3IRZg68cr8q67od0wfPpZjwAg0+
LOgF1UMpY6HoHBtzwCheIBI/sz0Z+jjMPFVT7N5/+jRf/KXNp2sYu4xY2zeiq75g
Nlp+XPN/iD35pe22B6uLAGHaX8c+2htRdaMe3cGxlCtII/Hr2KBxaDpvNir39UHO
LibLGv+NOLxrKS8Au2RtUQLdk1dhn0PXiSOwbaxdTed4sVyWAeRcJSeDMfK2iPsz
og9iz2wzcZ0xFtDLgHqbNs5AWGM8Wf4slEWzphYfjFhlHZNZSUisTtaClw6UzdTf
vJLyKi8Ocac33uEL8e9VGAjeYMXGdy8EB9gPRX5JUEKEkqXukZfPM8kD1QfH8dt/
zOc4kTzEd6WKoBUfO2Len1lBa+G0PlMqb69McM3ao3IFX3/48BpTJwjwkiO6nHIK
I/HQg0UXhF3a4tcJry9P6AAT8x8yMJvaEUfTkPda2XvGs0GU3IFtTnGUQRzvy0D3
xUVPRV2Miwk2WqpD67SpOssrr8sp8WJHCpOwqhQPA8rCyMjbFTg0gd/JPGt124OR
hs6PSfSS/DWsRi/wgplfqz61LhBZ0L+2VmMyjTYV6wFkoLUSQVrWitZ8O8xVgqjt
RZLKc/iS54/NGrSp0tVBl+Y9WFNeJha4FZmBFGknxdPR+u1trRPHPk9hwbWJNtLc
g5JMqLWJEj/+gNc3H7pvKbuVWO7XiyIOJlj4CobZoookqt+1gzX6ALNyfYuJwYEG
5lKDI9aKUfIhkGcJV0D4g32X76BcDuBtpe6Qfh6s/IU0eNoHD9RUsyR0GpCLc7NH
TXnyPc4DYfSdGNteyXAG/vNPKdeh/p0iN99wB+Qk6++C6Pq44Yj7JvkHsCBnx2wI
nSl4mbnpTVUa6YJfHpwGr/R66hYjjuABWwuEI/R/Mh59JhhrzYGDmZaJ7hcq2B+e
HPFK4v0R7CrtZujSVUKvgkYk1M2hnMIWkqyq7qHKHwcTIdvvSXbmC1ozRT+RMHQs
PIy0THvyamI1YBBFFRle8IjkGPbfn/9SM2VcK2qwJULV+R/HE8II++KwJ7E2Spu5
q4kzbq2WcIpaBG1rTJ1XFUiEZNCpg8xQgY+PW2HP3RkB9Udyk9FP/uMnFSkRPWLR
O1b8CTmS7YO9NUPLlCGQhYrCLjQZgvkpESbWqc4vmNzge/ldecKcEHcCzgamKonh
c5rAnH2F7HInAial5w/zRzpK6xOfOuH+iOR+9RIhf8P0U4NHKWEBkH6ODsNJdrWM
hpuwdq7UDN//annN26neTlcMGz7lqKK+qiBOsr3Lw5GPZhJOyLB6+wo4rQD6F8Ag
/bRYObOgDstsA7cq4ORflsZkj36xLBKnvVAv8oyxVp+/rqO9kV7HBMVDKk0H9R4q
2VjArc7tZeqlW+AV0d9kA4XSTSWiDRX5HXevrsQYaRmh6Ok87ZEbeK3HFngQxJ/Q
zZO5mvWt3e89vjxAdRiOiJTvQtHpAxRlyujyfpz4+6wAyId2Cizniuct8Hjj1Etk
Wwbjk34iEihFprTEXH9EfHBvPrBZLlUj5AunnwufCwAwcJDCvFzPloLZR5brqxF/
nUqtQtDuBLuIe2tZpxbT2yflECfAbSwQugqSlv3Ems9vlEO+zfjDQSbj43AjvV0v
SONBTy7Pg8WicxjTQWoXPk2oYfBU2MSVrq8efFmrpU0mn2OMjHe/fw4jSIwl9oxU
88IS2q+yIDMoRo9VY2hweveIb0jNRWONHD45p8OnmDCaTE4Cr2vuSzLkfJ84D3Oy
Y6Wk7IOSlk5m2Gfkl5gcKwJ0rYDQtrmWF8iAtIHaPwC/VOd536bttsjlwV6fnZEb
RJVmCPkRMdAkDV/7s8I6Kg8G2jIUTPa+qurBclmtfnjiN12ImMH7ROmj9/2dnYfz
luvtJmINanIrj77qw9c0Z438gEGb9t/ekLKLOv4RXLhjvPIAi1UI3elOazQC8kTt
4zUvHQ01o60yoGN0vdyXQKNfZmhn75C8stIXU8TmCfMKV/w2lyoFaN6rcIsq7RjE
33Na0u3VD/oOJLo2CDXAi4D7J1LHR+ppzj/z/ghFKAtQjARs5nHRkOE+Lpew0INj
Bw51Db+y0etgtIyJZEtnSRoAd2VjVDTPatp523aSIan5a0T+ebTT5DKY+Bml5fcy
kzTaKikYe5A4XoEfQ2QjbR97Gmk7y2z3Z9CXqmPJQcjG29npw9dHsPeH1+sAn1X6
3QlAthFboXnQnPQZIjFEf0xukFGw5xUP0QcsdO4VmFl1jSmH54Auwa8ZBjaMoxP9
ouEp3cuKzEqc+m1wpNuNFq62CyqolkRJVVWQUuHCOts6mHBP8rhpjMq+f7g+5L4Q
YPfzUaTU/1bhTd0yoKM0ZVItbZF5oRo0mbjvI8yHoFb+A2KTrX+nE69mjb/eGLMz
krUrfWIRFSpomQcF9KBhD975PfnGnIexejRm97SpUtt2O/HLi2QvhCFF2jn6Q4zb
Akjn5ya4/eXeNQafz8u9/db3x3Yc6/H0KxxH8e4yLjGc1DIYffhU6keW1J0L0jiv
IInSfj2pdCRKB8wyAdrWeuKabAwPwqJ98crH9R3vWjxtY0KaH4s5Npl3A1fAQd0z
VXD2fWjYXGLfS8i2PIQP+I4WsrJ2p1ICr8t8Bt65TGoixRGD5vhmZ38mJ8AafBhk
0qifpQYEsUVnWCDsTkDsMZvBuOuqALsaGjIyCvL/S+lR387jVNHZm69E3c+aUU2A
CQLvpi+e5TBjfXg1hvHPJi+lFVb/xu8qMi3IKfBcsF+mrQgEzrpZf5Epj9iM7nkN
1pWPATFnkBP/48xiU463ki5tf1PIv3KwlEzjPHo95HEp25T0hflGc5LSIzss3GT4
+MCT7qQctwmqiagHRUV0npI9GVVbWZXFn1q+0QzHBJVwi4qKggIbgzw1YVlc43Xb
i3OKJT3s7ZGSNh+k9Ba3O6wToGshbidM+4jk4kq1w7+prPRdLPlrWAI3kGbUTCWf
sAebnZnBbq5YbW7dhX9ZeUpDxao/SNzL+6KY/cN2cu6nHStQgZJ6hqvw+4erv2AY
e6z95rjez6XEpjTflKjPdAbOZmaKHOuPeQLJZ85XQzGlfBkkexxwTSE7E7AKCi5x
5TPeT/vjsKPM8zowLEp4VRDJKxsRpkmydapKeSwcLFaIHH5hiErhZjNYCYC5g6Ba
dDOaGZ0RRiEwl0WFFQOw9G0pCU9Tto7MZvMrKWn97MZyVB4m4U+0fkc5rOSvmGQr
NXAbaNfsvCdrMlHt0bXuwz0QQdvCWfwcgDK31bKBFN9hgOSg9CrA1xu7VzNJTS2y
fxkX0wB9/TO73ysk1Kji4Aqt4AY/x5CHQycn+ZFHwyquAWulrZYZSmJ2WCjLaI/L
DyXy+Bue8sINx816NCGtw0zg6J0wdw0mXrp1DeP9h2ctfgEufUl3rWqCi4/Gr2T1
gi3lsEZpvheUybDv1LKI+AvU64mVheqT78E5RXiqY7KPQKkYHZEjZu4SPCg/wBKR
5WsqKeM4v3YVqmSWdp+yL2PgTRoeuYdjVPPVlaTHe0AyrfZHJYKZE5/s/t8Vpai1
pKSSs7+60eNaWAcWnAnPHDvu6Tc9rNOwlsRkGef+oolmNfHONmMYTabFwMZdEHC8
aXZT3TVRJCgJqCghDzVs4v1hwRSOxdTbvL85dxtRdBqhOm7Sqcd+SMx1vDgFK9uw
7+n97nG0/AH9QHVRV/JMdJ8ltXE4mUNfo/rWCPor4RXQxpoZpGmswjxK7RNxWpSA
jcpO6d3ZCS3cXTxuqqGBKAGLlQ7QXhH5XXSH7xSJEqsGAT0gTCQUgPpKfDGvoiK9
J3cNTx/ibWSqmlb7U5B8RviSF5GQm9ulg12KQ+2y9caf/Q2n/WG25rG4GNsiIHzP
V7zr/FJE6fX41uJdj619LJHINLxhH14h6bAJGaxQwrxRMdg6uK1rPvHcth3KtaGw
yCgfch/lqr7Jfd26UYCiJg+s9ZO85BZj3HQdt4WUaZpMgcK3AevWB6regDTMKbxC
v5lqYUMd2WLfunElzVPRMA5QG4HcgAdfK3Z+nv18txJ1Fu24XrL/nS63qN+wUqVN
hgq1IBUUBP/85rQyKIajrXs/aPv8zkuykQdZL9excM+/pjsJq+SD2O55jkrramtF
h0oEC7/PZmvFeAg82Te+lBLXBnBLr0ukeH/NnDMgzWlDanb51wKQqzoQleAmV+fe
wZ+FwAqCvOu7UeCYgu+SpCxahXno+kieuRG8u/m0PdRbfk0oY/Wyc4x/XkppnmPa
NNIqhPUt1fe7ixGXJ5+FftW8XMM8Bo7as6ppfuHkcqhFHKjs7HV9+PNezJy8I/hr
3y21FgNx/N4dUudcK3MBNwBDYoiTTjMfWcrFzIdvFK0j2MGR61EtctRWRrM4V4Vc
3esCmvKll8g3HFsl9Er7yZLhlM4E9gKSeGmbI2jQskWo6LVYYjxRfqr1pGT4EpiA
CLm9wMBwsBdqfudF7Hq0yxxygMDyaPEl/KPTgMZ0SdFWuQaDVHFP9ywU9skdo/0k
iig511cvEnj3GNA2ZBmpF/exaXE3pfmlLEKYNIZVta1WJK0gmSBtaScWJArnumIz
1LGqY5MAuDB0RRdGjjCGzZ3sQf3xgYXH2SJq1l1snc7cMbPMUPnosHRQUQquv5/2
2WP8wD5utk9BC2UmfWoGGPosMrbAhtUAadJ34ff7WPeKBrAa8Su/dudV4iEV+iQf
NYmBGhnLdGR0HvHUfcDytEKRJ6l+wJbSDIdXruX2/g2PWo5ngPCg3l2X0LiiOn89
hMIoxafminRncFBLeMPpnj3dZJyzamgGmbajspX6cedNaQcxa+bq1G1Ja+SGvqeB
6KYXa3bgvIOmiXI00KnuxvTbwUHLDPDcgqguhIGu0rWJivZpNYLfAPH9vhFqDA5X
0uO+bgVFEWJJES3AbMeZzDSqJq4aJewDd+otmnVs361SUqW3LMVlj3+YK5WfaRa6
uu2KiuFqWnveFU5XUa60fKjWDVVwkTLDGBpc3TDyes9UGvSyyPqXo2pZm08q2fNv
0sr8DqAHkY5GO9jK+QDU8pVkPUY4b2EQzZB4D0D+xNpfCj3Jjj+8rS5BVqPS1x/L
+mg7ci0+isGRrv3H9jjPeZq+t9LDC6SN0Z3W9QuNF1n0hZjZTLE59koaNi0Ia+Ey
Tv8DLPzLBAg9fj+UpPw7A3LO0VMkVTF5fMow+wvKkHtHNX2yVRHX2d31HvONXEqj
7Fe+XfczHVNDVUTwhhBDJgJ28zxapM19fdllyKV6l9ukVGQ40Z6PhmCglqSOF5G6
TZWhBw0YKW/Oge3SoO7jvd/w5qYAWBu7tCAWVthGqU3w/XIf+U0i7AcJ5x/IwZl9
Yiau4MzjTWeL/N3jYXOgPszyIkjU5mCi7txj/3XQEysqIBKCvcETLaks8L2IkcKI
2Cw2CcM4JR3eicCdbeb5P3bPVBU34PbYPd/Kt7A4yVUWPADyLKKmJVhNYdx7s9i/
bQAwLmxUPYBWE9+ZUbAMDNgPNc+zVbdX7jNNbOwlnd2K9QHbfPZnmi96hYX6DF86
YV38akfudXlztmje0ea5vqwPqM3OiOTBuYcC7jptbIHwZChPGkNUfPW1n9ljIZ5N
CAxJQrtEZsk5gzTP7bczbdXqOpXqq11q1K2VEW7G4xunAxVGnEDxtrBK1GbuBpVa
u09uvdmMx8OLC5euzWwDd4sjizU0Qysv+k0jXv98Ua1ZRVxCFgTDAMULY1sKVSvs
IhzfodY+OnSWg8M6dCuFOopIPbVkOVNCh9aT7vKV1guE5I4T/i7R/PsQ2ZpHubQJ
PGMi7telnf+5MQxvF3ot316HDB7Vk29YlnMZB+wwB6+5+deFUyrUE6x98gxZvQOh
YAlvsKGxJBCDJEFMDU2owJxAqVDbEn0TFCd+JEZHBAl0D+iqlwFNofrUJcEKC4sE
bfz0w8p4G3/96e6/QhBodPgrF+2B1RvFNaETK7I7SONw6M7ngRPfEPyXuIVkQn8p
Ibso4kTQp9I8VeujxOVumhRVvkpyDYHXm7wtVTTHI7GXGIKDCE1Y3nPUxur7XRg4
Ye5rO9AMTTnUOcnybQnfrggtOGNcb8a0sN3RU4XQ8sQO/+Ytb1OwwJwvvHHg8aFi
bfomTA4jkitzEttBUFG0sKpoM4Yiq5+a2UZGX01pwY1SILFXCJvo8/OlTzCWZghj
DjrJNM9DTe82EDvVYss9/e3b408okUVHTN+GuNNKl7aykkbUf0ZeWIdfkJS/EeuB
mzwh/1Wo0EYwXGtIsiKzuxwCrJpgP3aGFvtkOALhZob6vS3CV4XsmQUuv+CvuxuL
9+LCcBE50W0QdUJ1BPJ6DZ0Gw65utl3BuDnIXhAgA3039EW6lruA7i/1nDKCJfyQ
iDofNDkek22fKJ4OQ5wRdWngB8t6J+5rbbFEwdrnQK2+7s69Z/MHqQaw0I0+RLPb
BE+WGV9iyGFKWc9qS0dP/g2BhEsp7YAtcTLsSylLb4+PGEIXs+vbJ+EVV0JiRfBN
VwkWDescbO85k388VIuNos12gvGorQCazRnESzPtfqDncktzdD6/RtLrePm856lq
+yDiqmF7YnUhO3ucvLvL5kFRZfyKqo4GVTysd3/FJB/tFha2ThBHLks57y0EP8CR
MV5sI31EQYliRM6kV1CXgkbiScds0V17qzXbDSm+dADj9yVi++ZY6Ag4i3U4BtYq
9MEM+Q07TQ3xRiVqk81wOH5qsT+2rXi3x2IHIS+HxsCCroPveVcELVlV8DyWuyD9
wWOYq3AnKutQk7Nn3iv4nu8QyJLUhm4MNLhy1AmJN6BwIs6STBsyw0Z7Yt3PuGvX
pPPk+B9ctumzTXas9w2vahxvWrT8Zn3DFqrYEfuqZ1YtOgaZZocxXQhgj2lF+PqR
Qyro4Ty/18uRgNsyXNK67ZP/Gs3vCXBz32+JLtYZAqIsa0/V5c/tRXqsairXLSMK
iwv11M47ucjevTMxSMLrdSBZl4omR5FWUwb6s7ETCeuNt7CbLU3tEbNbtSL9mgqa
KmXIoZGohXkW5RBit+8o0HIoBS8m6qddrZAJ5OnXRZKgtkrZWTn/kOqD0kSer//Z
2PguWNZHa0ygH7ICDRKimhm9H0gEYX0Fd5SRAT+b9dJvaLDxhjDaLHGtWTDA7ssG
sLUpkjkIZgMZsor0uxgDPxtBmlHnvQ+Ei0kkmQufrVg0kIGtJU7R/KLA+IsRZsNV
H9DQH1qpT6OqbuQk1j01kooD6IZ8j3FxoSvA0y5ot0pJ6sbLH11ST1+LjrQNGRlY
SqDvQbMbgXd8bCaYAw7+V8e3YXctROQdZtsRnRNzwshn24Iqzz8GzEJGFX6RdwDH
yE/ufnR0ZErii89I584hGugALgSsZOQknNuqNHBBjLct9TfnvGeFPC1Ai4iyye4+
Pk8wjcTJEBgZbt3td/WK7dRiA3IGpHGFdNvcnIqX+iHTCBBWgW7o9vnOGcm+kCNJ
KX2/pW8pOUFGisv+AEW5nho9f8/duiE0nkGFBajDMf0Avij5ySaBbXjfqeOYzCFO
qdaStQqQkGA5JmAzfRaoF+Kr02Ldx7R4VkF6k3zMbSYD81sM0dpQNnAkQW8TPadM
irXYlEWNIP5vdt8AMjvtfwqvrhtbJNs38BX8hpbkgTwIwq32h071PzYMMqe+gRhg
MQ67VRJPvE9bV09g/Haqtc8/PVjndVrCWyWMAwaFFZn53FUIR5Ka7cloacmdQ5PX
A/kgyC59lCco0u8eYUvkV+8OpmHgtLi/Fo/nhr3lL0Fqg5jTM8x3znCIKQDGo4tR
FymkY0zEQKGE1fwi99yqmqAtF0Q6h6InYj2eOJ4eVaP7a+7uBP1061UVt74Ux35M
iOU9vBNmL/yuGwQ9GQMbTQDtxdsrsEadnjnMQ98eFpk2rb029jbP3NREwAVGouCS
k6DW95p72e62sD+2Bnq8Q5pg45TLF14vnjYYhiefZka4pzk2dMcRfBwhDsmdMAZV
iwOXdOcjbDwqTzD4ZbyI1CTDmfH03KS7rBxRn/umISfTmyb49HStaeLeFD1jMtPu
RB33t7Oevydc/YGKpRwjTCj+S7agQqqKATXnuIQ9iOieBlc82tZTyx6YO2v84OTE
G81qLonOdVQpa1dK4FXmrHbDApVfIuScpUnD2siv4IJtagcruGwswRGUYndbWPU5
NDYGQJGZULfrpeeCoh+4pJfInPoFV5FlyEtMF1vfhLX1tDj+Pn6hq3c/uWGumkcV
Gno+axU6pm1XRIFlkIO7hd8u7k/UUWhgRRl8rEUwOg6c1DLfI9m4VIldx2ZF2jJ8
mgNwyLQYulLprXAXvhB/TpAXt7I6WjZC7E6JDrNI7fjncH4bGvieC7WTFvrBSQTT
k7EIJKC04wajjTnyjy/HrKxl2NzUG4FWsLDCgBM1H7NG1G9AiqfliDltpp8QP+Z+
ofvdw9AOhGd93F3GJ5W+d+JHil3ybod30d81r9k5ti+yM4n09rZ58qY3b3EdVzxN
mZVdFXXYHdc0ydYU5Yc2YgxpRvexehIjP8OSaZXY3O5+9sl5aVC0L5bdm5qDSLFg
n/3j8LTaFgwHGImIQQJtRcpZD4wk5hFKEATGZ9M4+pf8eKVaoWFZexhRXQO6Yhmr
kDMwJPR5xb9ABPVVQYVhewi0l4rr+SCfMyXWMwpVQ5pr9Wgl5UCMaK9CSu69ndHQ
/fE3F9K4mE319+YIUfd1EHp/gDZhohz/oCVNJzyFIJWlp0cXZCizVPkG8rfEupXh
6XfTAwprbKNca7nNVwi76uzuD+iF+HR84RRmPvqZta8Fvz38KQsEm5rX7Pe+IVfL
d3MAs1UcRzILRz0dLY2AF5ty99l4I+Fdu1dLJj+ghupqrzfPB+OCWOZ1BmOB3Mu5
bQE5E9EA48eR9cICNxhr43lyw9y8PgPGikOgu0zi79CeoZ/bdSx9BY7vWcPWPTky
8ZS5k+oaPCFJoq8MFRczcy/bYqGtV4MpaJHRc4lWTQEo19avpeIMWa/bRxBOR25R
aRLx5dM1M8An4nzITBQFKGzNEMr1y94rIqNXOY7NLrvRWo3qhg69LL0dJs/9TyhB
jdkAgwKNAdpFalWzrhcg6f5uYYzgrhULI3IlMwDJDPa+/wz/jUF+i66xKRqsvgfi
DeLO/f+TS2TwR9LwkO1gRUqSqlfDK7iOkp8HaM7QS2fhbjjWrHR0qJq6I3dTYuwb
EJ1bUIPimTzJ8BYawMmY59+krqBLKDtCnEL+Rv0SHBD4saxvaF+7ZhP6gtzbmI/y
QvtjF564FZi3cHaqlmVFucM+bUcO4A7M5D5VK2sqMYRqXYbtxKBb6zfpcrBPuSmf
Q83ma/tyuxmUNPRN11RqjGQ4+SRIHVYpcIZP00edZkyP30UrDuyI3DFNj1sEJCRp
+dRDU3YnJF0Udx2xqtV54uvL3zjJ74QwEsFWBiDfVLh111wIcEy7UKIfnxYBxgQW
r1hFABTFp2zQ0usaClHMw7qeX0RvCZMv6+D/lCUyN6vpnSFWWj+chBuF929PtKg/
8Um+7p+YoMMpNOnUkhro+fTxAFA4mVfL1poMfDNHHPYDhpkD1TLC+IcwSxuJxqSZ
OVFScZok6zKjrI39QIUM2pbCtE4hRsHrIkYi/qTrlOkfMQYfV3XvRI+O6U9ZEAEE
pFfKsvQvYhCoy5cEjV0GgbRE1P7KUquM2Zk/noF2T4xYCFKuDpI/VicsPejs2cB3
azoC7IPdhhZsa3DhzVLxzy2FfBReXl14uMi8A9fFgb3uz9k/dzG5S96fPhJhZYWB
DoTzVamtEAfZMC9ThT3j5urc2IY3uUG2JOWP+9UtPMnTxKlSS+c/5ml0IwjAPkR8
QH/RO9XyOONaKHzsQ3wmbvIF5P2kXQRex73Q1zK1y1JcCxH5+PAcVaIzUzF1r/HP
E8JZLRRFUroVJO7HjZ4mXFH55ntzkRewFH/KjZsTFU5jHlXaaxzVoX7tA9gw3bQ7
rcB5HPsJqEAZHcbrxHSseNPSkuydEXDVq3qh1pPbxvSF2F5TzF4bK8FIq6G9Vz8+
aGQOO4sB4Le9JV22au0wyfulzhZoIvDH1gLQHnZ9PCG4NHqGHY1YI6s6e/KWmQDF
MuR3nEBWjaxRGYp9ko1+sCK2PRRcYLDAN2PgOPhi+uNMCm9+cRzE29JBwS117S7n
WFK82LhRU9Lr2GcKAmeIRSUXFcaJvS9hFaQZ3OHMiVIke79cdgs7a0izdBbSPHuJ
8pSEkv3lS0PReunIUPqw8jokgKkREe69RBovAkDK/U57cwCi8J7iSJ5HhPp14uiL
H45E4d03gcOYyEhK/AeteS7iOcu1TjGA7Pgs7/uDXhlQNKG/MFgw+pfvChIHMuzD
yyHvMtup2CB6UU2fGr3f/xpZJ0bhr0SdLoGcLN8sK1iQ6RACqvst1YBZhs7Ml4il
dwtKSpLhB8sFgtJq4aYX+Ai11wjkblGNqz4smcC9pakoX1Aw9vzqTwFipzgqMupb
ZomuO01pvLAxKGvruCbRavi82W13sI58erKoWYuuuvpuyY3opegWzSorkAvqNXFb
NOQDjD2xc9zn81nu6tQ2K25712Xw1AIOP9Ub1JQSzdCCatKFZ+6/1bIcnM/5jIoh
90tiLsODmh/BsxJUmEq3Qv17P4OMacJxL7aK1FJOS0l0prwxqpSBSrBdYOp/nMnk
j1gljR+U8+9w8zR9vMwtf/R0km77VSLLgWzWxzUtb9Xgtu4Zaqas2wLq2Uz8yTB7
3jO+cizeKJbUeFWf2zDm1jBCkBmfu514s83yhxgO7dlYql6ARIrueRvVOsH4JPUf
Nh2GsOuzEs+cufr6WlZxpB0dChoKBHEngUqaQgCk1Q8PlK2YAiI5Tr6qt/xz3a0g
Nsm+9HWT7d5pkTa4monH6Q19Ga7d/JSP2b1BXZ2kxk3+IZA4+/RVIuB+nfOgMJ6H
3u52DkuEheeT+llAL9es05AYsJK7+FYkoRIOibjI5t91Uq+tUiexY0ANmo/QRHeC
CGx+31xQbWulOgVRCgw2M74dEtgMTB8HIAuRUgL0n8VYwmvGBOO5ucXbIn43SCwu
4q7onstJfuik9Izxhyo+hMt2F6Ey9A53gr9zUEaESBpdZStnhLaF686Xhw4K+zmv
I+L5+Rl24GbtIReNx3vqusomDzRIS65WNRKpxbaVzK54Xw/YEklqtvyP8OYziK0D
KtzOi99cEZ2e+AK9fTDQI/fD1xYpt0ZX6ccFFMAJ0jSWRL5FnZVy1CsA2DB4IfV7
bKAMT1RrLiZ4paMUtNPlxeDeD4wxr3HCViOAY4C4VZpAOsU9eD4u63Ssgh2dXf5Z
CztOm5m3hKzKz87lrlhBHicu0xLPhkMtlRKGIJsMONVzt18ISbOj6Q7/yom/lOis
R7ZGbWeIDnng/5dPHKMQ4/FWH6wMnHCFYC/DA1ZFdUOjOHkkl47GSqrDDWYP4YBz
0ZBxq0LomGfN1a/D/qlzWiGYcUQKM5ZZECKLMwzRD/Z+Q2ueTTyBbjXjZY2c+L+/
GfBLiNwDEqGzEv3BvEd5bY616+KN5N7wpnogXk6Ft4SYaO7dMF+Ueu2x3U93vlfO
JUIAKviPP9BlGMlA3KylzOMo34OuAkhMlmAlrl+zdZw=

`pragma protect end_protected
