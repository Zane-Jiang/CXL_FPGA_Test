// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h7mXK/qnBsCAVOv27e6XTKCu6xi/kMlguINo3TYffACur7uJaTzGG1ZRUhGV
7xYbCO+iDW4NUtuv/d1NaqBCzNh1QXMJmnqWUIWmqBHZrSgTn/xA6vSgGRon
kIGQHqZMF9/KtuHhK+QGJxZlIIW7ieLvYS5/SgLdvfc27hwc278xBlYLQdNB
A2XWsujardzN8CcL9l0g0Z0TDVXm9OJWYuJVau6PbA9dzHG/NhsLI9+XeGXh
QkpKhAA+DafvGgqZmOoWC2lheYZi7y6jm6AFyKVVd2yF/HgoTZFfyO5zLjeC
CZPuUHRL/Ie/Ya4OrZn0wHmaDztDByAXqCA3wkeXfw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VLw0xTw/3WTvkr8byYwBRXSIlSn69N7Aw9Se9EIQ5H5G3++3u6vvJDljEd9x
4pcw/afXQxzuTJ/yc/EDqhCffso9WL9VfPNuAHftBo7wdO14E7hdQJnJ/lFU
DugzFltQDR2ld5qtAQnM9aobYit0jn+kV7KYPVGN1w04qT3JtS3JuKlK3Hh/
YdJo6dAJ0feQfjnH9LS8ZyH5sWJ2lJqfp9FB+KUzpp3lprFwfpT+JWHdNeK6
OCdgvw7cWvCNYPFSq21fXekVLkUL3YcbO/VAGpsCEe/ZldRoIl/cgD/nA7FL
5SGE0X3cmGK+S+ZpcgMJnu+7Xik8RUaJsy3t75i6tg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZQT0xiE5/dJNFZRpU/UqZ2mbeciXj/mXWH6XOHp0ryU0uEVKgzal3GG3dVQQ
umL0aHVOHlo5zDwZhqgJYLZtmfV6uL/7PF/MCzfPW9okRTgBn/GqkeUohd8x
oJYoVhcjDjazPYA08yJbTH41yiqmhSsbrOqheZdkRTNOXl8Z/xdWQfQlPnOh
cCRLoWk3oLEHsCFY00UJZAMpCbUnBAIKRrd2H/LBeSnvJXpltWbYCnS3k7oQ
GWq/fhRohBfC3qvRbfNNo9VxnHm2K+kk0wLJ+znk6LBME1k53st9I3CuUxqP
IPAF10CFcfF0kiSHAkQ1W4V7Xb0x+Zq2kjQlBgguYQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qVT9E7Z5zU/z6PgdAlcGgWXbDzvhn6/d8GhCrMkKGSvh21rGqsY7ZhvXJu+j
TJVE/TcX56SUlrAlx1oaukjDW4vZHwhciq3jgo46O45ATxSB41I/T09fOn6w
AyWPfBw4/hrQ+EmgOuBs4Y3xUMVBcAVwEbxUo8C42oArKOuTXGQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Gapvxq9ndbS8yoaxVpIXjQFylZJFMAIs+ZD4GS6JFBg8gmhWE9mDwLAmAHJd
BVUVX7GyXZOPX6vbV1D5CauXL9Q4d29F28JdTaax3HC2DDPo8vER8zuxFRuW
eBkHZAi/cDLKK1TTN2PBRgTDF9vX6QMpkdPgOyJo+2QWzyZ5WB1CFnidtz94
8UoKRmaIYCReNxqOToUn7saQDMEjJv63HJPVIjflr7pw5Lfjv7Mq82oWwV78
5oLSq+XBKBDT3NeSMsRDdEPwi8Md/XyGJWlMyQO0yVX+JDwtd8TeMS2YVb2t
YF03C0MTWU/YNy24qVzSY/1QL2I9ePEoDT+n/xAZbNAJshaFgTbkl8noTAcB
4m8S7HZ6nQIHMaEeFtwvX9gcE1Y3QiZZlOq/gbYnWwJ2fm/jA/4LfWFKNzhF
lbTp/FkzTjVNIWx/NcoZ3rrQy8leEIqOO+LFPskdodSi3Q1TRh5jM4N0gdqI
ZZhyx2slJ6LH5QJWg6o7Ahxo+qvnaZG8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k8ouN8hgzz/cry9X5kZbIPjtFIdKHXQYnUxtqV2h6nLsEHnvQhuHyCdPPgaV
twZmD/VmduXOFT92T2dtEuoBu7fnBnAhlZj3TxHyP13NOd8ak4CQzBO0jwut
RF7L+77WMkw//M5s99aqrkqIM4F14hIBN3TsEgACX0WoQxzs78w=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MYmLLkRk8nla9sOdbZrL+zMqbAwjKr5Ff+XNFO9bdAQyNgFTAbtTsFMkPMaA
2jb1I8m/ssVnvdMyIJVNrHQn52RLiIhDDcFWIqPFZSTFxkwOwmyL02BOH2SS
SWu6mp6mmzVasmXtklYS1J2DDxilei5TcZI4vtuS+Q/S6T0DpQw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 976)
`pragma protect data_block
wj24A2kVNg1iWnI0eIwZvyLoRcU7HMoUQQThP4Ky+cKA8HKv9WFuoIs0rjtz
Mk1VraAYDS3noHTkMO22cf+F1CuISoqe/46a47vMJ9yeWW5VOyQDW3bi3+EF
zAXfhtjKtWKQTK2o5qjHEcOc0dHZD+6x5OER0iJYa8cr1X3Yhnm18xK77HcU
tUScSJj5MuvVxE1oNBfsNd0pSpzYP2Uqj6P2D73sCfHnWf7rlzQ9uBQJZkAN
wKsBQGR7WrMTVwYBBuj8gilZwoC1Y/YFjgExhW7zJAWO+zDlHYWVlGQIdZ80
U96vQiqCY/gWXINTuP9R+IcUVnm6j1i75KyHg/V0e8gG1kNUmLtRf8N2dUSf
xDBydwHJpls0EjjpDz1kD3wsIsunTjL/wczKZd8vWFMiwIUgNyT5poPFsBQa
tIZEiSSKgDA0OBWlPd7P2yEtdoLw3gHMuRtlQ1N0ew3coHBcmbEdwqLGtnr8
pjNbc4BYO1UYZMRcOVpZxyTKPlLqExBMpvx+5T1IFwSAdzA3B6uevv2E05xN
C5rcC9E2Uii1z0E76EY2hJn16pPd82DirNogS3ZwduRgK5dnIDaLFJC8tB1G
iXZ44T7yN9Jm5rdj88ToGIeQ4SWIPWOUnyuPD8Sh8MvCoctb/lEqQhPAEU5n
/rJh3FfQ+XyYLGoB9Rp44CwPNVSDs+lhWmCTTrUeLcWCs5bxJe3xzlGPo9CB
QvUwVFMVPYC0amBWMdTcoAMpy+xaEjX2+LazQ/GLSSi6EIuYMEf5MUEObuWS
2clbJ5ZQr3CCB+PM5eFdR0MiR8rW27caAsPXl2IPz0eZHZyZlju6jwiz9oNQ
6yoeGxyEQH06ERCWguKnwkynb29H8B7Uo01nFWImlifscDEyxuTh0RAee3O+
/hXKbvhslk739O8AXsGhU9qNCTR+lqj4HCnaST8kaHDomByNpoaUqcf6QEPr
27VIRQVmLdPSwau3D9n96yhX5myLXAdQNk2dmhuhl/C8o15SWaEOM5ycOwrM
HD5QiaAFDfrwBLdmAOhf6eTFjgzBLxF5aYcLA3SSPN56iZTNLWikYRwwrksW
LHQ2uvTKVBukGdd0EKfSsxm4KujFtsahq6Bh0oRV0LogsDYz2HnZOT/kUkUo
JNcZevgrNE+4LOmpfuEAhmuahKrCdQWK4e929tpEU2bvkVqydcu0TOPwPahV
HvJS9rsetElQo6U7cyruztm9CJNrqNjyvADMKfgk3PRtLcBaA1PZpOfM3wNM
RsfJn86D+eHoH+koj50KTF8sN66EMOm7Qzf5AD2uBA==

`pragma protect end_protected
