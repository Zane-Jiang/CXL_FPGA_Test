// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
dGRPMPCrFAK2qu3KnxYIuvYEC/7ewmgJxFPnCE8OHknfIcpdU/bzdaYaumg2y6LT
nry4x4jra+VV7LBjOJhPW6ZF15zkDqB65bWaLLnaEtgmEXiV6HV+PfBg7TSOJfW+
ohDy/uL2cYc8n2FEmwC6q3Nps6aSszgW6kN7P+mCYhg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5936 )
`pragma protect data_block
vsP9nNxzq7XsCxoJieXdKKM3CcEZFRXau4urpOoK4qYbf/og+C8nvT4WhLkrsE2S
pbei1wZubEwFHC7hR0PBlXcNm8YdToi4/1YIRGeKDTah4Iai98TFr3am5LhZ+/jg
VHTRU/WBa/94FsZgEXVCfn2EvoyTcLGo80ucUq1e3/oKUdb7QAslZjjN/ZHhajPV
50e9hL2gE6mWn0GDRGzt5stekmvafDFlGdmrF8obhIv8Fb5dV4NeAYzxlgYXXyv2
1Oa6gDT6hgKReGQ2f0TyysH96/Sl7E9luOPEPEtpCdxJIts1RNVzKkhPpKFAo2sF
u9LE1Z4lAKZhCrSrUk9weUepqDWlTU3vVatBNyOTCg4lqdp7uehC72Qz5kx46q3r
VmIG8UEQzaHlT1uGxlDa8sUj4k88rikcfcquoc1Esdp72gCtC0Ad/f3y6Q74FbM7
pXgfrwJKoNA5Ae2s037OIm2nMVIk0rQM+kcmCiJC0Q2ZYEyniQ5bKZAgUVMjAm8r
OwPnDTLsUaR7FPkB1166a93geN+3FSw75f7Fompa/rN//R7VC0f155daQRirUr3Q
i7oTJGr/fq0GSCgAkd/YRh6EzojBE6bIWHS34cR2gDhvuMiMFbDCH7ihdYsUJrpb
6g/PaAozuOjDupNQW9vClwOfMegUyiQtiqeMffaN7ke8fqj5piKHZniiOanScMmJ
KA1UfvDe5/xKcY8nLMoDNwr3tUV82IEB255Bklv9H564ws9mH05XASBU7KLTyfKB
0Bnkz53UGICOYSJxYoc6OhfIB5eHlqjOENz3S7+wAuWwQyNTm6di0FW312t0B3ZE
PuUcYLxrpdw2jjFEV1X+EOrT7c/zu/UOJOrQ7zK44KTuY1/Ymdrotk1IEdr8LIsU
wjRc9D/cjTUj4s2jijzj5U9pjBXedKxkaiSKWQn1vxoPVLBeqNlwpq6djpkywkQl
r0iOHIWWvFQNxOZRIuurSEFXY8WVm+2IjJGDmHercY2z1sNssKJpHmTwNI9C2ieO
6+zoaiV7l+uYntwFE3YoRtH/hah5b17Rd2uB6LJ0qUhuuEEvbB4HrDHCOq9f8Uqr
S21vfNXrMwIPM+ame7h+yIVYARsFBqFdVrLiNI28owF50pOhVaGVd4mOs7HmLF/I
G8g/CAbGZMgoEz7QsAuJUHyqDzI+bNeIZwhX+yoahSR289D3ZXRD6v/RnMQ+WW9V
UBWMO2uaV0WE0N2N1MUPh5h55NLnA6YZwl5rbuAS8Yl/IESbSm5UbT40HSKg98oF
woo88qjCPwtH+UL8inAlLCjxXXdXmTJnkuH24i/4IC8wHGYE+Ej71WYiN9qqh0mJ
8F8Liro6lhn18GAXa01X8mkkDtv/cEsiGG1Nizf5OBscW4+ipYuy2XLhD8AzBBlI
Gq9pYwlKZLKnE8wxadqVqJTuHJSmarUUIWTe1bfJyDJeA+AlBmpS/kNBV6bjtTgC
mJos4jRyKe66QFeKd5l/3xfOIpnuO9gO0WP4KFEiTQAjriOFkEvAAuMdmWtinaf1
J3V31zbQUP3XjLjc1WnogJoDfP62uKgzzJc2I/X/72cV1Cd+HG4RNeDq6pF91sFO
aYdusYSwvVHrEjMsvsfL6ZP2tj3NIBe9VQo/tAQfV9OmR+zQVoWtZk209zTVu5qE
TkRb1TcpNazbDzfB1BCfgmRXJX0vdZBGyyc6pD/4rtY354StTlYKdexOqSYhfsj0
+iZKodHs3IKFhAVx/Xy+TezhZiO4KjZ4O6W4ynH/TgpVlLHC4rP0YoXJRZrctsq5
YwnoYc8muCuAUfhAJdHgYqYCq1W+nvb+6xoN0p5NXIItJ2hVWDpHKlHTSpv1bbzu
KB9dliIA0CLpboCIS1/22MkhsDkC9ZQZ9kpXxHqk19ToNJdnzqJKep5Ok5OaEJ87
J5wScXcg3dmu29YYOK+lhK0qKmxE/X1kIITQUCeDoDqq7VBD5AGVslVAvuLrqxu1
iC0bvvTszd1hgKVeQCkUvO39EfDiDmb5xH1m73c5YGJXQJ0wIHuhwuVUtqN/1rWq
1kelkZlKcBWoMnMLZWbUm5Q3yIY31UKUkUHmilS51kXxDEI1LscB8GCE9UzHaDkm
U0onOjS7iDEdaAAzaYj+wOaAfLF7wCquxQHVK6xN3CDPq7X20eZx26zefOK4csZS
VnOwVfXOI9KvD9+oAAAKycPeX90nwe60MkiyMJy9/YtuVLd7frOzm0grxS5luAkf
jo78c0Qnsf01HhXeyf4xJa4NBqrukGnownhbIXgWYfPygTlY0GJ2IAcW+4TMh/0C
HduxQm2x6Hbso8skFX4BYC+vIg/oG6WvE9g1/JY5ImS2VgohwDSsBCP81k9PSFmS
YSyDDeS3+A+Kh54W2jv8w+kPcgnJE/cIIYBBKgAGYVuGb8zG5GNLrerUXOF6O8Ui
tdk0hi9IIXoOEjGKKFc0Cy4FQUDubVDuLxQzibvuGbf9GJQc4ydzPlDXg9rd6w4u
ERX88BPKnf2YGTKndR/Pj5yDm7x1kSmdmVRcSf+/Aki7nNR3Bn6pFAryFXlov9/e
ZKZyLgG17wkr0ts5HmuBfPbA/gqO2M3sHqgAUtaTQxQJzEykJhR7/Thq2SgsUK3n
S7/REGfqOxaQ+rkEG2J1f3l/DdZOpkp8cBzz+DNiTf7xEbTUiRrWPtbxDY6noBD5
Fja/934Mi8mU6j92DBaS9qJCMwEAsh+VW679ElzUXqhGtmThnZT7Ad/St3rdbVEK
+Pn5Ta6oTtf+jKTLTGQHEDzEjZ/SC5h/XwWnpUKIfB53144P/LrgZqSUavpW2OTO
O7F9VCogKkL8prUJyOgYNiOICxqIRNMIRJf3CQnuiyZgnP0P+9VL/Ifsknd2pOgp
o4LbQ3xxAuKSN8MEDOllTB9SQIEb/DdPOYxTy0q+P91R69FIn0Tk8kwaZScy3WWI
DC6uH1ctJCXSxtQXRtFuRla00G3OOZk2asByPDQhDNrt+ECUzvlwok/4le5KZ7/6
tj5JVuE9C95T3z+wlDZNJBK/GG0+pkZBNk4Sq82bmgVpqTdZQw6FMzNDOHfV9VNv
F+cLEH1DbPnFuCUjEPmtT8adznXo00197d+vjC/XxdSkZO84zYNfGuXMhMskjDJd
hksoAnrx/KEVeP/imN06stdsUgpibwWk5so6qByqCgPXWNi1256a4cKBge6lODff
zrxMlTehB6WuK3WVcPC1zQ6JT5ueA0Q1WMxlXLl4xkSYreMEfCW+XiYIErY0Cktl
PesX62nTspzaEmpsZHAXvgNFeIccI5/R1i4jMDpdPjd4++DF8tGuoMJhOM/0zMzo
KF+Q7PT9Qj2X9lnvSxsRd+I1SRVxdqYIJ6wJ2bcuyLUZjChs/V7S8IDrr7YgbEly
54KzJO1yyRrKrDEbGrJfdYPVva8P2D/j8aDtgJcdONK6h44l3LF/1LzhEIOHVZgC
CMkz8VTdDDWpS3TUj8XVd59TO4s27HL0FB4r9wRWyfkZv8yaXuEo4u+flFAK4+me
L96HSTOLklvqP9tcNMnAA4rz6Hf7N4PeZ0tn0Zkl6uHWxhUtCQAM5LanwuskRIfS
5n8QzcyUZiHSMo8rWITrOhf4BR4U5CPx1+uKtH7lwl0+oq2EYJ1xL98XRP4LlQVh
cD27efuax7HXgG4/NaLqxa1wi5mpqE57fjtYCBqbb7UQEruOzJ2wZbe/OEc/PJCp
Ry1iyQIt/pZSf7M3xIlt/IYEYXA4oeQxH9ISq81/6Et7tNbjgfAqvOITm0P2cClQ
j2XEs+1rXNeW/d9s9JHLpvv8CxTBZqVoBX2Clppf23nWRKfwe0k3ThfhJ9SHDWXu
Z9ophdf6g8nkcki+Qlu0WjXLEvxeO0cti7R+vma1WVbrrJCvQC0QeyXVbDGnpOym
gzJexHNK1UjZ4kgxRk265bQ3w19LzP+KHHTPT8TA7QKncF7FFVwePWoHk0Gqo6rR
sFV6KO30QX0RON7Vh5wFizJMZ26FSiQrYCBFhiDwUvnpi/BfWkJ/aba/e2mYM76d
rY4dk5mUhkTfv3lt8LhwdC6TyhSjuXOtjRKqksoDOjxAzRHcL1Fpx4F2fDAjStEd
e92v3+0IIk0r7tOMSOAB1+Mlfs6s86bauR50KDM/YUc+MW+tSeSi/8RyiRJFkqdV
sVdxocWoYP/5ZQrGSYdxH4aAv+nrOktbYc8hIkUBzm0pcbj3tN3EbtP1bCmvH9Xz
Ft3Xdc3P9G/O24qlRb2exxnbS9WPEjsm1jLWTCvBqDZrCjbp/IF91iONFgmC28/U
Tid/pJzZCVhbm2XpTWsEAZoDnagBv2zrqcoZbJxQJCAeHbmwnDK4ohKITniELHqc
NIsK72DjUA3UQayBJCtqkLKmp7M2N5BMb5U8uqG+fLp+pXj9Jt05gN3HK7IMkbTU
TqMGTRX8/6uNnrsWwEHy7KX7qds4OdJQHHhc8eRM9xtRYaeCrLDUaMQpgCvARzuA
E7aPnnP25bcqm5HcZK2cY37YBxhdRpKm6U1iq+BH7D/SZOn0vkJdryYOhTbGC8P5
wQKwUzvY9cHvQ3wY4Tiv0FWksKMZXB2vrEIPz6RGkJD8WGSJJKT4HgvVVWks2svv
XgN6HIEnukxzOS/TqfIflHHanxOkdzJ4M8Jdw2lkdyXb15i6GFV5cxUQAuMkdIvd
kCcPlY8Nj0V8jcdOpKj8AzrczJh5xFpPUaxKl5+VVtaEgHzfVrDy0zB1CMxY/A1h
HpXJ7pN0hsQvxOC+e0PdjZSLhj4MSNTTCFca/NnLawHHuBCHWSbV/CWbvcvO+FvO
GG2WeeXnTna4VEFWh04+QF5e6zQ5gRAQvPULRl/j3Up8FEXzF5KFAeCdWvq6Dpr6
z55N7xkPfP0tcrP0FZNMH38YhXj/BPBL34Stpt3wTIjmLDHTqowx8rGHqDT9vvMk
EghWZ3lnPYncjbNA5vJ0qx0yLwXHiuCoCBpKGwPx3eBpdoOb/+g/gZF/X0//UqBE
pRRL7VrXCtY4dr5z22UtnQwDPX6gAHT4jReTWeC1S/tt/BcFCun2ml1ZdjR4qiwv
JD/15/0oRvtR2DdnPaL38s9CSVPWbZ76tjZzYp7lbwSKhgxthNS+QXTQWw66T4Z1
pzafNH0GUaFlMDWiNOTJO8JqxzNfeFI1powUx+5L/WKIe792bicCgmlgUzdMlWwa
jui6D1Jdm4vfcIInMDC9V7+ssJbxverrz3pRlXLd9fD+WVeJwRlKveSRv7IJ4thG
69qZToxhNstW7Rs6LcAYz2k3/acDd3j1mUsiBsZ38ruu5OOoAAncjk0egZzG9IGg
xTj/nXf/bIt83HifExRuvT+5GxaBezDGBRav3+bHrfn1vsVQzF2OMmaneVUKQ1v9
0z8x+8qdvBoDaY8rfAvAIo/eVeIpzlFJElDeVX4iY8H8LUvklUH0QIwO+x+iIX0r
KFLGfajtKwoO+pQ3zBCkAjyvqbxB3eOcgNCEHHt+6EkZ5m6aXq5HAqq7/d6ujqWT
S/1DxGlSPppBNX5DjEX2u/cex4aNIlMCwtob62tJApfooAmRndi/kUiEPFGPBFSk
reOfnkE5iNlWWHQQoSiPR76XLlf7/7Nwu/NZlz2kdg+x+N+Mx7X++PEbR2UPDjJZ
34Nf0rftFc4HvCz9K6Pwje0B/Erz+3vZU+/7QW+gkZEL1N093/lakjKlpWCWFMRd
974XVhqBLoxvgXRlWQc6c3E2GyU+5E4RhJoh38zEBuGFRKAMcUlkW8coRjxsJO3P
FTzQbzS/fkRaQp/Q7M3wV7qa79D/e02JufcRRBGO7IrsfAKQDV6h6E1qyvGsV/pd
HyjXG1N+cTc9WzGsxjsI4MW+uJoOHkSgRngPY4y6UF2XGo7mmv7fAhu044wHVOOd
nWoJMwCuHQ6NN5VAi3wfRykYFE1bdnlvI/2DBNs+9DBmBm5hkE8lEC3eFmH1GGie
dsbZ6jUouCHTgiqVCWNZTleBiwyoG3CDYWtZ0A96dZmvAWR9Fcy/Z0vWSMR5HByd
FMs9euhnaG8IPwUuJRRe4QT4oaB2k9iJsKPz6kYwHl2bu6tO72RxAttdkqJzuEz5
9r1Um9pyeqoM5cTAoeeai4sDEzkriYpWgj6ro6Bcie08/kZMmc+WnKdSaeShrKit
e1YYfsWYIygSDoaEKSO1f6iFHe++RbA2yCEt6sNCcsaezFgoKpAzQBhLk4e+xqPt
ptlRAKY+mmHW5O9BxccE+6t+D9icWH3zk2Onwv15DVr0jcdJGIEkHIDYS/dTW1tN
X0CuPE5drjWud4O1cN8PoSErctirk6sUIdb0mpRb0p4XuVB1TnCKbLkQ6gRAaOrk
aS1oGSDRvZ80hUytlKP9YfFncpbacnsWEfGCTla8nuN/kOYD1gJgAUGUfmpn+ioG
z309pLMnpAF+hXeNSAwji0yO2BHoUpY3Nqac5jPaANgPkbf9nanKRgilJdX66e46
y4JYSTlVaDtIPpZpDTwyKYU3VSVPdH5EOSAU2Q/g6RRodyZfzW4P1oiP+Pn6fTOr
YbY2VJNdoVKbz3pDNvnm8LVFDWU5UQRl+45yCwue5KSVz9MDwKSjwBBbjrbssSWz
Gdi1wDfIhb+tJPQXhqzcUDUuHyMfsMg0BrmFa9SU5UoLZ+K1YNaq7443+w80bP27
jw3mxF4DyDVMj9ggxjsnmY23Pn91Xczvz8ZjkOrrCDugTPkk0RUUN7J62Pnqw8qH
gVZf35Yvgygwo81ZHfavVUX+5VFm9qbWtqcKUNXC2qfD/BBpnPBcKqQUroEiSROc
3PieZFddzzgewgl0rwsb6FObk2ZJ9zT53wOTpHmEiYAwzJxDYHb71yFF+Xcdk5uY
004sQmXtQCaZPEjErKpsqIf6KaOpRwpXSf/Ntow/sqIPar+DztgkwIroz59PmMZL
GO57evI3J5A9YjKgz2ZccKLf6A4jK0BEZNDzp29BDPHJCiGwTepwhwchHqCIcI2C
xV3SkK33miXX0bWlGcdr2XPtWg1cki+lni5isSQpm1/pqMfM9WDFlAW8oNwzySbc
RSfBQTdfY9/XVCZU+OLOQ/7eR6oHr0Wm7LCUPG8i915CIDlaL5poCTRB76VCeb7D
0tDzL0YeWn5t6bzg+FM+ncyiEsw0jsjIMPyxeKBKUvPk8J5I5KpbeooIgAW8cvLZ
g6vgvd+4QbvFjBf9WzepuDOM5eOIP0AL0E5QhXcH2GpD/UNqnKkN9VOm05NyDFn6
W2BAvArJd/i6JItFji27Km0M7g/8C28ypXOm52aU4+MkqlrVMwNPAJNv/HWlbi6X
Lw7UXYxCYutB92yMhLXAYdBeIEzO54keELMqTK7RRubk2tAHcyqYwJOmowbz53wR
COMHjY93wz4GjsDGyLVp7RMri1S+ab5hRsAqYJzsU67U0+pZzDOWG1An0+n/BKoP
Rp2z3aVvTE/yNFnGQLNxZ+ad9lnDNK90JCupTPleN9cj8oinAK9NO31JCKmhviuH
5j7WNTPl3wZCr7Q3JooSo3Bnxw2K3g+epA30Y1NkC88i299FUf9O7VlutlohFwbC
Ko9D46duQctAwz1pR6aMFNjnsg7AONNXt1T0ur5G7cRMOcMzDiPwSkb9R4j4cXjc
USL3iOUM48bKCbPSBoSlJK5fxv+IisuN7GvR/wkWSMKL5uUxEU3/p+eAQ3AdW7g9
0dzwEZxezln8b8lxXj75vB8wN6AfHGmzQs8C3QXH0/+NDhLDtXWynMkaASIL46hF
MIpERtoD9zcX1jB2P+wH3u9NknhP+SXb2HThpJO/qloWjcpkByI+X/yRUrTqd/7D
YGyY2aJfy7PZtScR6h/UqphhjWTp4v+yPlzEghRnzEOBW8T4OXsfSRyq5ScxK0rD
Yhg5pSpJtqO5znJ0Xt2CHM/KaenGcphdYGOjZAsNO+o=

`pragma protect end_protected
