// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JbSDl/Ycx35ZP1GUNJyW4o55OtVKXNxnS+tzdtO9JlD9L/ZSqRs0HXamUPYv
RA+LLK+raBRCWzMOYrFs0cK9fXKLWvfZZwpoUD1q8d0wPRsqrYpIgChpWOgo
zjPfvJoT0D+4WorijwT0t6CO5adzxDv/jABnwNI7uVu4NNxi0t1b1JSj1EDt
QscIyCFab9Vf5eXydRsJ3rte3EaBY/eGNrKNeG1FZqaQOB/pYFzQKWFUqdcn
H7w74YjYj7y/fxplJTczaJXTG5EG+Iv7huGWSvDR0VrdJ49S3ACBGe+fTW/S
+ggYnTlcU1/yvfXtdPoKE/4HNVxc9ynkImM7hOL8Iw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pE0Oo6JyqZSxjwjClWsgkO23tpy0QasieZmveHqUHDfBsysD9Qx+bsFLxAuJ
+svpm5aLe7ivUndyKK5C8kNs9hDPvFN12vvleUl7xbWM8cF2ewa/CaR58nEr
Zji7Hwj113anX4r0h8WqcMkfy+4dZ71C9o/RPKPHaRJ/eQxRIgKlyzJF45WH
jWRIN7kAPUo0rFKAoqA0EuuD6vcWeEJ30OnaJprzmhYHtKsKz/P/Mupri1JT
Ytnlt3bEpep245/ZT9tu39YAmJHQArf2PURwsVTXiQMH5FXklQft8LvCCkJY
GFYfCSKvKTsZbV0tyA/JTUBB42QljOZapRnGBwmxsg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ehaKUQJlCpFwcAlUjGIq4IRuq06PVLKBb4crQj8vFtrU5WaTXGjgAd6G9YYi
zTfi+6f04C7lKJQXY+X71HTbzoyCQ0PUvWyV7TJRrK9WoFYbQj9kM3uoU9lC
Vh7WQb5RfMAa9UNTKG30ZkSkvypveGSxigRnUBn3WpwSIPcULN0n+t1y9Mql
2InWkkix7JMeog0tNohKGSsH4c3ku0BEctz6eznumFwlS39pvBdJXKJ7hV6P
jdkp1CB3qU0d2j1mtNVlppUZOFnLETugfYe0Je8KHBENLXuH3QJpHMuSw8qr
Z3egfUD35+aliVGZrbKffBkCdYwjsblLL1sbFcMfWQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HR+c6vfORh3XTYJLjA+CyrQyTTx7yLArKh27wdMXfCYRlIQesJWazMaWOdNS
oiTmIISvYLxr8R9KSKezqDxoTF9T6PmGbH5Romdl8ZuXOjl7AeAIu5xZEpbT
FFc1ENi2rPyl6gCZl4uBy3itivI/4OTWGvJRTIdVnEDe9OHY5dM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rcon5xeOZ4Oejx7L7ivH/T9zwN52d0dCMKPZH6HN2+yy3wV6MmILZyYOkT2/
R9Tosci131uIEIvrCNLeO1aT1pKrfJCPb6db9auQoBHCA8fu9rs5tbDeFodJ
jpcIBSMzawM9tkkl97SLTEtDfGy9bw0S4poVUdv05ETfyO4rrWGvmy0GtJ+U
dVyevqeBGk8xVBgwBJNLfmPslMMuaXngngS1+TYnBR0Csric/Non9ioAsDI2
tyDX/5g23YAcyEsij1MlWAM4ErIp51EAMJ164SSR0UKf/zJF/KpTAiAIMuMd
SusFVgu3X8VwGy9LgNfPcHgVi+sDXBDwzzqxV1KOlElUvni5xmsJelC29tum
l/aIl30MpcxEPRHhk9z0jFbkWdxYO9/UITh5zUfoFXGtdg62b9879+/Ij0Yp
SPlizFWo8iTEjPSuMzMovWHfZnGtm4/3yO4Vy+iuMje5EDwpYPmfdR6RfZTA
B/tuTPyvaucNTO721azyTJ9C0q3W8+Ta


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cgRraRxn41MF718Il+VbChtW95Ur/Q61vKUyZs7LUUvYMYWQ1FthiBkgv5HN
PzffncXlTzizBUN3EAXjDtO19G4hddc+G8vFuANFtYBcz4OufBbu6wVpE68Z
HKThoSi8KeRS2onH4K8OkzdafhEKQN3nfm/7jVq258D7R8UcjvI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ayQB1gFa0qhgpPhNFUMUbN4W7dii8R7x3+6bT25aTv4A/ODxq/luT5fi+zcG
hJ1ebCEpfe2vTYQOhlCdDQOljkG3QC+xVY6/H70Mgat5vaLWcyIEh8i6nbDD
tmG5zCtNvfdPKFt92cJojKIO7UpSUIJZ0njWfaT3GyE3GIfiooU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3536)
`pragma protect data_block
JvHBsvD8uEjJAeV5IBzncDDP52wq/OS0NHWWp8YW/pdwgyp+ILPfO4UdOWro
rmkEBRxjTe+6dl5B1BMQ+hUoT7nBsTr7bn2hEY9Kjf9TavMu14NDE4iGf3FL
v/46r3ZPdCfEfTmGiQNLxVkrnzaXOUEob70ynEAzPNjP8tcN7tS26lIsAcKv
WKb3Ef+mOkN0LqYiWgPglph24ng3GJ7RJy4JR35WYeHE85ZuX/nCKE2Z+IRG
BM59GoxBTAe6pqD3sIxEahvBzLBWCe9PDY8lScI8AGK9W5JJkjim2Mk24Wwq
e3GRC3GVT3nirLt4FxKqdBlK8sqoHaw9UBVy5FKEKchKhoRhjcSegqDS+NDk
lOl3vMbPGj/hOHXD2wvia4YyKf5eGNYs32xTkqiOfJxqNRMDwCorTn27ZsxI
KGSQz/8Eb+eGsvhzH8yxI0lzlkeIrz8yX5EiBMd+9aCCmAomhPtgGSzbXeL2
sSp/iGOhphXSvE8xYYhA9QdRc47d+1Ws7h7fJtUsy2d1fMoA9yVeUGrUgY9Y
jNc6iV5/rQk2lZQYyzj1Dt3Y9lMZY9nCkR3dx2LlOJsMcU8NI7jfK6axMqSZ
24nJd118pIcVDVKDoDQLKdsW4wgZsnAe66do+g6ZK1V+/xlMmKMbtiKFuOrt
44KsU8Snx+oP0+T8UWCmBH9kO8vR6TMLLihbOCTr0zKy8EwdIlHpdlXzj4aG
bbO3KjMLzTThEJR92jMHoIaSUkLHfcTqSwRUkYTGAe5QeT4WKtqsIKbu9BnF
23mGlRghD0BEWsZyeGOhpixg8pFoK9+tgUQsnPP/TYOTFZZ1V1PgmbpVNdm6
Y6vW1XDavUPDumGWd8VRZnvU6kiuGOvfhjukfsTA2EKRPuBzxJBCC1oUGa9o
B0OeGg679peL4lrdsojBaIbMuxg5vO2bKbrtHNXeJp5/eQWWY53wpbex4g86
+xzMB8reHeoGu2nHHn3y+O1qZ5heJSU1huone3jT4Ltp245oVmkJpKmte4NQ
gq5eCNPXACk+JH7pC8ekhCflFx+bYXlHiTBIyUfZv/tmqHHwzK8t6JWZuXBO
Zkzdd/m6Ezj0x1eZwr0hAETfyIQ2GNhLwD7KfOWmIxggZhx/YbBquXKCgVAY
I/hvGq0BWhymOCqeic/SLcExsOj+HIZAZmKcpZguj7tTm4wgo0ZKJy6//r2Q
cU1d1S74bg63O0gCy3veoLQ7rTdAn/vLdUJYfgVbqzWUrxcSMz+jvG5HH/K6
RnlR6xrhewwg0H8pEiPdTgYt0STOSO+R0e0j8Cn4o/T+b/n0uEjmfhltSvNO
KQbXPh1eOdCTPxeYJNEaK7O7NasH/YWu86xWzo3kDoBaeTPK1GRi2s+8cE7x
rlbcUSTwOc7+XgjXSFLMgAgMw1ttKijyw1QuRmoIhgP6X7VSTt29yCejOYe2
5KCsQU8aM2TOhQWsEjnRO1FgskNDRcp5AG+JyFt9ftwniYLN2NMNf+bGSv48
rUsbvWcOjSfGeN8v+YfVpZWlw0UNeV9jNM/Ap6uhg1Pe/BmfCJ0pREhWIv3a
jHT1ahiWP8pG5br3XIIVik6RY+XT67s+XROUNrSj3jE3ZZqS1nJWG3L9vJb7
4xlrNSNZYihxu9NK3dTDwF3c7wdJgi9UP+EuMQXD5j1Rsd08XiLrC7EuWHeF
qMbafuKDhZp6asqma4LtjQcbqrM7VcVJ7vD7ejOsscT1hdL0OFJMojT7gSEg
sBpdGnS9SdKUBOZZ9jjjD7r8Q5QaZWGW6MUuGLN4OVzduzsM2qqb8HGVJX2S
i52Et+gFN8ukT6tb28YsQ9mjXOzzuWwSdUrrJsLz/GJyVc2gy39WL/IHtOOD
UZsXsCWUzNUxvXsKJilcNxFuPwpQbrugWmbcy2M99V5BJca+eTwU26Ma4qx5
xifIeHrEqMfic3vrY6XI/HMu8bEN8OZzhh+YJTXqDkrHcmQNJ5yJ/kWorhjK
2sdLEIYFq4p5XukwteX1Bg7wdEeYBicuvLpN5uo9wVHDdJjPw3dJsK8zV/fW
W2PIihDCj0fDFNcOHJQK0f8HhGbGHEjh1kd00Q4kh+eZ5nOswZTVhLmM4r8n
n5r6W5+pe1WCh22wUsbe6/GyHUGi9YdMGOLRR76bdgbeMAAvQA0UvKnNqx71
l337ICOGAvv9D/fzU8xj9o3CF0yFd5YghgHuHjSXe3TcK0Uiy25msaeqePcI
rrD21WI3SJUyHBzKz3xXgLdny3ECCZZ3lnvyIPbRq0OoJvR9f8UF3LJBcnpd
dX0bQds26IFGbFJwMmm9QZ9xgOWJMQgYr8yvB8/NZnTI2+2GqsLPvKTtsPAL
8emh8gR3QIInliWIQFYBhVEe2WPJoBdMExzfYbsPoFTIGh6xIvKiHZ80VDtW
Ez5u4RM4aGApNIHwo+tSpyj9Pl0qaPfof8HZcpVF81PZTnte/XIEqfcWKvHE
Fpe8D3RcMiFo3IwZl4UmXfa1gOrHx2J5Tionk/LP+kUwKsMKBTH9GzI8nKbr
IKVo4mwUotJZWGgxI5R9h75pZWY+MIsUM3EqN7WUR6NS9fQGJOWJI+MA2ar/
aqP+u2/zfn41vvoDlTLRxG6s99JldRTUr+i62jfaU1NJ1jUmTTd1JkCmkELt
bhKQ1M/GFMV4JKE10TMmHrCoGPxHrZbDA+amVfaJRbwytdwL2tIJLhPAeUn+
pa6KYNMCmAOB8p4e44gS7d4tDKbbySCMK8rn0pBbGeal4HHJWHnebMdbk2Pr
f0IitSWIrfvKA+4BQ8DgXZgEVXhfEV4dB4f+Ic5PT7JrJdi7iWM4LpHADE5o
CfZ8rYx8AW8XgKL8XRfAbKtdrkaZ9iAPRDI6by4lATVs5UtBC0Mb+66w0KPM
aB1VVpRrM16I4betV1YeJV2uogMUnoOkTNaHKQyVwEZ4mKdKkiL1pA8QQV89
D/u+go8C+z8uHLWLBxHTw5ThsKr917Hu3QGntvQ2vizqYThizsvNb6SI3E16
enbcXLTGs/J+mkqNg753egQ4/WHXQMSuxVolCY21rABU79z1GljAHyI7yQSa
IxJ70r/kXlSIRF/vdhX2fzjt2HR/TFdilVBStRt3fPR1oLZOEFm2nIi5eWqr
3sD7SlxDYut6y98vtkibygLanDDLs6LQOleIlD3nGVo2mqCkD9cAuqi85d5x
gW+BKIyDwEI5XRhjw2NopyWrLf5l43A9HyOlz4KrGVTN/7E2T9bMJfap9pNd
S38OlGpcd7CXVvUnTN1oE686Y24KbQOe/9jH7038D2SxlYKCdiprIHYxXZFC
ipsMUlAdkhI6Gm8uJ91k8YohyshGoyuM27eUHwKyBj/5S2uukSRPM1otOQ+A
g2vPces4Lvrt5JrhTrU+HQOdWIH12Qf5mbR1wpWOhdBYouTQZQQIgTUTIa6J
MGW2quK80wqFxHXMWLLM2Bm/aTtYRv5oMkCqfJI25WIEQMToxcSUhMbwyScT
svYvv+opAwcgvn/Nf1/SMqtuqF+QcTXNKi5LHDy0icuXXe1n1XxSfGgzerek
hzsxZlalVz2U0bfydY7HMbckLkWlQznsB1RkJ5wBOfwZf5GizzAM16bTz4a4
2LFoq075soJqtkzW3OEJZev4DU5kZpwIlA1ewZJ1t+5ECe2DSQ7DnzBnSJKn
WcCMectsdGocZwpOAXQ5dcr7lIVyyhTjGASXwfe16A10nkWRSWMjwhoBPfNf
R7ceUTntp9UB5yg8sxmpqu9A7xCCiXc4YWqBfXizQqVBDGKVU+8mYCPF1vrm
GGAMSdE4FD9rnCpLYyOd7fVUwcBLhDmBHWftN/Jg/SN9i2inC7Y7+ztZt9Hh
XgjYzKGP1B63FqKuZ52Lo2kFPDwQWkNKS5MTL2yDxkA/bysMm8aSYHLSgcW6
ztZERQJsncLXQbBGR0tlyaI6jPtzMA7UokMbS5T+xJK3TIYfvUKwGhEu5NvL
Nxe7RB1FQiIqPlvsCEAZLgLaUpOxcx8oqfgMfp9UmXZQGrNGHtUKXgD5plIf
5xE9zyRtk6UEqPdowGHpRTdkejHKTXfr/oEyS6QoL6B55zdcDz8BuEUEudvI
JsLkaF35/ooUe63asMueqdJlmZuyFd7qzLzNhkD/UF2Q7wJ1j7EdbVoH4AFi
hjlgFjCwmy+0uwM4zvORjy8Hbq2sv83gshzgcFy9Qn1bDrA7Sa8lvy+YTRxO
qLa+YQjJMa075C6L09up8DfGUSXig4EXPfBe0SmdIbKhi/5Hb3WcZxuy7ex/
sgZbHPNMFY9FZMW+jXJJGx7+2TVOa9Hvh/Q8a/s5n/OUb0mkRlk3dIFqUixg
2z+hH1HlFA0DLd7Nm38jrzTXovXBNxvl7MW8aqoltjgFCfoO+Qa1WHQJ8io0
dneOl3AGj2IhXkV40U5FCg2wqWCgMDCUbT5c3aOFWcbi/iG96tVqf7g6D/YJ
vaiZ8v6hsW3jeOt+kA9SlcBQ7DDffo12L9cPFYYDaiJoYw48Sw9cjMlnY7cd
wxhQ2C81dKmVtodLeQvR8s102Ix1C3HtEYe07mnLAln38ejchqwoqgnezt77
ZrmQLlknHu3d+r3M19+rvpcWNnyaUauhMYq8vYUGT9ynEaJjE8MxNykeK8Jl
kpjGfxPR8NVEOzIaoh3jP0eQv5PHurCu4Y7snt2ZJOvU6LRe26qZbON9As+n
xDVmowqa9R73qVDRrnLhpj7UimSKHpBz9NI=

`pragma protect end_protected
