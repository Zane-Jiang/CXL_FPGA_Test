// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
voEq1acrdVzDSPaLrXgNNkJCVXHGdKHDtLQdo53kpxRA06LyXgK5u0uvb+Sz
znzFM9gn5QMOBxYyEfQXa+CKpKs6Q2TCVzGHH0ZGjHbsUsRhTtBQy/v0K351
nh//tVbkNJrv2SCisoUg9QqmHZbeNaWeiRqskrZT3UgrW1Jg++GISw3HUECt
toSn3E3Kw+3Cb3vLx19lPGl3TncnvWb0/wXJW07A19lO+a0WFVGUJ/YM3KQa
CLvX2ZpECAYgTGrzDLZzDWD3VswLyNuPJM/6tcJ2v7G0l2SioSpgl27YMbVs
Pxka5zFgl5Dw+IW7vUnWDBQ2AFHnWcR4dQOaADoXEw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bMdsq7C5755jiRCreff0miutGHOjKQXIDal/ZkYKbJz2kr0MiVxLPxsIf25T
aeQtNKCPS0ZUeay7vqRaZm+9FuMwqNfQ7987voAzna8OQ7eMTL5HFFInJVWC
DoLGFxxxqM+wGUolznZpPuUtri6/9zalwLnWbw52RmbWrvkHjU7Qt+UtVVO8
vFTpQMijP1Dkj0mKdOpis+MsW/aUvwkxEX7LeqVX71/G6ic9MCeYkd5J2tfr
c7O3ctbwppV2BXnQc2yR+P2CBprZ+TmmtaKwuNPSpe4yhhI0HM/Ayv/eBkKT
kgqyk+9+Rmb7nkA4oFT6l09GUdQtAOD57ijO/za43A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hfJJ8gLMDsfB7EFJfONTCJvJRy6l9t6yFSgcVFW6kV8lsv8yqTds4ClUWwv5
B1Hmj3DlTwJv4B3hIg9HqEVLup3f1RHxyBpveZ9OmXp7L4n+Ma+ahmsGTtyR
ATKOY2Vczxz2gfOpDs3tMtsDiCfz5o2Gr/n6C8wBIZIALXna7XyO3lwbL7Xf
gOrQsGmU/D3bKM+viRXlaGhGjOT4ksPyFJIlUi40lkYiMwTe0I09a1KTBfD2
LWwSwYMQk+NQ4lSRJc85vDAbpAGEtp6U723cwFQ2nbpAJHMnbfBsyNT3pZf+
FECokicc8v60h/63IkIgZWKCT7WOIMewU+TC5JwcOA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GyV0Xn/Do/RwiT/xDHa0KTwcdzAsTYhG48aCQxGDw/CczLTLnNLfMX/ulxfn
ZOK3NL4oCZbWP6QH5E0d02ns8JaE9qwWqVNeTd8lm+tksyZOcf7qgqusuntl
i5rqcWXL+JeBsyZ+eFqsse+DyFpynyPPiRDd1dMy4N4I5igguws=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hv0k9iZI4bkqFuANgCUmi5cvncFs8elC8NQ5DooFh43MfgA5pkgf85a3U8Y+
pf+bsIYvHaU1b0hU/O0Uu/W55pnvDWGJWEcoewg/4yOe9yinE9GFWVEVG5Xe
owxSlXvhp+GLJRRHMqFdeEwQ7yWnG7rbYwDJkjCa8klS/hxdKX0PJ2P1VRfO
m9GmHqse1H614sNHDurt4OPYGvp7QqI04oRMemYJZGpYwszPW/yJwtc7d76R
CE3I23dAT8Bz4x5mlFyh1UKsSlWsAqrGtivvnr/0NLFK7+Rh7rQNZDkNeCQw
jeC3kwi9CickxPMENrM2algT+nRBbT9RpGAfvXaaTJxALMC7TFOFK3J8FMLN
tP/2ikMbcOhWfERDS1u5MDQVvdLda1plWqhcd+7u6QovUds96BLHtiGd3UY2
lGnlszow5vErPhqyqzrCs4pAoCHCKrJsxulr7SfA+K4/bVlkYHYpN/vk1S+T
5FTl0aolc50P4obRweUorNYu99XRJfQ0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IEio/3iGttQ1q6i1HaslP7+U2zkYGPgKXb8orY5We6dxDo8AEUYLEr8/Wv2M
OwQC6buRq8li96yPpDcFc6Kh6Qt86/m7MAYWdKRv3drXP0UqzOXLzdQ99KQy
UPfXi7PzaPPx6+74RdWagqpgloewBcE5vSeA3D3QdjiN/nvV0Wg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jNGvEapjpXEApqeIGUvFwttRJmv4GzU+PshTnhUgofs++9oAVZ1frUrlnvQr
KY1mEQPrZuavW9PwkSYbioLjwGhSq6KMHsP4XU/VBwfpmxIYAlCpJseKSwhj
X7sXLOLHqA4otRAcdXqQ5/QsyoNLCPkSqhtonZyBU2Cs7YpJ4ZI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10608)
`pragma protect data_block
AS5UVFdrDVq3clvbocOQaIwqyrbWHHu5Pryk18aSgkT1VRMQ6PbTUSyKHpEA
rU3zeYazK7H+4yRZYvhgNkvqlW3KID7ExZkCLJOZFkbc/ObBOeYz1jbhUlnb
AnhvH2sPImYb4iAJXTok1Bu8Hrc+m3h/Ah0yc1KlmFpEIZYjPhqKtTKmCtOD
gqrg64wC+Bzh2FHYnhupNGPtZIDvyyXIG6CkxWvPp784lOCCUOIPDALBAWsJ
YGikuER5iBcU2lNSztound8t1WMnPPYXzLNy1Na7embuhsG3FVpUXLN6c4/P
IaNl4uoVzTU+jSQKlKlDIU0CGaMkZQevCrPu8C91AJLUVqIEWkTsrUNomLAa
kefSbbe0J9hnFMsKhp71zFN1N3AhBdUazuJ+tqZRx/YtCUy0oqjRUrP5r/eA
4yewtMnrFZHlKbNOj0YrCNcnNpHIcegitjW7AP4L1VyKREjc+S0u/TlQ1NG4
ommFARC7/cglgnCrIcOJ1mfHThqZah7/g16OgrTrRBPRkVzOnZMDj/4jyja7
BdYLHRWdHZSaAiL2y7m5jyNNDKcvtdABEyaw4AvcAEzV9lhf4Uux9ul2N5wl
RszISSu5S882VlZFcmz0mHsAna/9brymys5fbuNfP3IZ0RwD2dNbUs7y9uwh
EHdlldB4i0Qr7V9IgLIMO/bmsSj725/bhsrzK4ImcdtGbiKCCKsSMnrXLC8M
1Th4y6ifaVxOIBgRZdFhsnaJHMxxDQJQIxemev68qpWBh6GvVcJP5aRV0QZ0
5EmGo8qEVGDB31FPMIXCgvAtHZjXJ6hxHe5Sq371lxoAV8iUGwQmNnICro1B
pjRQgjlxd2VENM02ElJC/u27nk+OvSVrp29cUdPHLWKKzBsqr3ieZiq5YZBP
sJoVcTyJOG8MRQ6AMZfyvrqiYNOK2xaGBhQulnr2mJ9N21fAV6tA72xw/yN7
b95j+jBvJPuaKjegiQTujH7CvLNUZbCD+oN//uTyjAQW3sccscjYRmonV2Jv
1XAy3rW95zHZl8tbN55hr8fwKi08MJyzyDz78q8DCePADsQ0a461LMRus11G
5LsMZGy4H4gEQcSyYejz+/uS3PQ+p8gcn6Zla0rD3QA/tjJiqJP48jm9tKr1
x2DemjHrusqSBcZbIAF3GVeIQ0v1Jv6tJf44kc34qhe4xR0K/i/dvnz3KKrx
SHKrR28FsZcL42U7oSWQwB1wsQ65MhR/MwzwbMvg/mp0wMdVJf+h8yGn+rNh
vQXo7uxLieGxulY3MuLFxavAUEPLVQhayn2FIYAMNnqiBnwzrydApMz8Jcs0
CB/page1DlWP2kE8z9NHcWkzOBCZfsIk8rBnhk2U4Ckbgnk9vTxh2AW7MhJW
Xx5tKsQ5eAw75ZuG+/Lw6DVIg08UveLEECYgbfTYJ0gZYbuACqUCJkAx5xsi
9M35ndtXX/PlCCF3sJPgcaIVwZXLlXoTy0HP0befJa/5v0HMuV9I5qWNlphM
bG183AYYQaP7RFV3b5HSHgrBB2SvjwmS6f+UckwOPN6y/whVwxtjvhX6DYxc
ujy3USqYFTR6BwaxMrYRggBcKdhJSoJ1AB4wdTZYuhOKpaEJK3C5abo3msLc
wYSUNjKVDVlGTYeHi/gC3aeuku1HW8OXZwbzJfToRBCgcQVkY7BmfWAKZ55u
iggbUhgfCp2k/HoKCcCVayvm1UCdkGmPEps1XBY5JBMcyMvwoq7PWPB8mXpa
+zLbBQv1QuSGRN3Ti8uu4sA16OgfgP4fjLIEuPCfKt/+k0Lbe5e5DzOMq4jb
94EbDEdZTVdSfj1N9FORmrAZ2MmYIzDm4fVOn6bhUOkZ2EgLEVpvi7RswtFw
w6WfMbCRKsHPYfmZt1B96V4Y9raePZX1xJoS9zINU63gji+FecM0maQCDQhz
L2tQFyWUNl/abV/vcAUFZrrutjyhNfpDdCrTKj0+gBU2mPhJMGlB5NnOpqbR
VyNo8mRDmJDoFQPTquAghobOocrZEt8ov8qBYxLF20fLSUYoj+4asF6WkwUy
Gc792oaVSkNEMSMKEzlTw3pJnVM16QqMCtiXrrgnATCtGomK1WfHdKpl6BC/
scz9G/V6tjS3J9ONWPWLpdHQBPuVn40cLfsQA6vtA2vq14UnsdygiK+YMRyw
oikIZASBhBvKMqScQNcaJLEUdXTwq+Jc0PZ5k193enfVpHqDktUwh6mvYpgk
megjoDdbFWGeoy4Ov2AnbS0Oyd4At4T26g8Q26VB9H0R9Pj6FuVsLVI2TVfq
AxBJGe0i3BrOxCYfoGrXA9TN9vGJ59Sqo3GeIs4g7yZRTEAlrZH6WBA7Z9Mm
D2na+Arx8HNb2UWymceRc0SH3ZSx/QquYf4jPYaWrH6S2KzBEyts4TGS0m4b
0B0U6R+XPQEGaod3gwTUvWz++BSxYp07ypW0HoOSNMSTeRoBG2f4LLf5yiFr
rCHS2UVbwOPThe1u7QUdBsukFcVg4WriHvj9yeEMsWXAOLGUIagB5DM7Z97x
I45nrov/BNJ56NwPN56tN73nqSDS9adtvWTE75eij0P6bkABVlz0Mt/vqGKW
e7otAzZeYRAKqPT/3EBJ25yMCS3EXTwGSDFHU1z/5lVZyJ1Y0W9eAWK1lur7
WcQLmLtQUveGX/po+TPF0jRdn/WWuN3BHpXlqqY9aW7xYMrbKOxDG+Gq3tw0
CCzKonlkdcQjvF9ltnYkI57J9ZfKB2zsmUWGauHlOvSj9/l/RY5yiRj02Phq
Z/jM7FQHNk1dk07cxV+i1Lw1PbexeNIetUqVFcg1+HkX5su0tV+OzvTHxCeH
5oc2NZ5tXgFaLdqG+ojGYsy0eDILpStxtgTBbPcf2k1UPLnbqa7w42zC0sQ5
UAcHHBgguTp07wDYsx57Ts0ZQsse0OT9Xg1OTsnI90Q7AVu5R9mEbVQwwf+G
vjFRz7fYN6QEN4KFGWGFIhfxcXp+wXm1is3FzhWqknM2k14dwf6UPvbzdyq3
20+1mGtKpiwqqs2z2mkEqCgsNA+An3qwqVYl6UYwg6c5av5bnNkAmysuFxSh
BC1tLdLHBWuHdpI8Xmdg2m67UViVOowndjXZgojVh+l6sNy6YkVGVLUEBUVm
zsU+Ih+Qh0B72Ut2/4SAfPBofw5cFhY/gSSA+U+mYgOIyS8njTItvKLf7Qux
nJWch8fKjWeehNn1xPI7pFpskAhnYDzxkMx+pt2EE0FNASWE0RQ6Ob/BbpdG
gtr7ZcJhAHJ2iTlK+bjD9QDC54ipOQXpFPXkGctlsvpbcA4bZIBkpEc6c7X4
30CVTk60QRzsathOK5YKrYJO2tPRQJbaJobBQuTIFOvwEMRlJllG0M9/cFbj
TC4cvd11RK9Whi9xWC50hOIl1iF3DqTKFJJG59izBR9Tci7iDcN0uNh6Zs3+
LdYKwkfvhAhvvqARvBKW2LdDgcFi+a6doPIWwgn77AeK1YxGxjZXiQ+lW4mb
zxL7hyKAk10QcJBc1hda6DqbX5PN8wa3/FDcViJdlP+B6ocG/L7uEsJ5lnQS
1QeOWaaijoBkWKITkbLjKpVo7M6JAHWQotcrC/nIpkx/e8r1hUkv3ZJSlEuJ
HkMdUP4eEqlaQBCL8UjB2ZMBf5ar6ZR006oRRhXa/UD+GuRf7zjadcddlPxt
WZUiYQu5K1v1a9legeA7Tq8Ru7NA8zrI8CbsSmFQSvXPnVLkgv7NGvgFGE4p
tR7jPgYI/ol5p9DgwB998k3cP2V/6OvVfmvYa40M6328B1tqHxEM6R8v2Sxr
kJo4JEJgCzAoDE4Y04iD4EdSaFp1vLKcerM66mhjVhQR+eqyxfQV1+k/Vk6A
trv9mjmsedhRCjfw0Qu0zmYJP1gSQiIPRk+nf44n1DZGm42jozecRHA0/1mX
N/VbtgEM4fqnRzsJMER2c+Ju8QKy0Mnx9PqXSB22EJHExQ7J+ywEB2d/X03p
5sNxOWuyjFCPoko5334/US2VAHkcrayFD0iBPVNgeixddD3nk0FnrixQ+AG5
X+iuR7S5rCZqX1ICZV6MZXO3qbosDa4OY+zfX8NOrd8sUEmIXkAvSDvBj6JG
2u0isI717h3n84nnZ2Gw0qxgNOYi70WX1+tHCQg1DDiHd1ZJ6paYyyZpOZMX
7Edi4xMJJ04yC1GPNSq+AmZOusSwMZIFxXgQhT22Cq3ueGojSzLmcq0DuG9D
2I9ICE43PmBEItXU9daLNzUbQEoEm8QjE9VoIFgFle7Ov6KC2nxoVsakJJwq
6RitLAvLyaIA0H/4gFgMCIvzJmuBimwnAjY+tBj3VCViBXhai1izK7zhvnsE
OCTKEH4xK7yNq20mm8B0j9D2q4ueg0YxaOCe8G7LP0qw1orAi5cHY3Ykfqoj
gtkXY07rW4sVIzgeLxgsoMcziaKc8nedVrF3ENDiH96T+OFZ62gVXfU4OeK8
HvUe6FNQxd6ePNOXNM7XScCuD2djCZPo2aOrWt6FQf4lIcSiykS9DkXqnFUj
i8x3JlZgSDeKeCQgZKB7C8U0FnVr4xZxx65cTcQs4WXhD6G1h9XRjDe7SyEm
yTINjX+WoGEG+PbACw9+ZWpjFQfKjLvprfcthS2HzsclzjJCoKG6/jsw24S5
Q+op0lTu4F5fm+Fer7nWOJFeqAQQ2DsItdE67cs1qMe1senR5BC13eU7sjH3
Ai8ptHZ52/ZUvubLz+8NUvTj5o1vhIjuh1kdWemXWDcHHiGYtTbeq9z+ADJW
nYh/sWvU89ZFWD9xWfK1aYMSCYhtVNYDAGu2rkAEIaP9rxicMoDLlUBTeGHi
MI+VxDhIQ9sEZ3afZvkhcC//3Ww2kI7cGrLGVAFmjYMlnQ494EI0t2ZmfFTc
gpAmg3LJb/66tIpOuN0foRuBh1WuhA76HHSugCpG9ADdD+S72oE7W67oqTTf
T4Md0podAX9jz0HVdkGcIqdKKy4+7jc4+cdaL+8w0LCL83jw0F7BhNLrQ7nc
7qRF3kRcCW45UZxxK008cOFdv2yEAjAyK5p0M8brasaValorNcEIzQJSOnEm
Od/pBu1ur6db+vqaJn/7oDDbkHaBc6eAmW+NgzEdTmqAxNqZDJbZ4H9zb6Z7
8MzypSn5B8xKe/hgTWeHlkrfHHGnHtWMDVzrNRawoxwHu0RTsXRSIVoyF4fP
z+posddeqV96bs1EWAu7XnHfubfI/iiV0GJWkI6R02t9IqfBtPi4h3nXdBM1
ouxcHy5/W5e89KQvP5+UaTLEf5nlShGnVdSkftxc7AGwnqcaP48L8+I53VYh
zx5AuW7MqmoNyk4xKAk2hnLLoxnKlUwNG834kenC3N2gZEsvGOrJpUmN+mo0
zJFLgs1AutJkc8goZlfLbCE31kqGNPcbNoa7Y1zB8aK95haJaje2xWyKpJ7K
7EgoXlGIZZHyBCvKDr8ygPpH0KQSWYVJ6lQdmp+pP0rFSzdOd5LwEGvSgvtQ
C7OG9T5ghEf0CMTQRKjSuF/4VWg9MKe6pdX3V7Aw8gsF3CDgjhsDD+pjrj6a
BEFQmz+IigreGOBOiOKwH61nu5L3//sH68x4AcfZSUMA8AiMbEhvxzRIjkAI
LypS4sXW59dyrxYI/bj4g9d0kOEUbrCado4M0pYfFFFHoyPFlL5U1/5P5Ne+
nSdyisKYxM1X5jBFTpn2kmz1X87MU/PmfPkP8K6z1vW+pDuH+K5UP/pjCc6L
LvOY54zSIncclVE6oLazMFHMt29WLRFc7yi/XeIengOBxXKx/3LkfgVVSboZ
4pbME+C47t0sN1c7NrWGGIX/gxRICcLIxKJFdJ/pqR965uU7iWjFyRKrHG8D
YBtmdC4SFCpZJkABHXP1vpv3VMq9gVYrt53IfARllfY5GKdM5rP1Bj7V3FIF
IDYxY9od2SbhQjennf6sCmCEc4eTJncWjDM4n+tRCdTl2ECv+Hof283t7xep
FQqxalf0h3ISa8MGmQtUZKQrdbKtCja/ZjRz50wDNsz7Z7F3QJyS/GYREpCF
ksqunThdZJWDjUo1+1B0TRYlnapdC/fpzUJ0g+g5N11D9CNaZc8gHfQJmAOx
PEfbNPfl6TcTOdNxRpoOcNozcE7d27yZ3DTomrPBRmOf5sO2zoV9hCFVJWy5
Z10OCT3596xvrFKo0LNqMt2ym0DYu44hOZyaoaGc5cFlhaL786vmR1Wl1hSt
cyPLHqPHI4YJg8GrGuU+sffm9LZfyZkB6IivPXJVnFkJ+MJCCH9XBdVURQaJ
f7YA4O6eLtPsDmzKkL1evwilC3NDO9fL4qtSlWJBn/jAamo+gxD4oLhk9EyX
qgKCUEZsh9qSgmZsCkUEYZBmqXEctE8WZYUoFgdCpyEGZjRnc819ZKxat//t
kKCDXXbat/k11yxL2jItT4FDwjdORKnVS2SS2S/EW/XhDeZ6716baxFipz3C
oNRf9bUf1cWUpyT9MRkKzBknv0TbaSZo6z6JiycENd2Qb5zoubUmAgKKCXtl
g84VB0WWF5NN1xqXXkztj+c6VisBLDkOVQHE1/KT+1a2Z2NoKB5ltky1cySm
0iGNggToCG5nmmtOW5v6Biw5yHpSiqwmOki+qp9RO4bIU4wckW09I4fVU4Je
yD8Ihzc9/ykz2RFV6AGmus4Ec/UQrJ6tNxrjJKgcTsROQylZi+tuZl0vkqKn
JqOKEYY0/jIRRGcRTBJoQI4LXDApNi7KzbhNXvrL86Nb5fYP4+AjrNpMMhsh
LzmMhDs9bU+XtIy6yVoMqMg/dNm6EfhUv3uN4T/7VNRjfYC0TaB/R3/AKiad
UxORNgXnqk3HMBv9C/Z4+NcdgSqTTsv4abWhbTkXVgraagv2V6hpbHz/eOPj
GN862ynrug+YswD4Ymb/ev5j/lftgbwhlM+Z/8mA+kqVr1tyUKx54ox1OmVL
T8dgRtSRooaTb2BCjOm24qxZ1iJgRe9ximb6ynFnVIfR3PRJZG9u/bQJJ3BY
Id5+JK/QyhI7qBSC2yctfnWu8agrNOS+YtfO53bd9+of7ujkPClKydZgUeSR
jTlfwPHSS14N+SjcDKa8LzikyHPuf9Q5OCas39aAqhNqPgjQrTO0ogFQYXTH
Ys6lPMdeNoyXopRYy+swTiuuRHugAlfSltPcUPZeIVZfGVtzetvb6TXUC3HR
vhkAUYsGLWNgsD0uINCLcFJzWpZJwbsgvj0JxSSA07sV2giviRseEpyxLjqi
0GPKyqV2/xRDFOxQNScxbRzvl7qM9pBPa1QsFaKJAKzLuMTMGXr6yFBnEVdM
DrRI0HKyIhOx5nbmaqWsxZKV0JqZcenHmsGKBz9X6OikU3jVyEq4kjz58FsG
FduYPUNR7tscKq5Y1Fkv6zth1kWBehZYKlPAx6BAsYgOuUV1ZUCvO8XUtu8D
vqqKe1UdCK5hjlFGQLDYBDStJuwvCfmBF8cFat7R+bxzotS/H/CHQ/Av169O
FLU7x1c1K4w6ZjEbWJJ3HrS2vqb0sJiZI7+F54fQ/VPshjI40f0xXq7dGgX3
oXzy7H1b2OMT9K3LNTcl/pETBQ46fOJHdCs8ptClfg0mtJiuCx3ms+H430b6
wD/007Zeh8vumncGn1O9T8Sxt9E+D37hoCz4XHJ28AeR4acGtcOkdOCJMXsf
yGQm/WLBJkx/cjkcN1bVirJ3H8HzpF59Yz7taK9fQoeU29/KHAWODoQ14fR9
1gl69LmLhI01vRrlzbxVtKMj3EYqTvhR6WNSVrKQh9a76HLjeemtzFK9m8aL
Q9D8ydexHemZZenQhPZ9r8edChLm6edR2FuQd4uFm4V8MIkLI5V6pmorY265
xDTU+dYLqWfzn4BJ1v8jM+HLyo/nZG5DRRwLAb5SI/dBFdu8z6Qhp+x+cTCH
7UH6NUJ+ROpfm5QRGBLVsoeWUUMVHzuL1s8aoe0W0hn7Vf1adDxHXAUc/PAF
bYU42ky3umM4kqPBJcOrYJ59jKL8JwMjwdkjAAShUifMLUo8WoYQoWVJtlI+
JZtoge6MVFEVPGPP0mv1AEAgLF0rRNxjKQSJb7Gl0UOfusL89OdxsLBsK0MS
uvHsd/8HMGPNHXNR3VdQcvr6l/JwDr8rkQfGKsMO8GLjDX5Nnj12kTJjJshs
Y5Yi3fcFGNFuXJM6WhGQFZNWFSlF+oonfd9ayGHDl4+1JSw1mk8UBokD7weN
eG/iibj5bPoa/kxyzxaFEmglVuL4rmHoobn7Pbh8XNjmumFuPdgjzyFPxp10
D32aDDP8128yZx/xIfxFJK6RhlSxLaS4v1R3XcrpW8Ju2JNEwa0J722vHyf1
SXhC3kmSCFWLxr1VrNhUDdo78rIOFzOBKhqoGLTzjh6WIlN1GdiO2nKx3Atz
Vo5qWY8Qce4Ii9X6T16pENYAt/2A5wb7fzpPVxars8VtwvnbloFGDACelPKY
5bRFhtVYoI/p0dDokxR84UgqyFw6fhg/lIZ28n/QFFMgdPnHgognd+GWNWdY
UCcFbFPLpcr8vw2r4ucShtYlvyTnHfisDaBF77nCW6ORIokPUHtV8vwtYWZg
AXlb4YOJiYomEjsJyVMyK1xmoIgCwMkrpBLEMYlXtjmLN4r0mKg3foksZ7ts
03wn5NmAUzwL2G/hYnFeTRzaVDoO8z+HeJkiR/98hvddVzdoSEJY7syCCQvS
j30fOTWP66edTCTIFUbk+ku/mMiXOzx6K78yiFMoV3wq/gGwj9Tf7MaqTWus
p0nrZlxBgS5pWpbRDzkFFnA9T1muvJs2n4wtb4ASc7ZfZgqItm54SzDLw535
h032KdBHmhZV8MmS65Vl7pFhRcNu5w2bxbe9Uzs9yhsD61VaIXo2V7Dx3oTB
qp3S31hntRonz4ZpkO80Iiw6DFsWSkSYSBeCbafDmwQ4lBO0TwR2LKyiZusy
02C/MZUZTATl63yhH7/KxGkLc+eMAr2Icl53gIOascY7V7O/6UB5U3IE+i7h
XWjBhhR+htaATnViHC5KuzJeN7CpPDr9xDJRkuInHutezP+Tpt+gixS+s/hU
JVh6EcghjO2o4WU0PJaqTZXuVfD0zvxSpvbG0/xnOzh7Y3pVAiQkX8/vZuSj
vYboyLuPCaA0cldOoeoFWnMJcuf2Wl1ABsMTCviqvraI7FojhgvANu9iv6uh
Md2i65DAJcRyFVJReqnnT+36/TUXtMsXqkAU7M7VF4V+Vq4M/QZGWEvRH6BQ
sNV6vkyl2l24zHNPbom6U4Y1pzpfwDCkcnMK/rM2ymQ8ARYifyEcpAB8BQBj
1Ea4RXG7/JKf5MhYcqp6RdtwKH0uB+SE2B5Ky2bp3LfK9tQXyA/2AeRVAbWY
kiKfY74xMTaCohhOOJd4lc4YTxcMYTPSauIEAnj7VgtoNV5FiwnxsRGZJlIp
oMW9airA5ZZGpfHnfgLnrDwXQifk8CCMBXzQfl27u3NqR6foQFO40CPqEIxc
qgfHw8+jO68MyPpkf7TKdeQ41M4b7GS0tixXAaLjuau3XCIej02cx0MGaUaO
tEdxF7TlpdojAP+G9PaCi4VAheigOQRI6fnN4LFKLnNdPacT/KsMiVr/bgOD
X2QsX44mOkKNDGTzOKIIKC90uG1xyJ+8moRFhYjYTDfAkN0tq7N2jiivrpre
xLQWegdL2HpnSWCH/RhylUFYRDD6gcydf45HRY31qvpWimz32uPEv+SCp4b1
UHwsScVDpq1/agpz1OINeNPb8sUAAB4vfMgJeaTddjbbO+MuXR4DoLXlomdP
A68RO+vyvtGzYlUJnW7yfTvIzwXPUFqOSdYqxygG9KcifI6lCWNpydcqq8ax
9wQcgTQCUwSAc+Y4DkdQUpW8dZD40YGjS+01sB3QwL85T5cFyEVdBipWWdZM
YNhaOSDhnNmjn3aG16e6FV5xZx+rMKEcvzWMz8kZQDwe7oLWOaxih0d2H81u
YcOg0tky1EW4lLonQOmeI7he7MfT/SJveIUAD/IXiytMTQDj3j90crPzwbYY
vRUJRZ2/BGOmcicUyvjbjlttraaJpMBxktAnHmK8HxxcZBp0mvC1t9SG87I1
6B7U6Mvdvu+k5MKxM+Ps9NcbTx4sie00K4tdKeLEMFM3YuD39NXaU4ohwERq
2zr+MXbcFv5sCNOrsV5giAMReFLYZM6D29QnJWdmnYm0nWsAcsqGFdLkXu+Z
y+A42D32rqg10obJ5DJ+Kev78BTBDivc2S/qEe4zEIoi0bxXFLAWIbRFKxwy
Ixz6uaXeBQ093FsTo2OlxiD2WMQxdHU40Qn7DBD6SrkuykYwp00WH9PDKQYL
AintWg3C2nNr4iYgTEAWVH4pcr7vLnzjR1H2evzbTlXyBtVF4xI796ep1I6n
k36zbvbUgKniP3xADTpI4QjNJOroiKNTaF4mmWufOV9NAg2dN0ZaB350Nduk
p14bVzzFuc4Bp4jugXVJ8sP2yKClG0AA5VMUpgpDCo7wAm7a3ZCUwazhdNp5
i0K6kXaAWQAyl517gNek+KuIm+sV78cFic3+gn1+z9TSwerdTc3E8cXu3pGa
dHKI/TnAgL4XifZQ7hQUSyzqEHjkYtgZleBPCEVz8Rwglrc8oeoTZk0X2MCW
MsMNXVfYSz3isg4NcQ4ZHPyXNOTsn7GRyXPz9cAqit7JAJkIEoghlgnA5rd7
HFIUcUoY36zj2pzrVxPiRNfQef8FD3tgBBnCgo4726O7xHOXGfyzX5T6Sna8
Zaz7aTdhMVNeO0h2HgScKwNe0WFNrDIRswFEipu/CSc+37enudn6aIaYNeQ9
XYB8R4TIqZadJDKbzMeL36cb+yrjufSfhjLMJgYPKFJ4C2cOTMSGJFzAeqhX
/jeYtVg12XeyZ1vWEV3wXlUQBdMww0wrRzMFUTs8EBHOjbEJXA6q8Mg0geCd
BP5caHMbP/KLBMUS+4UQ8PT6qz7lJJz4+lneGMba6Ir/bnW9Ttt4yFjpG5KQ
Z/dcUbDt/QpRiUFLtTP446w/mcI2xF6kdU11mX392h0Ta3TyxZjNm/AuA8nt
gCjUV+AwMoM8+YN3PnnxgXZKUcuS7okCQKsVrewNn9xetliXAu+/tiM91C78
CPt74oyxZOZQQpBYXKXdAqYSLnPFa4TZODsb0C9InFKpXN0wKtUpuUzLSQIH
o66uxGhtMOH9wg2tTgFnge3IO7MAP4B0++i5cil6X8mxPCm6fBRAe11YV8cO
ikcDH1zxSrHV6cv3HUvOsPm6lKtqprHhm952ypyKELnHngWhfYN0usF8cGh8
x6YuSTaWKz5fKV3SVIKOU0kT5sMkt+qkqP8i77SkvXsY8RRzJUyK6wxcyqf7
O779Jhzn7XVhUqZ+ggVApHvlzhzZ/CQOdl4HOZBRxfpTMhBFburqwAxTQ1Wu
8jkFmu6YzdJtsZMiM8evBE/hKpDE8K0LI3GFkbcS3L7or/ZCOTxXg/n0UNqc
CmE2F5DDtnqbgfCIZifj+SFipfFPr0nFcCT+XjbFDM2/gs88Mm3CSTDbe9J7
+npwF6wNjVQHRVuXOB8zWiyjewgknno70eyB+WkUcF/xab9iz4rTIXp5Le1X
bVHmlbtVlaPdrEdftORqFiTFfURyzN1x2iyN88rCnyG9pfWjrtqEuSmy/DMa
7BHogSuV4WXI6/qlr5LvCr20DRZzLY+Dudlt4F70PPgmCT5hCpbzeU+L4EE4
pnWzyUGRAj0/zIJVMqIUgsLMVmNkozIprhktAQNKoQnQVjrsOvkrLYB8m+Vc
Eiyg3oPcfsTQI5eo/yA6wxOjt7dNUmvELL7oveL2uUrfSG5bU4d7ZZ5z7nwf
rYI4Fmr+Fi26V6BEa5dxxLmmXo05/G0PCzgZ4uRF2deHj2jnXXEqFYgR0NCV
f95u7i47IhILdpO7vsq4xUhMlNVVz9iSbS2Fja0P32ZGNOA33kpTh6ECfWZw
+iXjemypIleKM1flCOfH0dlvkqvFJb1bbIKFb2TdNizeKZA5QKpGAvWAqh01
7nQX+nn0vA70Ggpp0ViUpT5znmGclk/hjbvKueQIyokQ+Rf/jrK22w/G9zl7
+kmqYrlz/WerIYnJ24zdJanmtVHTzRikbxl5mpERvqWHnQguMBX9ZxCeS5Br
TUFNF5wyQa6ZhacOcpDARhFbbytpl+RSmWW5y2F77LuhofSDSynaGNe7WIuo
X5tfxiAyrHaaoExRd5RqiekSL0pSj4BkBuzwK8+1qy6I8Wli0Jt0gKw66vKU
OW7pYSFbH7plY8Qte8waji4aW6N4xaNd/MQd1LiBBEUN23lEK4UXCURhiXJt
s/r4xUmKqy+V9FBgUM9oldt9X16Zbgk7ImBSrTnev165wlOgEbut6HSg4vTC
MVC8zFtmztTrT8mNW/ZsG2O8TkUKffLdSfA0Yp5WWhFcfrSni/HqTu2p2osg
RT6KjwZg4Ap7+6BVEU/m1r0SlIZQnm2lMx/H9m0xLgv01KWccGUcWXpQwmos
DZ6acJ5E/gR8nd8hDKCgZZWkLk0BgJHLSldQiFKOCIAgFmuARvKqKahFreHp
YLlt/xfgE2YqEnTMvG1QUDbj2dGDdUKSGMotaB5h6Cgf43BFcnwp7LviQV6s
0MAlLqSozieB0hZOxsVv09sYwAAMudRWCwWt3P66VFPw7mbJ4eC8gph4Ohbg
hUHvAUmPrtcTD/7ZUqbGngt4kKo7qEBICAEIJcwceq8zl4ZzlYXCv91kLwV+
Pc1zddc1UMPsByG302/90+QIYWAGaQBo83e9pHPzgj9VEXphU5c8C08YpoM7
dqpx0rEgnQaQedhvhbbOr+7fqIY83e9rmJrJQXEJEwOU13uA0qZPLVQAqD7s
Vv5mCAplgPt8KkYCmJt52VEYLeE9ziXnyH6c2OgpPWCsEW1TyUAqD2On/1i6
zVEvYeOK3vX68FcK+whtJWvJDG28ZNZQvxYfgmJJrifgbVjrMuSknsODDKht
vKPR48nxYK6bOGY2I2s9ONi55fPBo7WYf3s8rciC2kKhAxuD3x6yhjr5fGoh
E5feoGIh7ieA+S/+TQqI/SO6F3/IEU/XkGAI+qX1rqVnqtvGCsvw+5IaRH/e
vU2idKiU1+mKlkVRDFYKeWIagGRTiY8I07ulBuR3Q+etKOIpJwffEvl8D+VO
BAD4S7vJoroJwWVZWcT0mb4QbFtxZtTQYB+iLyCrEPajAp90NCSTd5lA4r1m
kmO+yJYezdRiSrscczOKirSzkDtFuHCiREmDJVIYWoz3vAcGOy2k02coaYQ2
oAqICgrctFEd8BHQiWfGJnQKklMw5EmwsZv96nWpNLyzlD4hufz5laDM2IGf
RcBfCqv80KoIsOewqB2c4sIGC45wSAzdoLtUjMP1N0uJiLXRsCaoGRk68rcM
ctC7u9wRETMAOs7p58CwSs9F/5qIyyFV/dz7gzqIkjmnPMkZ6vKDOd5KxCph
FAPWQt9YCWS9DKirXWSzBZW9umc5jE7OgrGMsNloq0TCZbPW0Ybr0hQAkGUJ
jCLdveJLFwvJCbgPJL++CZQwCXePP54v2AxYN6XUaSI7pNM5X5olxUxgYekC
bx/xVIb7DgEaaeG+K9kaZuQeBNhAsovdCpALSX0jPNLYWTi9y03c1kVrwZoP
HsqJ2M0rBN28LGG4X7yf3cRWPoRTRPOev331aV0R2M02kncrSXsTFkUMe9HT
bmQBLBcpnX4Rpxw0vaz5n22vuocjI/hYQsVN/1ZP+Aj93WTz5cKQ/vSUFhSf
XYXONen9V4AY7jUye+6z0PVqJd8QBrOXx5DarVPjJMrPDt7WLLAJg7VNZIBJ
Sf2uGwz8bgoai+VBjf2ejDhcG+HQYTXiXqB+ETf/4t/kJsokRGDkuik2d8uu
Phli4m8aLtmVnN2nQwlpfNlczMm06ntml+eq7mtK47dYSUrZFgYw+L3WxYx5
c9NNLl+TbbL/F6u4GyEMnIGwd4eFc4RcCf6B1THhdcR6hkSxuGgouRWX3mAc
KTez35G6iBb7imz8Z2AmPUN8EVh84NMiklZBXnCXFxPaKqdQaukPewFxCRt5
7SAgSdB2TnN7Z1YW3GfOINABxuH3N+Tl1ajYTgGNQV7X4Ay+GvkQpEHB/tQC
5g4cxCeeg0+Jme/rkdPpj9Qgf7as1GLAUIgV2t+7jQZoyrg2RkdkHrGZRSbq
yUrPJ/pwmNXPVOZORCrhUHxB/AazmITZe/aIBG4Yp9Jl

`pragma protect end_protected
