// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PRmnsEubW0mSOd3Yt88dAgpNkfdfFs8GXhoKQ+9kPR2zX07BiSLSylD2e1s0
WY4cywDzmFO++5OiBpqVHz0iP5pei6z3tsWa7DpWn24CNLwbeGN1pPZOTNMz
MolXHPUU20BmNU7IFhrl3xPDadSbdcKNrLSq9WRb3Y+kr8EMvhWvZrjT0jZh
lM9NUnSCwYpv+sySARafrsncmErSre3gHyNe0GwA5Y1tCzOz2gqElQoXWqVY
OUPzEp2/vqMSEsC7prVRzqf5ZYJkY3GV+uuoGu6OohUd1V0FOvBhkyJQW1Kd
0jv+mDQDME4V5RUjxJ/RpxLJWDMxD8dD6OV3c31EOg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O7i/Zn6DeRhX4W9YZ4KhdtjdGf0iKB/0N0YvE2QEYZSuGU0SWffSEx6npUFd
8TE7hA0Oxk66Q9KFwS2Sm37KJZjuizSsqMk3LfyQCYs2jq54qJuSuHCjDib3
KvCpHPGWIprytqKMjLBrVjblq/a/tqnW8WkVYSAkg7sby/+u0yBDRhR2hfIh
Gacis3SqthPvZs22zFdqesvmoaF7cPM0qKilS4TwcG8i8sk9n3YZlmcXAMAC
VpBriDdK35H+EuRYXj/NyqqUwZ5pZtApYBx+UYdvRvkzKbdgdg+ffKUE/tD0
foHMM0hRFhxVuoa6akXPDbANDLoEJLuSdUSLyXYY9Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Mu7aIroSG7uTBbxiwHamn0IOHNtZtQHzLkAtz386JxSlHM9xgHFL59QffcHO
+noAcpUXLUGm94/dA2b8MDkjtNagZSKeMaJlHqVbV7eW4Mhg1S/FIueIDsq+
XiqS6+8E/6AsRkhw/wgcU83czwe6JL3Liha1Sx53eNzxubZdwLsWs4rzXl4H
VCGbuE15UlpaumKaIvYAy/HQo8RxfUQT4dapnjtkePlM3GKuKMaEa04C+BDR
pPgNyHUoi2572qrepVzpYUvi1C9MWskDVwm5fPDFAu5YY5PRLo5mqgGwnE+I
Eg/MjIYjwlyWBUmeZ2AlvwoIPtyaB1it2xoV02d3WQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lmaoE9250d5Exco6fmQgCJ/FyCPGD67LVHRq6Ep1owlxXkE1rgbRnTBlKch/
DJ/3va5wpgsndhyU6YTf1/j3Oxdzcnar0XcCGtEs6lp2r1TzYZcfkOBi5tHi
TO3FtUhjDBc53ABBVM3LiFT8mZ5a7LOB4NwKTqiXshm09XR+kI4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LoftNPn0DOrhwUgZgGnTqHlSXgw1ux49Ff0u4U0uuan7CdpKpOxRHRbUr7Sh
yiRzuQJGJITPRDYLmCGbjLyO09uxQTCbYJP59W7Q0aaU7hn7QxTJfZKca3iT
cKyYcUWDZ3oWmEVXyl5/yQ+zihr9PqKCXjJ2hAcLcbFTQeVhJ91NnqbfW7TL
mldan6j7iuBy2Rb10r6MBm59xl10d/qRW2xkcb2tzjndEYdatfo7y0sukrQ5
q77qwFwv3GOdb4ItZLck16RYQwGtlYwA57xXsPVtIilKzZ53Wu4Nvv+ayU+m
EDap3gTTLYCv7wz0bfNvscELAUy3VfcXq0Hchy0YrxXtogI81faZacwhCvIk
0Q1oqLgeOOK8FjhE/RWWO4O5aMDZ1Z77qUOkRPw2XtE+yhrBcMAuQAWVpRFU
9dj4nKNWiaacG7qFXaW0Q3OVaVMl/Uf0PzSuft6x7GQXGFdxQPp/XXvvHBew
ruvGiuGMqbRDRoIIlD8pxkkXgwF/lEas


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XEtnK279QFZOlBfACqj0Hzea5pOjSQYRf6kxxxhOk50TzWwKns1fn9H+42ES
wseAMW/bJkTBGOCG3YhYHfaOsKZq65th7l9gzqHBMcinV0zDQJtWTv8F+cxq
HNJJDA/5aWhhWWN3YzkA4x9UMbDgHkzzeoDPoTQgLXcCtVNMt2A=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hrY8VUsVVRgJ+UyJS8JE9vSFeTT3TxYGHta+oAJHDPUD4hMcrAVxjPr6FKFX
cA3J5sO3wXK3UwuFteJC80Z+zI5rgFYQYUWghlyf//Ly6a21/t5knM2gW1Dg
Do2Qd0YnA3lps739eBtqPg3WwBu2Q2QJdBCXvoOyEJvplmaqqaI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1456)
`pragma protect data_block
Z517IJ9ZrenDlV5BJo3ZHLceze8KFutbpEUUEDmB7P/jLqSDX9mtM5NgL1Yh
ihUUcUV1+d2At/ZUpoo2A/BQgKiq4KGUdYjibYOnCLEilV5a1u80UL556YHc
MCFSr4ZGi8heF0nQdfHjMMycXNA3NE8MwyGTR6w5SJibtN4SGEmU5B5Idh8j
seM47HhD3qecZr9q7ZdlMMEvdXzst1kdL+72PULx6Hn7f5paDZ6o5h6mGC0s
u+/E77H/4wfERof7N+R70aX8g4B51pSfTiGT243l9dQTRpEa9cLigHUU0W73
wJ+j63P8YgSVVc7bBvv1rIHSp+wvDBe2QYu2b6vYTl6rcwioMm3lk2vUHLJi
bDEXjpo4z7eCDhuNMWegB7RWZjFxgkYVle1bpATT7T2ku5KXG3/YdA9Hcpih
dvfzK1xrG100+8fx1qD/Jg4eMsSO5FA+O7Q8FDI7hCuvvJFtmz6c6nsocxvD
7krWJB3mSV/tJbkwPB9MOC7goRdijTelu3YLDskTYr5G1k0R0xjTQ+scQ1R8
EIFIGHXfcfEu5yu0AgCF/WjWH9T039F93zdN2VEq8YuD0SbFWa5qH2cTLCVj
jo41MY3SJpgBmJNN6LSZcMRqrAUZneNLwfrKjYp/4ecpqbIkLaXp9gqCxDBl
auEoPHxLMS/1tHSj97VdvMi94MlCcjC/JuGe7mvNtEN5+9o7pJ7Whifr8mti
JxB7ULOa+HbifkMSds7VC3v7gNXGUP7CBwgGzMpk92Oc7wu7SGXBWF45jeSH
sjr+i77A5EE7O3mHK1O8jmROSTRAC0feQJqrnpNL78xsvtGO74pGUu6nwfqW
aaEdFlZy/5ub51JzxqjaYzu6oE+D8MrKIGmKPMXUDcEWLPIUryK3bChS11jQ
ui16KjMFJwb05lEniSv8uBbvvijIwq2ea+xywEbiVTMxDzKc51QN6Yyktj13
bnukHevoHQ4Fs7797E5VvZCWCBRd46UhojCBwsE+LEIocsAk6fw3TphPS880
hjuqYGGgThWgUwfyKsUJjezZKrWsIDsWuVjyvf9j9yZtNn+Mc7ha+er3NlNN
SFg6Lgb/kYaViGCi2nZ3PYDmDg/LCtJ2Xe1YrrhMab+qt1HU5JFSbjex0yuX
tPc5t5Wj0+/68fnPuV8wN188svTj6eMV7ezuUSFCraPrQanwLDjwvjZQ/lWa
VYZTBJm1cUONB+tcZ6P8itNGa5T2L7zJRQuCEulpohUOibJid6sxAj7+gD01
8xLWTi/48qrMCh1v80y9HS/QCuqTRxJubtGfF+aU4IHsV98P2CSMbUc16hq5
rmK8PKnTHOcS91STORO6ZkQOhpkujrWsF6oA3+pUGg+Od7ueqkEXsHrklfuy
7d9Yp93BhOF4Z87uPUls2sKmnUXpkzbQ8V/m18b+ysAhLKAXoucvR3qLen5T
Q2Qw924ccjwNMQDU6oT1rEr2hloh43gnbQqz4VOpY0NygJcsZXMdgdXSoIPV
Fa88VbnvN+dZ5o+NyV8PIlE2FLO4SLm0rczITrWraLRM6wq3NJ+Bd8QpBRf/
yJT2u+QjfRB/MZ1HcEHn0vwQoCHIlhDgcuFoeEvwR/3F2IwqM1g8bjmGDfFN
5WrOLRje/7UOSUV8VRqxvouSt3lY9E9ThqrHSMt13OA/+TwzgQ6TUOatNXgA
fVJLiGcwhpIUXxwkSci78N2Pbe3L9z1ryFc8gO382cGoSIlLmi29VycWGldG
UAuyVRolD4bHwQJg60IZCDvNNt9v1iU7v0oaZduNKVpkjoeUc4aNn3xd56Lw
jE+eeJQ974ghuH47LLDc2o7EoKd5qOtMkPYX/yfKibCO5Ldro5bE0tFAH3By
PuTtAwj/j4TCETQei9F4OzXCJCcSmbp3NVp6rWjx7tOCFOiAePm3bI2C3uLz
tqcx3LQicG0TOo+o6e+6hg==

`pragma protect end_protected
