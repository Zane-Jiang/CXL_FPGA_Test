// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1kqKYl34sDXCvDnIVMKs0ONizjUGNySWL0ZUBGieJc/Rh5VmfpL3MUXHJ9qizOdD
3Ii34Yspc2rmYfdDwq+3+Cn3yP7KNSL342gYxCzacTJ5e5EWOwpphcdPfRdzMaW/
cO6XC4b0HUyDXHq1T9LMcAofT7I+JzKz0pdkzm8BnCA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8416 )
`pragma protect data_block
LwN3jvKzv8Y1YljWBefP1KDHrdOGf3U4v5PVpwRYzk4TBzPmVuJz67or4rOs7s5w
cHn1b/s9VUbe8YuTpKREmV1vgMYNeIEn1uyKxqjDR9gbWnJAKOzZHnqhZk/aiTix
QLjkPTsKEY8H8W4q17QEfa1HdNbPafP6nuPLE4lJosadxBcppSX6St30kBAltMD8
D4/DiS29wyLkXJp+b5dX5zmUd0Hmv6R6x6zCAjByq/BORyc3TI34B7QWTH9V4HK7
m+6OHBjXvKGE8RCtijJaAItVvaK3V0F1gkXwne1Tf3gfS8lQRbH0HMN3q3SmsYzA
OOurzPuxSVsSY1UQii4KHHBj1z3J/DHz+y1G7COeM0XhqnQumf2b+yhF36hh0Wpu
cYL9X1X7D8kT/CWspt/nh0XsOF2E153cEFDgMIkKVWGwBQFl3hmryqSCixnVFyTf
TQ3EndmG8Ext2Jg8MFkrJZVrhFb8t27Mgc8huzSoxtKCptf4k01nNRlahyoSVuTy
V/k53wh2lmc+/GlKqOvn9bAzfLGv9j9lA8/7BGSv5XwZljAjDd92qQuRE0xwGFna
0bLdeIwP9G9yRPV3K5rzRZn4uiNAqTOA4uKpCtnFGQyKemg+7WhmyNt7rZdsHDGH
VKK3a+35dbKG22Ihv9MFnMKRQM7MPsXmCrjHhVhJf2AffFgzqT9Jxd7B0r/HHA0O
v/AOFroVixPBr9pKGwRQj0uP8zwxksl5LML1290zN4WpNCMnJbzzRw3IeLFsBBZ0
n2jhY0jMKCSlFdb5Rlo3IDJ5zebb960FFvePmvuvlwEioT+rvzDrE2o2K15nAAiz
gAtsm9NCiTt15qHNaY+VLJaSjYsBuSNeAjz71WGAopQLlOyDGjUl2MJ+pmbyTnqo
lTs6P4iZq+FuGjLtsdspO3lqA1kj1dVfsoULLWEXtt6tp/qjOHH4t+Oyd8MRhihN
LbDZX11nJlB7zttrUfhw1AIZdfGwQeS3t8uyD9yBX32YZUllF8lJAH/lHOsP4ZsI
zXegoK7I2H+d8FEObLzqabdA3AGk8Ai3Oe/TzTRNRMmJJeg5TqBdEpD2fu24kvUa
3Lt+nMrSBzZ/zh3RZ2aAxfRYbECCBCLXWq76kvS7ND09O0hITy9us/cMQi5DVLvj
kZapYAlr0rGAECvDEaIB4AoHpABKuBJdIsH+36hV3tvbdAMkIP8lQpJIft5tLrN1
F1XVy6u/Bpm9yYkMaYE49dbrUNslvsPM6ZHGIoNckoT1Uo98ONm0+cEREUokELl8
9rh12VpkAq5LUitsq1X90ABj/C8QIYqQHcd7lNMRyoht1i2R/eQwKseNOGjS0y9l
q9CTxLxp692dulTJXAU0EpF0T4h23a8CgWTZ65YJ9sh0ifwI6sMiGN5nNehi61N8
sOz9S+0iYbdFxGRVC3HjNavz1gjL136PLHyUfTYTtLHRDx84lHl6qagRZVcqFu8h
QDMgtzs7juiPzGZDf7Mfmagp5xSfP0pDDtTZMY+VsWJXtTp9miw+Xk5ePP/8nmN4
IwEJ5orLS59RggbqxGb6PUpjRWuBiWDL+bMBcbNw1dCqRQ0L+sqLyEAmlGCdX4Wr
Ml9XoyJ0NHluidfHpkDIglcGXchoLiVvkmoti9E0d0WwktyXY81DCEqzEqX5DAXY
gutY6qUlSC45EV6HiNnu1QsW7DppMsesZ0pC7B+acSPXGAsC605c/eFkbBQosu5A
yEUHYlFGioYq3JLPA9eYh68o3VKtVK+WPbsMbR1PmFPn75NCrtOVUJlj8dQBRPP3
Qrv6UAJTZXIczYuI3Y3AWFThsHeH8zJMYmLntpvLcOGSOgbebfeoXRRl1VWBDafu
+LAFU2OYfbA+xQhW1z8v+UCgNxh576EKglvzp03c/4+bb+IciRAEYFApw7orRL0X
zj2yJvh2zvflrORh96snXi7doEWc/D60ua6IW5qO5ixiFhQwbZ8UmUf/TkNKN4en
2oXcyf3rpsdFiXISnvh9kV4vK4dXSN0odHfTZqGCyl/vWo9e/7YjV6GpuH3ynBsP
eJs0aTlVLJB1R7nmFsTCEnhUWEgLvSgTaGEtaDJKFRswIZi4hEZV60m5t7MgUH9w
DhGVb/wXPT5Qli4QKgSGMirrBmRs50AbUR5KCCmXD2aAJoRb0XZ8c/Y8V+BlIHxS
t4dwfWA9TvRw/DrW82Tkq4Of6mrIKew506LMwKul3J5i437UOGnlujQSTd5OzNRK
E0EyUIDk8/VXU59bzgpw1UrrqX/xyYaEgfUCg+9YgQRDS5jQLbOvwGV8wD8Duk7W
WvcDUkvQsAODla1NvzeExeRp2akjE4kRR5uDW5CED6CoRG4rO8UVC84wqrFdjwMQ
RNSkRB6miXavwRfNuR0tIAfuFvR4bQTPXVM6zXEqAxFQhT4afwgu/sNPeJxnTpsl
eJti/51RU8oP5aOXtsanZR30qxTHK+LgjukgqKwE0qyuexEgGVNUPr7hX2MrCa5U
EbQnyLmsuE5+t49PT4/qLlD8WOQGAWcj1llbc+agENApt/8BElfMob1pchMIgqxg
+6vuS8bqOyr4io5cSHhyHHzbe/N1qe3NnuOI+kBFVjcuwiTO1mzpb+FkM4X9Tyss
+EP50eCMUbmQp1IYNUN7xZbDNfS4TaIeaGVd+DYWlKZAxn3D/7w6PYkh8Khk+YGv
Pp+NsVXc0R1TC5C4aSJYzI/q+K2Vb0DpYGqwwzNpSw24Pbkpibb3pkhgAVaLWdJw
W8f2LvJ2jSvwdRjHhn+yjuDbHMb6p5BIMaHJDfWHESdWwbPSLnBMITpbgT/8uYsW
jq3qXe2ZUuNk6emkYvFTsbBKz4ScU1usqvoIxkpq7uVI0IqVM4SNJFkZp+MsVHNN
RqfN11LKCU+bNTrHMEGYnOROEHof+JMHuTb1GHR+0mOPmz1X0nimYW2wKFHESf1A
Au+diEJL+2p2lct3k2o9IANuCna8pnRQ0bELEeMkcPRPyLu+sdrE55mCUYMmRWyc
vw2E7xSL3ArQm3p+QhHMdKMTdmd3sxE7bvmBVN19yq38JAypX04AieW63nEH9Fez
63GJfSe9JhXqpdxL3jHTBhkf2Y1uCeh2JwD740IlsNld8avNljire6X2jMoIHdue
BglKcZlYf0AS49gke/BjRMwt08M9ICN88ihrNpxlY6K2qBhzic/nuDjVW65vb2wq
a586FPomTJtXmUcrsI3GqdSp0xT0UHe9Zelj/hrDwGj0qq5olfRxbO63eGBRYZ66
LjVFkY2DVvT7FoBZTrewxh22JnvU31JQ7YzJcIKHHA+SFpHAPVgMWNkZUaHHuAa8
6HZYKrBGuvtksh4iKGFiFiHgjFoxXhFP2qNwt0jQDqzTwN1KHYQzYncOgfblWaGS
q9JNH3zeEpa3wUlAO694ETEPySvD5XLbAizg3zYuJJiJONkYWEuXvT/2OOrEIQfZ
b481x/yXws5kcgTfmrNceYuIDQ6b33Ne4Fsttra2S494rUfxi3Y4Qi58DMggxE1T
D89QD6aC/WsC1VEScE2NwITAFdWGl+ZGIdJDrM2kDbZwOdYs36u8kmIAVbV2aAqV
5WfYtOFLMjt/OAnlMiuhYWWHTdpwtMAN/7fHvQIBWX0yq0EKoJsXblu3XVpM2/oa
PjIHA0vzhDcNqFRGgoLOCnruxg0I5VwT0n1ymgFsvSm+wgMZVmd3fNZTOBcg2MW3
Md8sN5KJzLFQlLv+kIwONsn1HicMpAl1uTn15X98qyHm+zW5kwzC2Fq3wDwQUo8d
ZTAJl2w2q6etSb6XS+3tpUid3MgeRQfx/ODbQpbMQ9erXg9e9ebwDKBLPGePVBLL
J3disiBe9Ddx5Ktr/mNDc9YgPdXNCLPETnGaz972et9kQb0VrsGLUMLs8zvrEmX8
8pjrM9TGtF19vK7xsepHR5PgHr8ECwvcYM1mpGtwcVvdRr/qb9cPuIg49jQ+Z+fW
0wXVfzVVcFi239IHnGAJrAqGy4kl0euJfqiGTh24ScB086MbVIKDTMu0tkWNIrE4
JDwCCwcJFnE0NN8nxE0ynk8EKAnwod4NxTslMVEzwr3dZ/EIuo4umyW9ShU+EJtR
mfybc02aSy56cxhvHuTfg6s97KXy/rB7NUgSHtWWa0rI8WOhXVGnJQGNji4VyhYW
GLtk5r6GX/DMIhuSKFFhWcFIdHk31ERKxXZg/+6WOw4ZLOcVrF8GuTIgjOys47G7
6k10rSGnK6++bfGaG4OgyTlHp0nOHwSN6v9UN02feOKzjq3YO9SWxjX8KIr6ZRNc
pA56snYQ2fYe+4KoCEMpCavsPzaH/iAj8x/cI97yCFbGyzJsknpRhaQ68vAJOnBB
EYTiQEi9lBc2ofRaLUO+Qx9Nsa7NWe4RkXvlIILmf8S4oaQfy43QpRLRmclJ+/6E
UCC6iNQd3xZRWTc15qme8LHD38ScpMUYDVQvH8C9TCh7NiW1Jl6OEZ8aG/XI1xdG
mfRqF57EZNSjv8AtUW1mY55hxvT9ir0vknvOJwbhZLeH3jER5QjGLoFk01G2Rs+G
ZyG3INQEX3w25BtLGxotxrYArR6KPXejFHWA0LXjX45Q1sBfiUrgvD30MgmoIARW
03RjM/cJb6OQCa6n1Bp5FK8XqmLEf6Q9T0bmovQ2ZWP8AKuQo+Pk3B2P86hCbeNM
rUV6n2X+BII4rtOlq0GOYioOxjoKnUPeKpTHMWvltWVDv9ngP7e3vNYQC/NDx7zz
sXROPFKXp0zWqQwsjPZuRuSCzRfQBOpDEFs+o0FBjaMmmRWO4rhL6jFdfGjTLFjo
e79pdiVSjhXD1SCjsYkyewTFn24jiuzeo8KPuK+qfrl76MdL6r5znEe8rDzaPP9b
rxn/PRc42YNcmIMhUYKEJzbBcYjhfVj8xWSDtsIEbM6VrpTKChwyqG1HRGF0BW4K
cHirZIuuim6TdDAr/1c0YByDExY7wnszClVHJ5ao1pCb+cqB8AwWDAcVmmKwiJVH
UhvUdatqnGVwwbJLZi1Zxit8GKEhoNbdDgfnDUcqgI9t0ovlhm880/L7Styl3G11
jdX/m349dDS2cFCHOjYfGo6Rp/4yP/lA42ezzi5p1kXSO2s7+yuFpcjcnZ+2AKH1
oAL9YA4Oyqm38A+oNL3LxDEh6Bq3fqbGaWKXs7FOLE96Gr+c9R42U48UfJltmsi4
kPFMohO+ULZ2Ivl2JohfPVQQNQwcFFUgQUAv446hYvKtL8LjWAJ7wQ943tut56KP
SUrgCqsLs94WNcvrcIA4TXSPOkSIA6qo6C1qAtjhxQdrDtqLUnQoBgca3S/ZBG6R
V8hIRJBwo304+cyo25nbKg32dwYjlTiXXuBfv2xjOSmEcie/XsZGNQT73Vccqq+1
azxOKTCvw4QeQLxxdj7lOxBBNL2pDKS+srq+3JlOCo4ONq9EWLUD87pfFuc8iAiw
ymr2uRRdj8eV/mNxg2Gw9jQxRe9nCcczAys4P1JVVtqpnAf+oqQKsRjM0ZI1rwZp
G3XirYGwAnCgsNu1DHTfVxDGaXinKwf4elZXxC+pQTT91Q3nd9AvaB7iRTVhLWNz
GDFkN1rpjSCh5O9bSXqQNEHWEHZ7pQqpTpJ8Ra0JrrobdUWdy+gw3WJIzSkl40kw
mahCOrdi8Q/tN2pkmXLF40CKUrz+FjW+H4vPsaF8wnosrK6UjPTbBsqTrS64Ys42
o50qK3GrvxePQtiGRHccqbxKllPmQwPSHDYffeQQlHBi/MY/5+WI5IgAVeLJN+/l
tVcjrhzWvbZd/BOnjSSQ2foCL9rH4aR2Czj5LXF8o0waIxhZLxVvMvKCHi1cN+9O
Yix8PPPcVeJ+OVPkpEc88FsuRBvFAlAS2w96iaEF8dL/VbmEMLXRBUhXN0PS2RM7
J5jw/sNuELU8ZunP6Uq3atxA8xEuB4RIRwnkFRqRlfJV0YT0xjoG9JIvsrF7z0n4
t0WhL99XJq34RpT/D8Z96qNW8HquCRU43rXZcRcpFVcl5uQwrWe08mvVRziQAx2x
2tRryD6ZWj9wNy5IDJBe7idlnKWTc4NBVJtpeuokDYcbGSni9nsv8Qz7XJgrgZbw
g6BncoNm9js/VLZvH3EfTKe0U9K3xS3HEG+6MIAhcnX6BQ8pKP0B0AW3g3T7j+lr
W65lPF+ely8G+h3f09q9ialEQlJtaGmgjKVfdhREOZZskkrEGES1rVspCiLgOrTv
lOtK6bEqtUqBZ6oM4Eft0/EGDPOC4i4d0l0spPkpru3hSy6NuG5RgQy2R9PDiI9T
l4EnUb0fRub9iXcx7qhAZ+yqFhiRyhDXPqeFaVUw2BLQhmThVbPii2Bq6tSWD1VW
3t+VNQV15vCMYoqJDFzRndgjkO+pBB7YJX6QqxFo7o0NVCyeoYs265yfrJMdDGB3
b51Ald1vFLgQ4ZS0ItWSgA/o24Twn9G7eRJK9nJs63R/566m3EzP3ljl+UOFigfZ
AcMRUIXiiHZpZjMoYZewyUBxYe8WHgwGF+hHzmESYTcPODl1O3O8gWmwmW546muP
+YnQ/MHIQsHKBSpIA6Z6A2fXDrJC1HQokZN78UtMkkjiU01t4txuxlAokaPrls44
eQr6yCZoTwtJxkSJqQRcZbn2kznnw6MDP4H2jwY7OwstKDj1+eF0nzWBnYTNyadp
11f1tNTEiSn7G340RYl4jlHMBEoLNP7iAx5rTtUiLLGkv5bJvgXSpeQIN//g324j
FQNCNsQZWzOglIG7UsJYR9cCLgXi/ETbyKAkeasAAltYrVs9glAWBx94su0VTHZk
rnl2pZ1RTNMxPv772X/5E0G5JJEKAzBDqTuzROBEWUGMQvhK7aYj1k0iq0kLDVQ+
2mShZDPtOHVheB9NefZFalnfSbMCCPe335u+cDsr59ssI0tsUgmLk6yq5rfTLITu
Yta6imo3wTnNvFpyM7wYSfOBOFqRLwFQe8lqMjBJKMaao3ROZMbiOgvMvA2qHOhV
c64BmGDMr1Cdn85483rLHabBe3K6lHG/jcJPlc3C+cXLP0avvwBvejKXooAwCzzt
EyAeEPAl3LrI3VjcPE8X5Q1GyWuBaHu9mIZwjHX+JAE+zTxC/gTydl1nY65MztPQ
BIPVG6pU+IVEfOw5uc8J4pY0j2HCCipGjEq4IoBrCKDW/FccI7nY6Xgc6DckTlZH
2NbV54DRXkz01jQG+DdN5Q1jJstPbOt8WbY6BscLK2dXGV4ESTdDtHBrMnQpxvUH
xZbZhzxGXOwGoKIc5CJ1Sc6zW5aRAn/boILisNGhi+Y7Y5iw3wSClyL0vmtwId+x
9XnxKg+3ROcePIalLvLWShI3GUwGSgp3YhT2nUUrcnP7ZIoFAQCeLzXA9JlvXIMN
9gVShVfKyrEUF7ccE1+8GDjW99Jcga4y8W0YrgjvnvBnyfidpN0SqETLHOPoN4K4
4Oh6NLtAkpggkGHwyKxJ0x9cVyHsLyeaLArRUknu17AVvd7sw0AiB+tkJL/LRBTk
HiR78+BBBq0wtWja2oer2jBKoN//BV6/FJpXaiDkjysnLtJZLCON9CeByeF8vrRI
a3HfIY06HSSbmb8QWzYE8c9iBgnI9p60O3rQ/iKUu8aoOV+ZyxAOloahjTsUSMF0
10wFIjorj3CV7pr312d12X9Fp+fVqYzoltsnFZAKahcj57GAAEpVtb6C9sBv5WlI
/9ySpa+AhV04EfUVgZkw835Eb1mc4btK9Gxf3X84MefRJ4iCFQRIIjBbn7LKF3n1
pkrnGtqrJ45OV6/J/LYYAdAdjZpgK0xgHU7EflLQYt4sKB1oZbZtIvpCiznZ3U1n
ypk1k73yNPPqpPcSCFZmTIhqY+FQS5f8iZm3Eku5HbcxnfFVqqd9YpIHmm//+x+t
hsxh4plhqjdHOFJy1Nqm3Hr5+IFq5aXH7rwzv4R/I83EaKMufeLwxmAo0PthUgeg
BSRr+kolHELSfM83MSVMlfHWvv/Xrecf4DO2OvDdQgWFsXqztIc90v+wO+N4e9EO
RhNT6AdRjDaFD1Bwbkfkvs/npDYwrK4HcKJsMeMlLZL4Okn8K4y4aIQH/kQ5/Ywg
5P8mJ0fCg4+/5uxjHQCcbTLG2d51yFde3h1Cr2bQvbinRT9goxLuy9Z+Mz8nzAM/
c73+V5rJMREIiqdWtu+RGYW67w9OJrYSyVnsGum0cUCI6JV2KZ4faSUYLKp3I8cW
LngZoNuD9RnnV+dKAGDIFurI2m43eYMPCn8sTETJhLp6Ss+IAMp+QxjcUmN98aOb
dkwiHyFVOjNNxqwRPJbCK5aPm0S+8hpBH84whM/Nf/PZJHiio324FlmoFBFodwbk
jECFFI+qNzZT6vt/136a6kXClG3F973fepgBdnJVA9zljTXQCkFsrenpJRYQ69cq
uuwZX9K7h209M9TORJdbumf7aDByOcitJHScyl8qiwmFwYPZXB4mD/pDmz4waflo
ahqF6NpofKV7LQ3pTmNCy42tC1rqQ6hmdfw+CX3M4IUnypcM+agjjEbAUvbeyk1x
v74AssVhdY4F3wQhO676TrHNTnvEQuyj9twTqIEM4DiU1TDY5XRrGJ7oAJnsxyNs
8d0h+pxJpw45ZpkgsvBYhYGehS17M1M4WMtPjz+9UJOdJjzYd0WrsfIABghtCR6j
9ku+1RrxZfDxAi2SePeORPU4AaheuJVKVLjvqeYAHthHMUjULoRvPbneRyqF0jzl
VjfozM7+3ToJW5QYl+qMHdD9w6aIfGKRVjXrnLxSrnx7RbRiGoKFQISJIlRRACoX
+Ln4Ri7LNpkMR4PbIZ/X2j8q4OaDJVmajarol42Xn8osJ0QynKXZ0f+5myqryNAV
dNMJw9ppHqBds4at4UUeJkBRNglUgsDQszuVD4r4i6LR1MDdbtkCPFNyhJa51rDD
2ggYe5h8VX9UL8wFyqaFMKddwyB2pNB14sBv2kHs8EdnxAISuwS2oYikfhgO741S
CHV4X9SOxjkhnYxqNaI8dbrlIeD+u0Rwu80HllyyE2TcNkOV6OXsMlR8reT3BQKm
KNgU88jbRQ1bwynQY2FZ9fp3gLnwPQ0K76oGNknIrtg/uJh8UG7z5iXlfS0xbDii
wwwY2VaP4k2vBJZqo3QYf+6n/i9UMF4yiB1g+OeiOKyJSQcndCNOnGYEap9KlFdK
XMDl6+gZ29T5Z5dM35QFImReuv8OdH+q1qXw01cZkhFQGGk0551mExfTjrURjY6V
H2DgW+1znyd4dsXlIVfcqumXqnQvco4j8jY7dBnBea2hNo2/bJRddABwdDsMSE6f
MrCOHTzMqSx59poXPkOQxWqERjc8Y85bu6dE40aN0tLwZWTut5gZibUWjqdFiSUw
rj9Yk8AZv75ea0WpE122fR35+WWR9XSVT6P6Yvaux788ArLF0inQqMG2ovBkePBe
3eqHVy7c32+WNI0feaxV1kzUYKxKwrksCw+SQFVLGlcC6gP4iokFUKAf1xPQAQox
AH+35kF+yiHACqZI2JU09BM8ZoUCF9EWJ1cRoScpB67torEenZvUHX7xURkLyMSU
R58+OWTBRndMPQU+uwZx0toLKPaTCfzv6Ig0qVAI5qbRILmAiBGNCQVn8yeE/bXV
JX5C2/Y7ZbK0WGeeue8Y5t+7NktcYOaBpKapJyHpMkrblHVstrXY852yxdo9/k99
h2Y3VYTW03Q4NTkUUkjYHaKMsQNydMmG8GrACeOHOM91Wq3AKNV+zRqJ2s0sRiGp
TCYDYa67geTnfD3ubceOF/pdgMnRl0fS80vndRQdnt7o2IiU7GnGZu6wKiUGkxNC
Yp55yqQjA9T0jHcG/3WqTpacBCCe6h0mRf0SyHQRienNOxD5RVpsq0Z4jiK2vVe/
vQVETie9/jHMYN92uUysTgIpRe+vfV/uIpCUJu1qekWthd53ol+BQ78zE/eounRS
9LOevbiGsYYw38rKMJkbJl4DT+KI4IsFsanoQ0HJxt8hqqtdua57dkdzGHn5RsfK
Y2tlFExZfKMjGBraI60uQPTHAs04zLm8Xo/4Ks0BB92+TJPqFTdxgAq/BbTXLeBG
b5cc1BJBJRJnZdAMH80Qgfbny7ojifco8cpN/LXjgSKqVWMhrDLQCkdWgkRCyG/u
bj9VRD5QF61XgIMXGXirTNx156DuXlmeIyzLALysp/qHTPLxHRjG4S3oZTa7yUQo
aiyKngu7FDcqS8duu3vTSB/X4FkrUtrtKMb+mQKOJpBPHXW7f00Uxyv9hRE505iq
pDAOUlU2EvhsjrCjRwW0pR6Ia7NZnzDflRuB0tt7FalzHB2nRbGZtberyWJn8xC4
X7eaOVaMSP/GvjDWTonEyk2AaGCVPDPJsggbpKKxtqCfqTI7+AGxkBcYHz7EMgxl
zorYn1KGfScgjsscQW9SHI6DE3zOBnHe+K420Szf8dhfTPADbJwwMmzlEXiaGaXg
am8OlaESxq/VWtsu57Om5AWe01khNwmpUNsHTJmUuHmXl5yYr3Jj7+dCdCx7bF/p
9vm2RXs8Y9E45bP8R7WOtfrry2n6T/ysrMDxFr9AMz5ILA/7b/dhNwn/phzXLN+p
mf6zXk6FgdNCiI4FyeFY0l3uNi/vsXsK4UsUVJd3CMi1KvqUQX9uAgvARZZqlhat
B0kNwJTJ8qqyI8i/zZG09OBsGz0lidZ8A/jFQUFJbtIjLINhOpbr7oGF6+AlIymj
SntBsGoRJzOtDk5mq2W7CzoBaG3JdYzCTCfnZF7CGLC4oBZDVbVRXu+n1iB+iSmQ
0g5e/uVlBBVB3RPe6Fcwy5WqdENvdU0PqjTNO5XqnI/uSvvAcDSUBiGJtimerEqL
mgZND6TSRRmbHhUrUy7L68Y+DQXPVHveY3uVsX5Op5WPyl+8/Zzc80CHV42pUILg
1WB6EJ3Id2A0uR3Jj6Fg7OBtOx6sCUDUKH078rAy/rpgZzeihFN6GjsWHuoN7et7
wb0JpXjxqPBLXoClvsoqgjUrRUSSrP7vqquZUn5Fa4KNtJJVacs4oOzYqTgyihPy
PpO4gz+SL/Asg7lYAxEG8l58TZWAdycMHpwx/aiWJMALWg++XyPivqkZEloQaFYG
m/4bggZNB86/PnDMvs/22To7AlVDvPWHCjCg9JBebur/XvWki88WeBdnPH9oqCty
JuEHDb0AMB80Siiqt/veYKEREy00UO0ZCCdz0kHakgFdogaiP8CzXwMnalsvAXx2
BuMenXLMLxftOjn9Y2xGtw==

`pragma protect end_protected
