// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qtxdW3mjaKiwO9erYJZNtwEgSghxNESWGwIvdQ5dbg0xmdch6XXkQRzuqvCGL0WMnwmCC95vQ3da
jh/S5crFAlFe6NysBYaKJh902XHDH6e1Oaa/YNolOhHDPbpL3L4rDUsnpG2aBiu/ZxIJCse5aGMM
OMELZ3y11sU6tmLTHFXKZaTPXAB1pO2qFbBpCz/en7p3Su79XnxwTgjzcHMoN7ooCW+4cDrKPbFk
MOGqrSmWMHxCtQ56rWug4XWLq2FrCWJ+sbTB+4sv9GoEohHzhIOS7j/0HzlhytGHA6XPhe3R57vd
EtBIWGs96Eqb8gNpkBAZx7Jn/l7/iTmuPpkbkw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13008)
VmFWaeV/RFpyoG9vZEu0QUclVGdsJSm0wDh0bdKoDW/g+85rEdHZlSPYikOIXawodTxye5Nh7d+a
487x9700HdRQHDhM0N/kPOdmw/Dqq9gkufTHxcOy8fwV7OMODIewvc2eCj5zsErsenNersQFkGzA
ypelsVNJxrLgEipvNHJLlNPSfME81ddRQhMS8Ugv0d5cWtfElwpNeZ1eKv6ejCBTTWrrvQz8a3wj
MpGnkFID4BMZOIHpRp0ev2tVouApW8qzc0BujAkONPapj25zgfCLeI21uQFMAi66c5QolVzXu3AG
vPPPpjDKwulsEJ6xSYhBBbfch02JVhNoGPgAJjZOwquhwJKVXmBttBIZL5G5N121VYPq+5DKJcWf
QdCMx6dkIJvzmQGQt4aMp31ilceNaooYHufyMV3UhrtoHHiOI/K215DJsL7K4uEDBUcZyI4f7POg
LUaSyNAQQoOs9BvNXXNiVvaULnBNYgLRsu0/pzRtnu/50j67HGN32efXjpqPVsWd12djgQpgFUIs
vHTYIZyWiZOpVDv+JjgAaEDTzFTKRnYOjPOS/7UVhdu2vC7cLSMq6PhkAEvral54lO1uzbQj4hH+
bM2b49/Xns3cc5V9+GBgGfULuJENs38+Wu7mnXqhZ9vNcQxu9Yctc+xx/rEu1UPsFITQCAMrqNhz
8rMu9wFSXm4Lk2jHPkTVwuyokEVxBoLfh8kEbiiYaieOOE95zlInUvXsCqicwuxdzw5fhnDdNau/
e0Kv/nqxYLLr6W6mut8GVsYqJ6ouQm2laDJuqp9XWAw8vhHhCQ8mQNg329hGHeHILI5jH2EjBL7q
4CnOyFzEHRbtTB+mqqE42Z7+a2TpEgjPBZCIsC85yO3i2COZnUFimMyyDuLGjMOu6zxvixH/4jaJ
1k1tKIoy2Ht12SoUOXgbzyNLn59RebIpR1bjpx6Hhft94GVWWIYz78rcTa8SvD6sBOLPMI90cuIU
TBRiXOgSpHfF3bsvT9E3PTnMj3k7dAM5nOs7+1fxawJ8w/JlGWuBGiI+e397IBR4YxEXpswe7kvF
kzhFHgpUK9cbiA20kNOKUEOiwSEK7RfHsJSt2OZvcVS+pZxz48+epHrvGMaLTOYRDnDaQppFzdr5
CtSNU/XV2zLot9KjNlU0hUgmqHAUUO4RYrrJhDTKMqUSguhI/ROneL1NKvZnNcFsaQnltgfXhcSR
GyVOto9q6dfX4GMFQALy8QQeLfIPDiH3mPhxV6ULvZX0nAkGl+dNqqewr4cypg8KeDDNqNnlkyL8
+ynwud1BxqPBUDl6l25C6f8KKFV9Ow6mWJ0/AVuppmcQsVUYSkqG5IHpEtSKrxY761rbYsBIf5wG
BW3ilMK+pX+7GNZ7KLgEOl72gSVx65CfpgNMJKOQr+igyyrXBhn1Bu12EH32q/VJipiVYqgoggnS
afzvbRziZ+tkekd+AL6aNodyNdfL3mMWTf8YTNLz6K5Io6PFvEbJJFEiJE1Hq63GXSHjWm8ggrx/
Khuwh/TMs5oqroxLAOG4x9qyeEEwKzt7qqvNuW5GjchM/P7jV3El9Xuz+G6Mjb0LGkWnMB1Zfczy
V+Vax8zxh9htNYVVnQ14WLDaxA/Zy486EZPgxdes85rsLaJjUxMhk057YJWJdEATjCUxPLMpi8C4
uNUbyZIxBr4XMm+uDHh+aNBqZATVb++DquizGeH/+CCwqT5Ko32nD+AWAdY4dtVYs3VI7Tyhb0TC
/rZmdcfvSFBlP17Z3JC4jJ8VYD3B8E0ehIZ3DzVUmMDO3sE/EzO15q4/FWLQwOe3E/lGEPFcwQdG
BQfjrMTWfsIK8jIfjAblPOMMOa1LO/jEmv/ysBbhuoX58jBXda7cAXZQjf9dJ3FPx9dYroc9qDQl
dSvjiT5fC2HF/JIveKeApJrFtzyj6caAi/LnQiyFM9BEpesec/khFBBJe9pdBru5uwCL/Cc3Juyg
3RLlIB14aW/6aYUu5ZhxZqkcBKKPnNrjHqQ0NQbsn1ZHZgJfv3x2mut7rtQnhk43h1g2ytOzpptb
UxkbnpUcPFjLK0AviLIV18SFByfT+crPouRL3jg9sb6taZUWUsekYc/N77EcsfQTqjHxazL4Zcsz
UJc7NIvvsqSsaZcZtEeXZ3quxbccQQLaTbVIud/kZVRBYV0hnaE5e/0SphQlP5V20ISV/wrj0Ptw
i/kgB/xXvb3VdGg7QoYkWsEIg3a5pl+2V2BDa03lqwszDOrmHlsa2BEU68ibJEBSBEiKkVL36ez8
UCO+zylk8oPyj3ByPIy3eykeTGSz4gtG7SPszl62cwYYJCx2sEw9EZ19NyakwyBIMOLlMv05hjZ5
4ABisrbZFqAvMdRvReKt0XatLzp+xh7B6Vy/Zx2URk2YSU7eGzIEqpvN+LIMmaX9yQnbDN6LIKKQ
VgVxAvVfD/5QO8IkhLqaXP1D7xEq/bBG0r0hmJClg8ko6PSTr/s/YIB3E17hKpWotu4FIpML5bzm
GJimxHHgG4ClySDIqrB1REI40ALmSnZLXFcWBNdmcEl0bNOyNLp7houJdO0ITxRp6dWbC9Id136e
T9yq9LVh0ukAehpe5nmpQuWipra7rdIb68kEhup49O3woRi5Z5dQJzxlxVxei26gTC/06hOaZlbR
7VonWUkPczOfUcLPkU5+2z5O7QCNvE6RHHPjn1zWyeCbzXykQV2fZ4wmyx9UoMeLhRGrvcf7xH33
oii79sCzrUKF/Fd6Led+pzYMB3RZKrZRXY5TmnLSc1l2sSmqKoawuqzEqiPpnd0Sn6luqq3ljk1y
LVlNki/EBoPsAjQdQ4TRwnXK6BkIS75tdHyURtMsNj6RzSlL5k+d//Ycw0L+4nOvpMhe1JJt2SPN
toWYlL7S46AzqHMn4PrNURPmXj+caJNPtlS9YZECeMOg++3GM0bLrQDpKcxIdvxH3HoAENHCxRnT
vGzs4l/BfYzy39PTZn3liJLDO1/L8ucGgLid5a3rAj/WVCbZ1zkbq9cM7xLsMgj7V84IC2Za6GYQ
fFCikw6iUUYObFrBTC9i0/zjcTpntxWOFWFFGrueO/6vr5gvpHnA2wuJZBLYvk1Q4ali17wcBhm+
+ezlfR55Dy+Z+jtJiGq6aCpGviPsWr/zZzLVKMMNyUj1ctoxFbhPo2G25APfi4KiFS43LXCYHQPW
ie+AMY1fzVfmouQlnxQwGsiNE2mZDOCUGiYhCjlTFPIx30iHZRPvn1b38GCeZJzZ6pGH4v4cauBy
vIuLtlYmNtH8eMoFoO/BG2dPgFqvr/L5wuR6vYY/jdczx6vwMqFiKaj74OulmuWwiCgcOLtVLLr1
MForZVa682Q1TxmhziThJzbE/WxdBwijutz46UeBnNBpuHpE9G/UwgVUcadPAaqBYUzW44eUgnxA
OIEB3YGle/k7K8l7oLwqI8u9U0WuYcR+vTXfS5RsByJJyYxJ/H9mw7nA+IWRwtCi1e9JOUJ8bGhh
RfsfpHKNxGN/FRUpbrztvjsao1R65ztWDqmad14B3H88lV144DFitt56LbBAwqjqciAWglJbTdPm
cbLcDCY+DQZCuGr6iKmM7QOEeUa19RU23eNBD/rmT7DG08PSYwI+xE4dht4bru0cylHcAmDQgBYR
IVNqNNNbpNapYnF8hkECY23bB9ZcXleiWOXWvpDncbOekz1iok5987KO55yyDomzryFCAw85wovu
eQ2ywT1Sd2qrpANoEh5wVbM1dNqL4MCtpg62l5FWAp4tlRDazJEJ26Sdt/oZF7QQEGueexDt7ZmL
RNaJxqxxuKizObDU+lPbbLM/iULRVS+Lmr2uP5x6qOm53Ht74X4IC1bmpQSBSSXwOTfzSbDwcPkr
YBiEymRrdMWPwfHLp7HRcZ3QZg9ajigATdwR8WFDiQx4XLv8GzaQ1tumaCYG9LJ+79AeH0KiE9T8
hBuS0bUvNYVBIfMUhiIkrrT67P3zowUg2a0Tsdt8TIgCU0yUv5tDz4t1hBQOBQD+2uD5kr+mAbts
GAIri/Nvx/1XOLWnbvB0IRQ2obV62VBIK44hy9+q3zCl3NoFfurYqmQDJ//CsSpsJ1awccIZtWDS
x0calOLc1JoP+qA28db3xn5ENYyxix5JHvddI2ddrVHp3rHjsK1/cyd8zuACWKeo/J40eS3v+snU
yOIB3cK783PwzYtQcP8uW73nFCYnPEQaFrPobEfrKFIomyjEmTeX+niwW5ONj4yAO6MZ2Lnj82Kh
l1uxmK+m+nDqagmAr5PuA/VxiDeeRn/aXVgDvkgyMmV9XBCbpgIq28m3wMHm7uVBRU6tZ0umnfoR
Jss2NxjsX5Cms41yucXIIF8Yrrj4AWwAtgC9mTQVMt8h96cr5Swmug5VIP9GUEMi/zoqksV/HOAD
tWmzjWzs1JoU6K1XpFAMA3KthkaRebjRFGqGv4xCGhTnV19MeG0QTyfgDKNl3KJfMnVFMdeVTxo3
WM+fEOIH6aujgJg3/RV2ZfoU+MxYWulvv7pxR4Qu7K37J4MPgnUCclfrBKjCkCPwXuAp7DPjn65y
4hS78vOVeldQ9Oqa25wGSkadOEOx3tohI8DLJktCXYthN7jnC8q8c4f0TtMJjIG2h6WzwszYxnok
35eoa5/UcJjyZ4G7qYZltELjeYL0kmqOmYC6kFgXKu0CJTmDKpt2ORez52rqvJ9PbGdTP7QFxCEA
TjCtc/syufnF1RvFTVV3jW1iA6fpXwwWa0s/QkvQ7yCN38tB8NNfB7nbVtGgvgrvmYUvVDelVfeR
AVPkPHfGyqk0iQk4+P9E7IO9mev1kch3xt4jLRqzC4mxeOb40W2nWHOoELp2o9hGjseauVFsnz8/
TAkvpCmFdfx+zl4cRVjddeXuhq2GMoRC6caCyxuM6tHpBIvdCo2/Xien5hqQQ4YnULxX9t4uqNvR
qw5U5fpMVk9NBDPbzQ0uaEhnd4j2v1iQZTDrIeAGl4j4TLiSKAOY2OYnYAXtJhUaLTuG0DILacNn
bWFBJYJbXTNc5edQTF5ICNR0xLcjSTQbYQlEvJg/OFJIeBnmV3ImNBEpIl4LOjtHyqepoGFKd+im
HQazZR4T6dWXZOdSvZSAqe90pMUNVxCjmc10Gw7MJuYRJ9uERkNAdAsC4Z8FS7Au1Ojw1G2seXmP
+r3H1GMYw2u0CPDJS1GqvH5FyUNtUza39nu6zr8khCTyjUwKVvdouJ8iVFzqyBLOV4Edv9BmAXAY
/hRiaPQ/0LZfodw2EWyMkc4ziAAJ640nNguhKtEAyYhFNWnC5rZlyhDYFl1g3ohsW3TW8WuAhR4t
9wECTW4wi2WKlwuMG2O3TjLZ7TBXSONNDeMzRV0iSbtdij5s3dlFqa0NWlYqspJEDZpGQDK0Ljmf
l5iY6lGnJtuEKk+AfhWdvxiWxV7J2/ksPPxDCW1wRwzQCcGYH3qZgh2JvKkaU8kcWDhdJJ8HmTOj
lRhasmxr5n4Kjz9G6K9z2ZSxkpf9QLqX0nD3r0ftG322gO13LwosDSXulTALwCsN9gLeJbQtxh1M
GAWlHU6jdq2fIeG6teV8HcG7cAlbjPUQFGnp9QkYf0Je2XFtN5g0PqKtT5pXHPHvgvhapBqTLhef
DE0CSFy0hABpPiXwq2CgoWwgfBlY5VWq70X23oD86cBY/3Xt0PL+Y/JmViwWUOP2IXH8HepNZ6eA
u9s9oV8Zosfvy6GGIpoWaIuBsIq1tEKly5jexMSWHGNs1xPYIt6pMIGGvVSIR15yN22EnLMA/bgC
Znq4nUJ8u12Gi/7YRR9EPZ0VzV/D5DMei3ObuhxbkxpFoowXTGs04M4H9Jr5j2Q4id0SSrqbpwfd
nTRcN/7q4snJmcbLuI2rR9mAp5lmdtaVN4yGWzrnMUtnM4eNSgbaiRYJozR8vdNKpmjFJrU1S0jo
pEfPUJ5PnuXU7m+TulSLB8KFPXARTuaqe7vIaESifPJyjkifZrkFvSNRTiFDymIpFAJ1oxfJ/r2z
itIwJOjjT0AANN+RVlOucQjziIHo+Hxr1xyB1Kc2blr+bVVKEPY4rO0LRAfNGS5MPMDWFvIkitnp
btu8yP4+ZdFB1GuoQUSYRTvMEiIIiKwOYKxHJ8wKAZtEMgsmHau+wlOghAxafqo3+wL9EbLAQtUS
DGVv9Fs8IYYa16kOELArswybaQizfMe7nk3cWS8yZCBGAP0CtcTbr7J3wcjtqvxG0XJJlgz3/2lb
vCEF4HOr32UsLq7ft4O+w+FvXmdL0ewbILWJKDH8skt8F097ujxkX1/Y0JinA1aUptUY3ab+H4Vz
zh+TxEykVgJIHeO+OCLNa0vqs9DYtOhIs+8PGGPWP/mFUxlksUZfgYY453qk8tmgMmn5YPHlGgYU
+6qWJkVu7/jjyQz3oKpOuHW8tWjWeDTlYbNQ/dwHpatRWB26c0oyMQzyjUvdWNuvUhBYMcAWkQ38
Z/XGlXDeUFVGM3S4jCCONkYrY1sFaWyayr6rmx1/ww4wt+FsiLSQhGscqsGCWTH8n6+a+rRiHlnT
UOYYm37rz3yOY2kcg9gNre1OzN8Zwk7iu7Z6sqC8E7k4hCYAsKGP/K0LTvkwQh8HLvEvi5py4Kfs
V5jFAA3diKLuMBVmXY888fMVQfdgU50i9z28d1MT0zhuUy+vA6uHU9ASs4Ab+5kuT1/VLCxDhfxa
dPwtsfcIhjMTox8qf/HkO7B52AxXoptNURiG7eF0fOAu30/Xz10sVV/Lqg7vC27TKEX8kx6Z7Dol
bAwGkSG6RRlh6TFxVQrvg/dmpCxTBS8dVckxFzN4LmHvHE6xXAv9K1/NYWkyUenISY5ZXKgtZCDs
m//dOZNvhvpoKJ6BzY0WxiKnCG46glC3v6uJbNRy83lAo7GYGx2bPlGULg10U22gouKGys9LmBr/
Gfan6sIV48cc8/Owc7NIfyytnF5Io0wWJeiMaRidrKeQAXgCv01pB0fo8mXFOvBrFSZuURAR9vR3
0nmNvjP957h1ekBxstMIrdI7NVerTVKrT4MFmTM7zmwdBkFNMDQJdOGPR9UWEP1oDYSQonPEE+G4
JZL1LoWsnmq9MTS8M08Nu2Vuk4kE9f/hY7Ech2EFLnudhr6w6eLaJyDq+FzqdcO2NZNdy2SxXK2i
7eRmS89/KGV5O0PeV2er8UmKRoyj4he19J0CN6a2fvHsE73T050JwtInYonhg04SqdRr6wy+a3Y3
amqo4bcNIahbpnpz3pHzdAL+p/fOQX7qLWxITx9d2E3tWT6l4xJPVTYRgQOhn2M5NB7cWQH70q1r
LgY9yIJRMxEWHwqi50zlRtsJKKLA1ri55gQ2aX2IjJYgZHRNcbzcRIYQiSE1bNI4icbcEjxzQdG5
GhvgJ0NGVvPaDAXu2Rm3sCoSpzDv2qkknYoE3b/YPU6qhYJr2fXkobYnFj/+Eio2n83hTPT50JGs
TPD4tfGu0KMES567v1soU2RW2MWwuqEVbpgPulCI1zrQ4V/P09V1tgoEYekQWxZbBKhRibWoh6NF
lTAA08fRpmamxtPpNfVfYlx//P5coGV2brnMnUKXaxxpwVsxZeuxNsUL8LaOFfpPmBme7QC+OWb1
t2U6eihKdainXBtZCXWJu+sJQBlupxA9s763A524sYKJOOOlkD4iHUkmsjm2uMXn+eY1t5tTw1M5
wvSdJP/a/5oP86YmvZTV3v11fK234ulJGC3DKpwnO3xHPDfuQOl4qGzhmRaWsd1Gd/SUn2vYKt0U
+4aYkcTYBmW4w1TYw1z/AkTPiRA461Xcq/R4dbKZuNjgy3HfctnZkDovpimP6w2rFOud+i9CVHoe
ovuxOogKxs7Q+4M3t10tInZNMblAsKWES5zGQsNCKNl8D9p4AF+lQg3sXmT6DICu34n/KDQKcOgU
VNLBHSgm+SwC8Ry1DLJSxRMn7ke/cEZCZ+ZwpA++FjyJk+mdpuGjHkSm1iHwyt0z05pGbIF79DYx
wtfD8nsseWwBbv3BftJlClebjeyFxw1p0TD/HofvrttMJbH+9qFnQ/oixY3CNw17/kGVSBZU8D+I
pBN26agF6YqKRFUG/qT/Uvtmo8XETq6HGphIiqsVNpy/QVQpxmFF392/3QAmXtallV0j3v5JdSfF
6qLcPJYI1pbSpLowVHknt7TylK3/mFjXTZYn1gOMYDg4iYb2JC/Qz0glKUsI0pfPNocw0uFhybrQ
1RwxsyLueeg6JOtgOBkKe5o8wYr81Tb982yZXEGv4vP8mz8a/DIzoFPs23lB1SZhFOJrVa91NFpH
cnlRJG86OC0eTiQ9fzwghh+YqiaiFTddxNUrvcekQ71nucQlWQeT6AUdWfOyPgsolgQoNzA31Kd4
f4859/jOGEK7ahMQ/dcSEvG9ki8akzowmPcounNmGq7Efb93Nl6mF6JmOJiZszZ8XS83oK4ux3Vz
i8/+Icj3F9FYfO0wLm1YX/ooLgDaKtpQgBpg3uJojkY/Mvp7zl6W2nWdryVc+ZIJYy+QyrV9k00k
XLZIVJ0MnHVYIXtAJ8uyLJrAs9VL0JOrVzJ8KaTVQHDN2p7MbagBEp3L0YnSz+X3pTyZE4j+FY0o
k1EqdMRgoy3bKY+FTPrnFaEhFWIRwaUWG0aLIDNyQVlqLwXHM5br24tlDA5zQk2PlR74M4kPJIjw
dp7OxrP68IWULBknnksFuIdiiXeSqWxClDxtsaekyGwFHL6MB8sTzRAYH5jr2AMj5ZJR5jKr9xdZ
cMByi4ZGBHpktEs2QIRDh1cNkCU/SekRQbRf7cxZtxIp/l1EWiVG6WqzsKra4RXg8MFH5h/uJwIw
lXJdju5lmmd4zxkTyQf3QUOGBiQKfShMaHzKdNQHURGsR3Pf5rpH/PBkIkilqqBKPzzhPJRX18hz
oIGk1RyiD+i2LFExwlyYkids42uw67f2gtDIHzVx/eWtQ+AhM82pQ2CLYXYajl3oFffE1FEYgX43
BlInxS72A/C692G8wbiTGSfALIK3nSJRdTl5MuTUAcTGiICoDcc8gJnUfVvFRBpQqi5k/efLRaPv
LB97RlJckweEmHVH2YwuW7E04dqxoTvbSJCQKPn3VyWpJE/M0xErYEEDJELNM6i3HMJTiTwOqE+P
KwNY7NayZhslYiFt+DTcxP4iNxqTGQyO/jSnd8EaTeLG0bC45IDlezw2pY9kG0QmsSUk34W1JEaa
LhM5jxc6FlLKXByMwnXJxtPeXS1fNdOPr8M0QxkSEyekKFN0xyd5x90qqIUOST5cWz8jUbE03xpB
vtui4PuNra9pP5i+o/sJ2LlkN5kR83qRK7yskodT4hWzhuLHlwCyMsuAhc4IcFwSoiYAp8AHKNa2
jdCsmVIeaqF6TB8vu6P7Lrt8/4vm5zj1onni5ATOfNiV+yrjRBrDCSK2aIMr7/zvVfHlBZmcVlqz
GQBE0mlAP3MV1u5yejby5rvc9xe6vDswBAMtKPZT8/EH0TF2g/NdIy23/xlGKl5JXTfCDTUHFfdx
XItdmlfhiA1PVvhTMXuT3Ujw1darFhDY9NjX/GbfLwmnPnTeOOp4uwGcBHqfFjyIJN0wpXJgBSx9
NWbeDAUdunuw4fW+5K1yOc+hDslOEEBvZLNJ+jLsN97TI2eLlXX7TVsqOqBuidKcVqx5eDqvKzCn
LYXD9y4zVq4exiuECaFlcWqEyfxdP5TmJ2kfEDUqlUFKw5yXUIlEvncefHQ6tZHBNtllXcCDjrP3
Wi9Oc8YJkzb+LzzV1BFIwCXFrRx6HU2YXO+4keh9812+hsl+d/cPXuBa7+JQAewGGpkmmp0o2mH8
mLOug5gHKXusVtySyavrvFxoQMyC3WE8OdKlK2BiDubMes5aVL1kMr8HM7HCgAqEc/MnaN1aBcn1
qI+a9LaeODi3dJjIA2k+vsgO8ZsAAnhgSaSwrxTtuXVdIJiVyi5pcAGmO/0ZeOGQpPnLWbt3LiMg
vIGIV//+L8iML02A7A9zZEc4GwpiH+M2DCx6Nq7Qzc0xfgiuI3FPZoNTmnhuDddew0PaFRU3k87R
JViCS/05iyLqnNh5HxwheQDQNUhQAmw80vM/IzYjP5rbngqmnkXMia0Fr5R0likoPwQUB1mFDg4c
jBjtn2c7lRjRLQwFZKAHKQzx6OLhxAXL5wGgkTrK3UGrX1amsWt5ECgMI65oVjZdW7Ez+LggdXB/
5aUCnSOICY3ruqlcioavgX9vA6M2s+PO7cPbNiOzSQFAUneiri2hQeZRuqFLQ8WK6R+TvidLLmwA
CPhIkYyLQid+SwmtowP1JsbucjVcx5R43qSPWLQGyQQIsOPhDraFjKBWRcHkoUF4i2tkKPdnnl/x
EJ5ulnSnv1hjQDWcYGTH1IacZfXAmbvIkk7Xtn1H0N64/ho4kXSs6YM/h+x7s0Pbh4rRvgktMugV
3jU5LE9P2ZtZpUZoF1iT6DgYsKirOeMpdwni63B+smbtH7O8STPm8WmuYNAd/kA4bEeIJl3Lsj80
j8zzM7w5c3m/XspZSS9BkoJUWSxf6Jq3e6z4cpzeEhUifrevuZQ7bTkfMZzd1GrPsQNEmaNTg9z7
Ar97o0hsmAAnmPjP0XhsyEj0wwnknaV3keGIQ7CGWsn3BXft66VrUiDvxJww/fm2vcAMJA7esmSc
DjBN7DOd5reThe9E+THjCE7Di2XymzC840M5xvoRAuyVQNrcnYrgqL+hEiRruO73fgyfQ4U1q8aw
+Mr1Y7Ne6TOA2E0fc8q05H9OLD21FdmDdC8gghGBxIx5UmVT+EErPwMOA7qpWEjwUvkBtwvF8i+E
V2Povex5uhKCjwzpAw6SdBT070UyzSWjrm2W6CJ4vqbYqJvmtBCf11alYJR6V3DsDUsHW+aI7JXi
Vi0Ga0UwIC1QVllw6xAmtUEQa77QoBN7kBpKhQGqWWn6YtUyYwq5yVwgqPE2/+haCitByhEruJml
6mPfYokFUkwFnDmB7HvRRo0UiQGGT9an8gXiBV/IOnfnQeTuwjFW5DyPYDSIZGZzWAh9bKx7VBs+
IKoByRFsv6RDu42Tuk1jFzvYCJKVwlB4xnmbNWNh11PQ/2KEPuq+WaPJ4OKUW9fewBoBlLHc20pt
MI/AbMtLTmQmtfNuilhcPzxMDgckhs8xXnmZaeIfFFza2oo8AjN8mxJwhG0ayy8j5BgKrmpwrzso
jLvAaB/p/Xl3CTG9uGliwQY4Qts6edqVDhz835Aa0zBOuIYnam14vk3y/BH2So3Tuj04ws4XBY4W
vxYIcI4ET2zq1xaYDnR6IXaZdxks8XEN9K7FvPYoYJq3OPNEuPNEGaMljKQw+7jYBkg4T11Ayuir
pFqxtQCh8af476SiyXumcBU5QRSrzaEKGKYq3p+JnoRgvH5LyrRQ80qS42WCNJvfAK+Qinukerg+
2WBmHx8wyCA+RsBnjq/HHDVQfRuZl4TFMr+gtHQ/7zX4Ig497cwrMg5o02OkMSN9Fabu+AxDKCrh
BgXUevcPfFnY+4QgHJ1dDSlp6/ziiY6k96pM4EfEBRhrKP6xy0iymKpCxxlDFCQ7iimO93G5sGXy
WdG0NBZnp7x1PKFAitbIuVYDhHGElB+qRi2hiVtrBnMj/SCsguipCCPunGprqLr8O12FjUyUUP/z
0MPIirUpGshLFMBF0XUUUH2CNOACvFgxpeVcs4Nr4K1/RU20xW16lSE93tYc49Rygzmvj+JsxkcC
LnnhXd36mr9AjNhWCoRWLQQZkVcS+H9NoucapeuBj9Ddg3RQIJFLBAah4g/NOSyZCtj2NJSU06Sj
debaWBgCGA53U4N4+Qk8GytoMhiZMkr5B/xvtL3lr0wB9llSvdGzadRHLm1/vBQ524A2S95ZiD3k
U+eOEtTTJnrHEmUwZ56SR8A2EoZ6UvOIWkNBNPMV0z2FBKLyb0jhYy1+KYsRXUMUiRuugTiuWe3/
i6BDFxfdyjjnj4FZfblbcyGjNpeU/wuMbF1eaHt06NEflj+mno0BK23eg0BXhYchys4P4vYYsTH3
884gGxzbkq3jJp1kxXT59+bdGUpCtfnCB8o0XqIVFG3ipkOv1gGtVIlWUQ937KduP25kNfZw16Rx
lfuwOJVI8wX+5vrZN0KuYMs0CE/XsNqfx054B+/0YVs3LDTy5sOu2PIT4bLehwkYAl+roKBhal84
lZO7zGAPKXKTbknfV7IMPgdC6A8xidpdCtfFQhL6iql275mSfYRru2GZRgwq+j/iuiRRAnTdt1ch
EDcaJ9lDdVZF55cNtgirNVzIPr90sZPLS9umvBP60gggKojJASjPvWZCcNvID18mMel+r4/TwUNQ
H8NTBe0pW4OL+V6IVFclC24LY7kN2jvoHElqYjZY3Gi7lPq+eOxcoanYZRJ115+yI7RfNY6heOTI
+aNhuMXqTeJFebIl0p7fs+HHH0ZBk7p0BLxgo8Zo61+D1TCkHVuBOB3AuafLHW2QZXne/4R/MSIg
EkrDSHRYAjFTY300YVrNTAUmTuk2gBDDtYCRDte4P3yPDl+FNwrOSmWs1NN9AqcNu015quYqVPqF
wd4SLx3KKry/koQlpLhrP4TdfVH4l3El5R27rGwuJ+bMLBEuLn407Xz8G4c9ZspeAmdF/vUFeSdI
2bl9pYaWYfOLCVYiXB4fmLnRmB0xhxgr/zxHQTutzs85IeKzUuDauhwxGgjULDygjs77+05R2b9F
DNGElUcb/rjawEGWVsJ0GD0j/SZXnwPcH3W42kVFzYwxNlt282Oet0//zwQxysdiIZAF7DPT8WnA
pe4Uj1VmXUmRbvyb6OT7DJGsXUZZveqoeJFtnfg8XdR9gAhTGKYbstplZeHKd5WYsXIVGnjRCqPR
/+QUoN48smrUbhPg/9wum3sDkA1pkziSbdadI7f8vXO9kGaBLIKehj7g6vSBIAeTg+tUTBp6+MKT
Q6uWAL/102X0ED9fg9cw77qH+9UYEm8dhtV7bttyhd+fjgElHKbY0b0wDd6G4UhBDZOKdKnjD2JK
wfKtbF33EszQHKaKd8ZFvPUxiZlUoOQCX9CF12w88bTyEdltgMEgj8wAAPe7kaHZABiMzSMCuM2q
Ugk6S8MqtrxYasTPIPPQQH62q5DqHnw0GQb5iXcPegnyJsOSBNBBceyk9+47O/tiHY519aaBM4Pt
rVsSF0sTkxHyFf9JdnrgnFPuC5ruzDYR+HSmSr8m6ivtLqQw/B0S+FSnOzcCjyMnfqKLS2V7yZ3J
AZpBYsJC0PO34B+0ciFUnFPveIiadCth/B1WsGfIgsfH9GfHrMiwTLrdpNRTIDOzY47DS4VqADeN
O1lQLJgSitFrGczJ6bgLevGj+e3ofzyUvGKHm5hdUdUBGYMnZp9kj2CSbcf/d3TiBHdi+/il+YUN
omrYjTiguaNBRVM1jD+bTpOMZxK/zQcTgCw8BgjIxNDNAE4VgryN6pIwhCEaVE59K9Xfz6Pp6JNs
VHr7JL7owtmTPWVJDvpY+UHB+ndZ2s8qkprFsyIyPDGGGz6WU2V06Jv9ulVtixc+Fw8dXu2tgzOx
UY6w89iM8UzBnhyxsIQKH1auyrWX/6UpcgyjVcIc/11mNxLzkfsphjZBqqObac3fWOUZjXoflRPF
By+cqgxeS9HECIg3NenvtCksI48Fsf8837cvvAHtO94gBF86Sj4eGGkfxMjmZbk0sinox3uZae0m
YGM3nBI6GTT6i5oaFDxR5xvoUcizl7NM9MOzIl4UfAflDXsHWXpqf48arKJnCJoR/Q6lK1TVLHZb
AQcmrA0ICVFgiOlzdEPV0w5tkTvhMUO+/iig6iyhmGunNMiAK3SVvNDKDqZeKe1Y5dmH0CL6ydfE
SDsdHJMUT5NE1QvW0FMCLLUrtahRjOrqh9UlLWVsH9CfNVi04MTY1EyNo2YbGlxLO64/wg6w4Vh7
hOw0880u/z8NRkol/b8s2bSPvJO7qxBggxSOibV7hqGABOKHUIcGApDPegkBiuuYj7uRuNjDuaP9
rwmjbAVGcxJQ8dhhj485xj1ZT4fqUO4aqJL/YaaUzNa7Cd+x53IlUDnfpL9DiDsbqnKH3rjSNXpY
JSZLTVcuIv4LRjVqIIBTmVKVzZiIG1u+Btoxwy2ptzyd0zrMrLmWRwhXr2d2m0y9qYyfU/PJ9xg9
PvcFNGWtcwP6pLrqDbb0YqqEZ5gA47VgS3lPweigcyQUMRIe01H9SzWgveO4MZtq9PsTwX3To4ZQ
iS3juzOkmmxJz87GhBCGCNP8h7Exe3/Sb0Krd5TkbOFvF9Pny6C5U+bcif/vbymu7KVxYy1jKUSv
4loRo68K6mkQWsEhglNKHUlc+MET7hOf+x4er1Te/p2EsOpUfPL8Cvb0ZwCCdfgwYdKTUV6D84mh
wk/ysA4a+akULsMVlQeDhY7uh9aiIXP8SqjOEMEU2QpFk2cGt9E309kIwDNqiLPYAnHVDGpfNnV7
EC9qak6HIlasZ8mkTgL5HS72vGf4Sv4+ddPqrLBSMl11SFDBH8mP7cB/5+WDjNmaYrPSVJa2NSpi
Q+JWg9b0BYlh0Fz8BajwmkYVbFLBNfktpgMAGxwYMklUZxfcTMa0W4VeegFIL1rErc/P194JefLF
uNkBPBuURg0uwgve9r6WqupXJiIYOLxD/LHsTc7Lo+uHpPyAS8zzuDwPUzKeA/FKwXGXD5dPrn7a
Ngp7n85R+v0XaHDWHnSit/ZkoanfqfgesJXugQhnvoqMvJVgwb6RfRMSn9+yLZDsdjFrwPYQlb+h
HjLWgcMKSguX6SbhgpHBYnIG6tnWeoqjX2hQwTq3JLtqP4UQFWLa+pYcakAe2kIVK7tEHcnEtePu
BXjz3kMtIe39Oh7HxMvzgkKJ0Byv5WzUKg6eWsEfs3vYmFdeVfPstrxDXnnTZYEAJo4sTwElAEvB
02S/hR71ntu9pVjw+joBjMAO5yItczIicEfjLzepdhus+8qOugwabTzCN7/iZpQ/ABZHdA3DPBsE
UkhVhdG1DwWl8PR5On7PVNGr3B080IcbX+BWbZM8wf2ecdfSxhoTx8WoxdqSwZxqP6HFN3rv28hB
tcv/DO1hsM7zpaqTQglFM9MlDT57iR9vnNAHutV44atNZqiF4qyw2m0FnlzyVyhUBANha7AdaFs5
NS7lzSNxS/egJl8SGARUGGILIt1e0NbxzVYQMDiSEoqJGRrlwg925ONP/ojpYNyl6mbr1OoDdOJN
SNWVZQAWsdszIOozRlifS5Nnec/vPxCqK+PMjoXb7uonGzFUxTfLb93GnMsA6DJrCJ/wrO6nPbL6
mzEF4WFlQO9cABAU18VJMDHU6JwYqGLrDbQAlY5N73cUKpxBy4ioQBt/yyRgJM8QHXMBdPoG62uH
qW7sP5i5mHF0d0W2ctJSX3EogdmwkXkGffiiuK1xbI0L7/5UY45u+qt7PG62Nh7exGtJeyFSpOxz
rWUP24P5T7sqX1QVR5XYuC/6nd8UfSprM/egYigxeC3Uno8OyL+0MGceAo3nA28m6bQ1Z7qfXL/X
FFGKTiNd/3zZVdZzwqY9wt/rS/RCEMe3YlLrEzK8MRCo4MEiIWB+B+ALrvNa6kMcLyHJNrJYSWiu
2SwB8C6R47/4LQ+Yz1H7KzfIEcFPjpcSzD2iBNknBJRhYBSgcNr/yUhinCNw/Mh379zs16yTVmci
o2+JSqcOkmoxHg1CDVNOAvIaunFePTaNnSkNqTXeELiTg7ap9lQRMS8A9Ggs2S8TT5o3+HkKs6sE
Keg0hEBfwfJ/D85YbVkXrfxkI0cbxC5B1GEvyFU/8IAnM4gax0n7RpH1k+T9kPrBm231SQ2MOvsH
bNNedOfhmjtEKWMCtZOv4n40CaDpUKKL7ymarqWgYEKayIc35/5Fva8YLB5ts3k//Bb1Wi1xR2Mh
tp/Gkdz8TH9zjdzaDayRErWdWzFDDH9gBGoRWvwXMP8UwNrXQBgBEPrnzuNngNE6Wzgo7Dsvt/ua
Dy6Ay5Vh1tc5vrt556r56OlMzRlar238aisxbYDR6/DqcNfGcEG88DrbE5ZLJ77ffVIbjtUhPs+U
EygUGp2lrA4TA4fePbcnxsN45mQleWjnqCHSXrjy+YUQ8IVcvO/Qj/FJNfFBP9y64VGnhpANQdJu
tNoKTplSk4O31+ZNMhaLrqrz8zPefAnZ8caA7OgUrSYSw8j1i+wBhF3Dxqe/S9QgC9Say/Av4Sd6
+Z4AFZne6HQwd6UfIpRP9fJFv0ldZkN/gepNMtnsWDvJ7kMFjdfjKDJmWmIsu4wju4Fc1zvMWftu
XAEkmqLBQsIrtQGCoePiNQM0mZJ54dOimC5V22ZHaoQ3NNDYh9yshoyBw4g9yIEyOkX/N2dPlyNd
/Bu77XaJuEToIHWzxAYGgZY7l5DA7AtbNCUjGywr3xGLMvCiYuQ/Y9aGgCGJWCNZKnLw58sXrxYX
jg7Gr/e3/dOifZ45XbY9zursbPiqNm3h+aydke8fdvXqx4V3OdpvscK+ylUjHrDSP0xMRUWBZCsW
Vw4BQ5vNqOIHM+e6CQDeLO0yGWz8Kp36HJRnn92/dyazf0FdGZAxKG7o+lkDjIYygCH+WSmlJ/Fr
o+X6aNLeWwnLMu4IH/XNdh2xbz0AewWUYzVrPlIngLBty+ly+YeAt0V6KAh0vTKB+lqEzxe+NH7Q
Ef+S/shKuqqASpcGO8dkWrLNXSZSqNsF0IV1ggF3I0PPLblcotOoAcYswKIftFiEli7H0YlVLqkq
qjHIlWMkKrjBeQOu3hGKuBiJvzSSXPsvXjNkoIqFdWcUW6p/qqZlgl0x2/r7cDNYV1UrO2qINCUL
fDC1aBewJpcs5Ptis4jZLPdzQ4ACyhhPTS3DU1R8CIQ5DeJFD6le5TddXRD5k0uvxywnlaOeLIxE
U2/fgwFE2ErM2riDGNNluZmkx4IjDkN8SpB6loX3YsQuJj+nLDkl/RN6aI9SOGH6GqgakG8nYFt9
fN3QO5A+xN/GDaVB5KLI6AcSFsvQzRmBDPq0Fnrwvwu8tk72HZqTxA3gCxzrjs9+6wUkgIr6iPMF
tX+oJxEW7Oe3/WmmU0GOKV3ZPUKZNb7XaRvqPZPa15HUfjG/SdMP66ciHmWcKFjX8c+PaqnziZVc
qcSohr5QzdEez/jb608gprnerUGN7MfFqnfPmc/lpiyQWmexkWl6ZfUHqkQOpJS6emzD2WXp/jq0
f8u5UZh+7C/Snsra4o3aPdgoUw3gw9IocFKPpBKQ9QRUH0Ixd67MZItqIJOmcUie7C9/n1dSac3i
vuJb7QGHYWkIEuX6FX0F9ujTdWW6OWoZz7q85RO82UcFTSN9jITkrfE8lgWM3JodDjLdVU+0dwgm
3rcjdIO3Pkai8omM
`pragma protect end_protected
