// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jY078fRyEt0LXjTkNmbx0zGNx9g3xkaCevyTlZQWG1HUStPB9f5crXjc1ycI
ycFleje2I+oa35y9e9DksMmmcLvlmnOoEFLX8ol6Mp81G0NuNj60iP+W+kST
nd2HImoWq1P8p4kcOyDwDe67hWkuJZzVY+KA9BCHxBV25+aCN393hnCZ2HiK
5B+prN4RhOoaQZtcLNDTLxEB6t8jqXOtmxAFqcJNQYzt8UgchTgUbMcmH93x
oViNdce2PX/9FFuchwVu16TWISXyysQktdEXPLcbZTyP9jf+1VPr9n+Ch10u
MSoFnG1dy3IpN4RIcIK8mRahxfpwoAj/TvHn36LD3Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YTreeeJ/osqphxW4OuxIWu0q4A2XFFcJ7Vka6hff4BWXRi+hITBY2E0ucNWn
OKGIwiq3fCg3Juf/z27RwZmfMddmOWs0LvgDMb+3jVDDEx3unMmN35qNWkmO
N6QoZDh60hERYCnA9CvqIa+Pw4ZTo2ZRuRUMIJdaD2kLyWPHGCtJz0vUblf/
iShJRnkOTv+ANu0rDiGlL9g7rtV/w9SxyEXEbpwIgRmvOpVWLFxHbdxI3clp
QbkHWd6K26MzK46PD/QasZum3+11x0YJAVxBzsZhvXPAl5ECvaMxYT4TOVEI
7NZ5AvIAvvQaojX8rmqrLanw9gt2w4XAGsd2wLaeeg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NxcF2CgNomZ8eBsGVs26Vf/UIVmfvR7bgrSNPHpa41oS/8zJFdE/VxUd4iCR
H+SZBsdB4T+LIK85SiLKJReaMAsc4TQbf5IggD0t9N0j6wCLr0ijjkAxtO07
yljnGGHsnVNvFpz8lVKPHHxzJqgpTkuMevXmV945G5TgDCq3YqeOKkGmVAeI
N4Jl80akfHK9nGFVm7efNbygoBHzvfvTv/ZVraaRIGwO/h/EnQ3lpLsIPEu1
49gV8ehXI6pju6+VxciZ9Seyn9OZC+9MYNPJQi/8hRK5518nGVDPEm3zkTUo
6esGV3S6NCT1YLHuqs2+8jQDusgqowJ5AiiQwJkgjw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rFE7l35UoYtnSZ3dPsdzLc/TnnbHhD9+eJEujWTML8YoY0Y6p1iKXMrXQ99+
6nyvZFPYcLGSOsmYlj25PErVuA4AFDcOXSXMg67xgUiMyeN7N/5CfK84WRYD
UoCHTPB9wPewJBpR8TCOm1ojGrDi0SfTyXQ/cWzKENiuza/OMsQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nVVOPZsDGHZ2X9lEoS24K+szwPGrXy5fsT5dKuOpESctH4SA7iva9otcMkye
2BHEYdt+Qs9CwH6QetbDzwsTp8AcBq8xIMpQDRMwg4mmuhsE5MBRxpA2yrDx
qkahVNr8kC4cSwLUQRb23VFvZ5O1ds9Rvejk8BfA+62XUwUKH/d1HLegVcuz
aDWS8O+YmnA6Pa6kJQKZIUO+jyZ1YkcS5oKdOtwjZRTFyTpC+74MDI/IamVD
bnHEYAT6crAPnMZYuegEu35l3DBe5BO2+ZsGpK5NoGQlGRroTQXl03V8hHup
5lLFghgY/VrnX7Cu/iOv5Lc1qDVDpkcfjUSPKRVaavm0CAbnqnAticN94dK8
h4+a6yHtbgt8QMMdInjjXiULD9dIgvCx9lLWfcTXPCJ14IvxTPOXFragi8jp
81M2n6oyQF0oI5045rs6SW/IygcgduRokFsKGd8pBzE/8DTFHEHNrM+cDKmp
+XD2+yd+7p55py4qFIX7Bib3GlQUNpiB


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uxs/qREajiSBVU6XAd3JxSe4uKKrd51fbXQuGPRAnJq8ROF5hky6LoG9HfKQ
bFdfZeIHcFMcd1va4JEec1dBNHOeQi4M4O7sbormQ7KBLBkjt5E+Hqn2N7zU
LTlQFoWItqVN7Dr04EOHwBZ3WypCuWcqPzwBarX12/23/TVMBNE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MRJgX2K3RqlqG4DL7rPdpZdhsQaCZZBQlVLGSC+h3sxfs4p6o19JMeLVyE6k
W74EWPdCrw/6ZhR2XExO1xY8dNobraiVmx3gQYxCjtQ9o+hnKI0siPjj1wdT
1gqB1leVE3tK0ag/Xk6Eq7XgoPTVJ1QtdBM6Ilb1/6MjYmHp3Ag=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8304)
`pragma protect data_block
J6xnZRjC+rtjw2MRtSllRcxg/npLwlMowSKqB1QK4LAm1QFlXOhRHxP8OCRC
NFB4Bb0eIhQX1ppr9LOFe10ylQc7l1h3cOHwSwnvJqA/Z4oKWT30+mKLtIxt
8so3+tEEH8lBFNkY8lYlIz9GDLiVy/cQqRu41qeJlsIEj2LJGRFgsPBAl6m4
UzCLB3bW5CJkCYHT4loz29c8vIqOZ3NUAixJky+JNpLRfaPo1pD15Er0uZLS
niKjYQcqN1q6tvMhJ1hk8QviJTyOGEg46ho7kcWtXGvtvmYWJIOV4wskLch2
idqM0FKlx6VGP8kOovzCZRL/Azs3ZJFc51jwWAL/tZHauvfXZHOUa35J+yYn
sJvVwG3cHv26tQ4xxMsI7Yk9Yund63MaIulkxRpr14R/Je1wXyxCjMjIvMC6
MY3hHS2SO+LZYwUPXoGNYyT95yiwC8iZ5NmxHTP8PBGGN8l6KqmSgBOa/EfN
v66TsPluDp7DtJOEIkq7UhEuX2lg2CU/UwYjsrR3qWWzQhn30l3o5nt5FW7i
uhYlEmiVsfyNCjwHMeRG1ONi8EBlxodPwKmBYT4yAGDhIE1NmyWfy/e4vkTX
+G+zMy5xNaGVv7kWfjd477U2HCCPnIgUWjKmmtcWOeYCm1BlhEFmk+SKlL3C
bmFO6PPucIBpovwre6lA3g5u4lFE/kbBFzbl5HTMZHgUfApGXAHNG4OxfzVE
C3Z4+MkSctbcaMQI0PIHFWxQFnh/6glub15t2tpP3qV1OZFbTibxnjGr8N4h
3ErsF3/Y8w6MHHKyKIlEMvaFVzIaJwhZbFDVSg/vGNh3slvT7cFr6JwifGaY
++b8EOFz/o4p8Ww4QW9U8/6n9OSd4KEwJnoScPAdIt/NsvzwCqOJ1KtE23+1
NSrFTXCxXnhF6uUGJNruqhXsKfGYhbE2ncavLEbSz/7p92dYPcUgHKwD6MoO
U/pVi6Gn8RY4MRqCm80pXzwwXPvXxQ3L4uCnF3EppAdpbEqLzQ1gA4waZiey
2x/KAxbRXKWSOflYhV81rhxOefD0NMvlvjRiIzpLMuhmqz4+EulD9XJfrlAS
jlqSoqIg0gmfJ2ldm8vSGSiesutUf7q1L7AxaDBpmQ85JjEpKFSg3U9ag0jR
Ae9Nvqk7YdnEE70PYvkBfkI0KsqIbqOjYTlRfDYqCmuySMNDFOSKUozfY2Cg
8ZozSMNwqu6krwpUkqoYA8Yv73p5O0T/GzUHHb3kmRvwGWl5h/yRvnPfa6wE
FswXirjrdQdLIi2RAAsPyF/RQ8LPh6ESy3wezXFqQwKhu874Q/1low7PuF3f
bGixwLZ9rQwGxtchJKpw7MJ1G4LV9lX7b3BPJ4OuJ92MuHOtsLiKqnB8qtG7
Wa9Nch1+7etZ5mgio8+bZ5RHZwnPrUse4Xl8UChdBMyKO8TdC15Hmo0Obisx
15RoPS6XGewuJpz28DzMFLm8D8I56nad1W6MyvTTC87+2Fq0lpZm3VdH2s/N
supvt3j8EF/2IfdupQ6M7V6m/BsUToDPl573/KwYd4GB1rRFBalnhOeNthun
3q2Zhw5XIn4ut36JkmbqjD7AeGQuvpXTcoascCdsVkV2i4SrZwVJdF3PFhWX
/pXJ9FTlG7ul4ffJXgcsRjJ99mvyis4nbg2JCU5CRaSVpXJaqPWvG9DX1LXm
ErAif4u+mBkVGqQ0iYlY8syu63sT1zDB7ALJ/Pn06c0JJDNpuY+S1q0ZLDyX
HZvT4nT0uRthOrMLDUcoRnDoAyCy+5nUDdt6SKxtMj8YteErUu2pCj9tBCKu
5lGuMPV1c1rzI0ZCFwOdR68BYNFE9iEPuQRDm80xcFfs5OGuNcynGb5Yi/6u
1CEeDIrWqJ7gWwxbY4J8uHjq21bCZajBkMkXvNYQP3yl6KX/3+OHEIb9VNHN
3TIZDrPzV81ry24TQVQWZGK3ENCC9ulWKvrKz+7CSOav31P0YXG1XpwaiDwM
SjPzC4AvNdZVTmC4wGtgaQtytiMdEK8/KJR+Rfj2DmAUzAgVig3md0CIr8bZ
WcmtE7x/jYtukpyrB9CMMYvGNPdk85Y2n/9CwUAKAppODX1ze4+DxKJgqtAY
iwwPkqSM3vxsX7GkgY2ImeB/nbnqTXAMsebaonhv/swv16CqYL4zQ9dYGZen
CbI6wg+LtYynbGz5cRocSj4aq2VEbRDJ1v6QDgfkhfzZykX0XlvYP+W1WoHd
pqFvcsKM+2jX+BLplcRh0lCwbDRGGktKkguHyh0cFTfti7Z2BpoYnHeidrYO
ShX+KMjAfrm6ew+4r0V9FrUB+xF7HZG2cHxfv/bY4WMi9OnavA3ndBqfF4Rp
ykAerdsu0lizxaqXlqssyzsSMvCYuXzWPa6EhX2c294X3T6do/OC80JwSP7I
5lej+gOGHAbuX9iFbh2S2CFrVF32szriGWI9sWeLX1BXJGkIrwiOTCkevLhJ
x7NrFCBzeWERC1X1CwJVAJfeR3OON0sL3SLp69TjfFeoO795LD1dIzPn8j/G
ZTJtTMjDVJahjlRqWQK8sHYbJNitH2ZZAPnnFSV0JrWw42VwOFfhaQgVwRdT
niLgx5luiQJgJsqntXOs9UwzooRzQHVTcCF/Fa303wU9h3+KhFi9X9qOKhkV
nkxVMFDoeXhPX5Mx/MP8gTU8KpOO+dnHH9CGLweZ9liEImqQnLMEqs97vm6V
nbnHZqS5lVtV55edLumrQp1uudTWHxJca0WjbNzlyq5nlpTllM6Idki6N7pk
WR0W1hfKUxJ93UFzALodwypAqN50njPJ5FvAIX141As3TI7J4PhGxOos+HOX
t4AMk5yjuxU0BbKWfaCKEi1e6/VitMj2nTBs8/h+LLmzQlEH9rnxR76VxuWe
EOx6uMWvSA9qZTrxiUWZ5KE7ROXvJTSpEO4B0m2YY7Vgj7dqV16DN2r3nHus
Bic+skBnJTm5tMB3a9+iJOMvZ+zWjG2XCLeE8EW+yIx34iH0swEKhZspYJ9g
6si9h7qWPbBDQMgeZeAE0JejnpHkjFFH9Gj122x4CaKi8oQCoLYvFlcdyAtN
6FapUrptgNja1OisHUTeSwW7y78wtdI/rw1LaZeWBSMir3HvS0BGDvhbORu4
s3ivDH1q6rlOw0ftBaShwB77+nOG3V1K7Ph0bOuLFUlgWHYj34hSDgqINw+L
gi3fgQ2b2utkKFkp4agkluhE4z59lxioNwFzV08Yo0R+ET50s/Q8dSALvYKD
dzBWOBgFlFautkELQu61nmRbNQXh6o+/BQVvEQlw/ZH0z9P+Y4EoMX22ZC71
qzMDKg589OxVYg0LbvsKerLbDLRjfG05o+YPNyW0DKV/a+l3u3ji61YI8atg
gIE+AHANFCgFeMKs85OR0PZFUlEllkEOm3k6bkV10DcZ4NON3Z7LacVAq3FE
GpmNyB/0yiTQaXL2j4eZKlwBQDlH9XvVEB2A7ySjpfNwIop2LH9qMNRFfwAC
JtKzJbyHpsfb6g4l+gNV/Gp9rpubWG+GGiWpq2PpX73mFCZTF+13je7w5ZaH
ot2xjvfaAfSjQdxjqkyQeP7RzqwyPrAuDa/QQkLV5SbEQSz4p1p4arWbFhxt
CFALVDDlP2WBzjcW/XpHBqKn9mGzFVjzUeyR4QwG48prGRg5i7xNcdjbu618
CWOu1OluCDdjovvNOXWwNaonqxvIihNMfzEhjKHfWD1+OhwnqbwTiu7SyCnz
cICbZkRXri5EaFYfUkeyQ88jfxy4fmHWksrP0Jik+Zp29BEi5XShOP0EGPdB
Jk5pjyBPdzUiR8fdSsiLVP38RUyCrkeTEeO/Qv0dDFQkjIvdlW/y1ody5Qcy
mKkDu3IEezMPUAE7GvasM2xeabLRdq3gZWHnyBDnQk1O4ZBh6bGgG4LtYLOs
jDLYiCNF+CVNSDoHFnB/Y3zFR0eA+pz6eE1+kiuCxU5ZJOlOCxfftUCUStOO
llFl8MW/JitLIWdbgeQji13iZK/PIw+mIz9/uH/QJj6Yxgpfw9xSiWfHiaQu
L+qXpPMeh5JeS7oF6Br/mEJXJuAbJcXNGCw6xKjBiuSpxb+73zthmX0K4Al4
cwuy4GGMoUbXGAgcEkXFwsUit3HnVIRJt+IBFBGXPBLp9yYSOJ17muEyoku+
4L9hOy5/1EpCbshg7T/mmMd8MRX4x9OvPczbf2M+6J+lZvGcZNlbhzqNqdO1
UwowXFAd7ZzdlQiiO5A33NN17B7ZuoiPkj0UMzIuIOo76z5w7B8Leac1zNTC
Ge/ufpRZqWLrokX0o3opF29EyOk+v0mjGCWpe4k1Xvwf9GpB84p8ZHou/xel
LHlEAW/azOGtljIklJBJ2B1uWcVhOwxIXbqQxgVJk/isGmJKO8a5Up1cBJOQ
adUJQ10Bji5urN1RlUJjhxPp2X4UG8zCzymhFxM+y+dJDrTyitjcgwbkChoN
/LIGiHqme2H3xpl9UckeYDdqfpcomnakY3IEbGuShcH7+6hz7JrtSRHaC2SP
SmyowLbpgh+xH//PBM4ex3TtSmyvBLye1hrKr9jedL1HevtIWB/9CBQHAXTv
9ax+/aD4b2NqM66wCo3waCQBmrUU8NHqj0KquBlIcRWs29yc1HTRBdiO0Xsa
0Cw7C76+0vAe2+6p+FDdN/gD0aTPyFcDB0QJhuekRu5ofqualgCCrcl6gDQj
rbs+YZePzemVDnTnP280lunmJWI8LdU9tH+mT01sNO+4tz0PQSpnmaq1V0V3
sdSjPXcOW1wdgJX9Tm7euyP/7jp2pfIoRQuK38CLfsWJT+J4m7tdtjaqaTJr
AVd3+JXp9Y1RxZEAH14Ldy0LueW2DENBrNiKQH4axoDB+qE4atnUkp5tfTAB
5r41m0hCKRqlbHTlzfbWu4ZPbzQJHucUKsmn1qgQDBUwBtvnOWd0/gIOW//n
NYaItd8Zwq9Pm5YhdJG+WU8j2ZUC+c/11KY04QDFtT0nBiHwFvIWGYW70BHf
VqL4TnDd31nDtIwAdWUiRbhJOJRo8bgaTpPr/GKS/MkkwcB4VnH44pZItxzu
OhuKJ/YHvqri90tAkJftXph7/BaV0rhDsTCkrvmaLRxb454lDrc/86EclIjt
k6Z6IuNmVtg7jbigtWL5nPfr/lhYbuBD0jhjHIbU/3b7l2o7nqFQ3VnIuMRf
nDYnd54811xPAcx0WR3SSoiZ4HSQBgVwloNAh6fNDsr6qw2aZABNH4rr4m5m
L6BR7mjwgD265IuqWU6iUrOUNAX6BM88E4fCrv0QIkXzDiMPSg6Gppos1Evj
CGQfYLup7hpRONGVQLRpnONna9OKZa/sq9gldcuaCQLD5sYcAZXw0gUx60Jt
TTgY+ulmkmXaMSZGI9lRbc7NHe0hJ4azDAyq3GbVKBCEZuRyEyZPcuCxQeW+
xcT87FflKCguhW3acD74q2c0NiXVR5YlcY4OQXKgAJzS/UtvQJSZu8vihcIG
qZyfHojuMl34TW/Oh/ipFWiBeiNDdYUD11eQ0pcz3tjsfUnKiRcf+1VoI2mP
sbGA+BWRFxQMVTQxsu+wK2bBQuTunjVKHvEpFiQIoW7s6YeC7IPG5wvQFW2M
+90FQ8nUbbx7DFPlWvMlskUKaa79H0uEkA5z5MafxQJ9bB2ZM9uOBXkd9Bao
o5CYc+nf2YSADlF8qUVlzg4Rf1eaVd301pgsQNzu8lWehNJxQ28ryqxztq3n
sTFTOIjUG/q4Cnwutp+lXbUep+6bKRlLBDDnHUrbJZEgkoYg7QemeYR18iKK
29iYvKQe+EdkwkdGc96+QqP3j8JBJYOpCJ7hc/bYN2VElHoo6ATBWIkGyceU
8YZPEZ8SqAkoeausmGgTEQzugzpQQXyEA2p0OK5lB+JD6GWkdwYcExPqXvvD
AL1u3oBO5COyoLg+ZjHQMgb3UqLGLaz6MAhbH5ccXBrdWGbtH3/dwNBGMSWn
VUP36CFlL92VapD7HDRSCr43YJ1BOnCFxLuVusP/54nR8uKKQTiJkUoe4DZH
46iu2LcRVPRjzD/Dj8BFgmpAU+kyAVG+MQP7kxjH5Dzju67YOspm9e1qz25+
6x5oZFy0JF07+qFAZkEAyj3MQfwGFbq7fq735F5EkQn04JHHTKQzlCL/HQ+r
Wlr/QeIs0Xm5ccNYpUQScEc3z9zQTUrCdUKNuTHq7krgO4QpiukAQ0hky340
yHqRGgkW97hwz7yXgl9kVUmaQSwmi30/LhW7EmuhTI+04WjHwWjepp4OEPi0
q2mhe+8zCRKRyKbjNuPCWdkjTMsIo51IiaqA8GYWjXPyrEB0abvDtNavZUK7
jCXbHKACdu2UKOjqZ0kjpzP7FVIMvOk3E2LhOMhhXMOEcFTRULylVuxs8IuX
sz00pudyuxug6SzlhCct5mfwXnN9xn+QWUMKFtxfVwzoWcErSl3pr6Xu3lGz
HlVDdBIsmbpUlo9wVU+x2eRTggOzlNx715Z76VSk0d8Okemvy66XiXFuoHqm
dGlg0MX5ogvlaV49Qh+Jpv7RgGPVbGEPTGDH1Rrll4Mge8BQNek5cEZM0IFL
mgbhtcg/YF/fFTnE1/Xrlz2eX2+GZQgRbQITRgt2uw+nXFSUswTEMoRQ5uDv
JEeNcsqYIuquKmr893hS385NgJC+4iPQ85JQNm6cyhppyTZZTPYGzTLe1S6w
JrNd3LFSOZkXmKsxl63AVXCVm4915Yzt4OyqIOJr73z08+TDD2eblqFZwc0s
ufq1w1+CvTalPErQjvP8/5YwOmodICajaBzs2W8zbwztYgSece/0CEreQPPk
DeUemIvdG0wJfqGXQRJ5nLBGVOyJ++cKPak5WoADpQLZaL54YROBSLYG+I3e
BA4k6QZtnos/ENjhY0OGRSUX7nsgJrtVh1uVpghwQCtOM1pWQjWz+Ltdn8hm
ro64pU01xna7EwkvRlsI3QS3xC7uqMC+rVV5tIlIf8BhcF8bim619qt3NC0Q
1pNnm/nCMsmyLYFepuub3EfOnyy/NBqNVkGLenWlofH/+XcG1m7JfbZjc9Nq
4DEe1E9dLJgoFKaVyDGShlyBZoU+tmWdLVQ+NhSd9smGcDK80Xr/yQB3jeEQ
m8OsmHlZTynyU5DHzb9v/KAvR4PuXbAUTwmdQ4QX0CNaAyC2BCduvgWVALYv
+fY1uzYkWwhN+D1SpM+E2i8Mw0GmU2KJ2wVXDDdKBZN3RzL7swdICPwg7Qp+
ETN4WXnIy12g5j4j4mJy7qF2eGX16pl4iHBQJXk+jkEK/r7ODe2wvE+Yb9xo
I1bs8sZ9xbAVMBFN1hNhARNrFJIdtZigqHQtfmFFrAxW/LcTbRBzuWigx293
EDHfX/8gDqorjjB9Ic5LHdbwMIHamR2CJlM/2qSqdcX8SIOctNb62oxDMQKE
Q70F2rmR5g9/nb6cFzBa1gkhgZXqrbS2b9LqSTrQZKEXdKEpNytnPpMvK3xX
3r27NdXUq6ukQJQKTs5wmZQOV4Tk8DlGITv/5y61IWlDfKQWhPpNezpMqEau
jx3PvzmQhtFmP9/0/gCPL7RTMw77ePurFwcAdyQ3KP3gfe96p74LFrCu/rk/
a8LKAqtB6ev4K3XN0QrzDQqBJoVdl1FGZzHVUjvHMTHkF17JbRZhkoOUyHHO
cLUyLh/9/63MehHoLBDELW4OSIQXDJa7gEmEaYt9/4JgfcYxXx/4+V/VDDht
qCKwUdSoHshTmLcfmc7jt8SXiY8q7RmHi+pLQRqLh9YLSLQc/AISHfA/tJyC
0ADe/I1UUga6aVOeXCeA+95IkOtDpbC/gyJ7mavPPf41cRvTgekZCi038NPB
M6VudMXJmInfXyTgLyQFSaXF3kP6wXzVYnNy9/9ZQJbo5zon1V4Fp/IKq3uB
SQsktQ5Sqysb7PG6Ui6KdcmnZYI9nxfCb6/Htp132TaW4i8QqNcwTf0lMvGd
EluEtQ1CSSGnfE6cyrFcp0nx67Vpexi7QLvDhl9yj/IZvZE471vIFmuyxNC9
14h9GQPJLNF7wYGGlLrN+AUDF7oADE8A1I29/IY1mTS1f1J47YaNV/r7Lb4L
26Ci+X/Neo+tS4MLXAkVfU1xqXjp/DqfQLkG/nQ+yWMxkYFhIoDK1VgO2Mny
9OMIH2xXlZJqpaXNW4Rvm5/Ubixr7hNsGJuugWLCQaIiatN1wOS3iIo7sVor
A49DhG/ssZd5Se/xIYlOs2PaOpclkkmcQLBTUJ2W3h4Oiyemc3WjJ1m9qnA1
mRSgfH3am4G1vAjtkZ3OmNFVJI5HS5a6YHcrzSxDU2DUGHhaFu8h/Rgspb+y
WkzlYrTq/F7oskVWI/fSfXp6a3EZL4Xf40rLjX6HAFuVCbRhItplrZGCWJbe
wADndKWG6SaZxz03aAKoSX3s6qHsLf0sqaJn/TRXJTTUTz0+nIGSNohJiJMR
XKzuf2eNhBNoTH5M75KT/1qZZV/ck4/zlK4TTkTyVEiVHpBqoq0v88WBeY1P
u/7PcYpuSEff2asHwCzwqo/NfbkS+ca3Qojizq/dbAEKPNXbDehCdyv3MvE0
NNJC1cIkacEWuWKWBqFPWORRUU7jrrEqNibfPh4JgH+oLO8qNiMfBfJP4K3c
y6wkxbDOofEK5Wd66mue8/hHxocU9c5W4CDxaWaj3jaGqEXpnMLhIGGv9kIj
+SqLFDA6HBx/Iyymtv6CjbdRN2vePIJDo4EwTh0Kx6GiMuA1Vt5ULN/Uo6SO
QejMDhFh+gvlvx0OoPTVyXztyw6/WVHrfeab1E2yApzxWwi2FQUrgDN98Skl
0peXDUJNPQIq1IJ8WyURMy1edOmSCjhgxGixK9a57Pz2/wYth8tnK0o7z167
ZgxVibJJr4jUHDidSeacx1rxdqgv7Px9JUhGMRzYKWTbKOkdTwwoK1ZKA2Q5
/s5qoDLIu+qmUMSE2kWNO2Bq/pi0z/VYuvHZh7KCbUwDMnd1Zc1+QjHSFo3k
ZTJkvtzoOyIqdRMx0XjEFosqk5qgg1Bh9GzAOxVza4c6QA2L3KLhRtZmN+aG
6MvEyP7B34KP2bIlH4GLbwXS2X1nGbTAY2tojJwA/eo7zj3vQJU1Eq0qTpRg
kozuRfnLf9768puNaagXezzpf9RAyvkgpdol0xjTtns8jF4owQwfhw9j+n6F
hKrfIg78VAndvY/Jxn/OeOQ5FH/Z4aDdxxZJKp0RURzAHc5tLcXKXkp8X9M2
+bqyyrTjVb/uFHZIwtI84CkxUAUVQ2FpiitqukgoliADjXHUe/olZXMDumoK
Vpzia0hoXQNPhAzHXpYkOY/Ro8wT/X+eK/IyJJ2NKxRlT8KzheDR/OSkJd6G
Ozv9Ch4I9tqq3QrcMcImL1S/0jRpmBAdtIpNu8AeS5WMDR+c6Z/m1b7+VECY
47Thp/pTacQMIekMpeK3jk9K+At8JUDiclHFLTl3+Pk9hhfuRwLDe8IOJs0p
UaJj80ijM2egvTZw8c9tQqvvkHl3/Xeg3hbYf2Qzs/gs4NB/OL2A8b/bpM9K
OhV/AzMJNRAPDzZEOiORDxNo9+gcJErvU8r2/PhzwtwVgKKJHBG3N/sTFAfz
gPtmcpQz8z1SMTxO94/7Fo7Dzm2zYsEwwkqh3VQJZmFEGg9oTw6jmcaXaizI
U2cNF9lAbRUAragBJRYPN2ImQgekyoo9Xzt+Ydgo2UA1/5ZFeGHJ29TTKVwp
lGr6ydafONPcBSyLyt6hQxqo9GZwvqt+Zid9YNlvFGxzGsxn4YQAiBtwE2vx
jbXSFCVDYPI5NSTOhfjn3CCkqhQUf/dVRPRAlECBA6WqTvNxUzXvtYvqmNaj
+7/7ZhPeLVURObFBoFOfsp2TgEx2pp8t2VDjiMGA+V/Mjie7wnQUiCWrO9CT
2zUEB6IvOOnxcx4SfnX1EzBHqPYlpdBOZeKs/q7gQ2uCIwLcbmtX0tG0dC7m
6+VrZCzZDaZheYEIcZ5PSBZIw8YtCTIUqtNHy6z1f/rPgrJagHSUcb0inoKh
B4Khc1DlOoTFBa5M7z37qbXB5jhxovu/DGzp8dVo4O6pAj1dIdUPVd2nK1g/
CMprR4cLvto/SPS8T5XG81GfBwxwEM2mldAxAkC3kpJ9GAi+vU3o5jyQ44Pi
QYpEa0bh2ZvNmb2bDJOa0j2n9IOaxVGa4ZxveJcisto1tmsRfzCE8Jg7Q7PQ
gX8ARRhyFUmPUReDSMkz9lznZpk0YQecoM4RiaHrYkd8b7SZx9uEZb4gfkrA
4+6oRpvKBlsowc5rXmUb0WkZMNGAU5+0wPiRwD6mljvreD+3wISVwLMW5Uzx
aP3+RhSrBunoFN7opSxGWUXhSwFAG2eyTD4RQC2BsSXXcLGcyD3q+KzXTJXP
vjI0THdr13/LnqF3/VsjbuSSlVjFzQM4iV2QMo8VjdSFGNEx99AiwzyTtD/T
7KTMjiUl55JjZ0sB1DXPi9OjoKV+7jBBFZ75Wev3lObggtvJRI6HWhmaaFRo
7IX9JT+OAQVu8LSYsOXBd2MwvWyvvtZT5WPBE7rkRJdPY/Zmz5FhWhXRFvMr
tF10H+oqWpG4JIqTfVj4O9pFQG6uXMwQs+aGMu190LDFr8Zhmfdoit5P2EMw
pXjgcSes/XotHjX5odHRZY1chd4S6/1cYHuGuiL3LrvyffARXKJgc02vZ7rt
PyGEni1kv/7uuTj7P+snGl/VPE0FVONViTDpDgG3ca9QONxROm+I/cVWNRO8
r6uiRrTcrJ75TKbNOgUrBNUiJdTte94cJqYherF1DIFaLOqviDl29v942mMk
cxren//h5zbx7Pwr62NP0SOTxTS0LiNBEUBqCtYkJz6Q3LOZP6/fX9cJtqZW
Bfes9Y67bz9RmCuUBrd/co9yFRKZQPZoGnAJjzEQ+wG+wuws+qQ13Oyja2LY
soK9MAC04AUmMbUrjgCkNEq0G4D8N/H3qzeXX3QDLa9xp0Vmt46fTm5caFUM
wNwKZpvshiO2IcL8q1C2qWJn3CVtKdfu6RvV+jZ4FYh62xSIkkorjFcxB+La
hc/+A8xgTP3X7mtrmmD9ebgeGtq7/koAc9EjMLjU2CAoY01/QsQAvwYneofI
jisoQcUc7g1tN9yqzg8exbzrxyC9TC+W

`pragma protect end_protected
