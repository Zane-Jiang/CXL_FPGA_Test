// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HzA+q7qBBaiQN4tqlpRkoQRHHQIiXXZZayMVXgiO4dMYng77vBXoppk2qqFw
ndgrWwZkd4Bo/Tw5FDLEbm4QCmzPdprQysuNrhNR9rSpwZ4C4b4GA7nmRe7t
SnLNHNfTKPmHojzgx+3tMRdI5/Z2HQJZtj+/BRWBi0sFBszvC/y7bNBbQqJr
yrU5X1/P0EXoWNaD11E7YxPUc2H5NwePp8wEXbCoBMqXnS3c4RX/9zC7TZRc
yZgM6teO/H4wxO7ymCfW6bjZ6Fxl3TnHsq6bHGYLiNyHBLuWPizXuoziGvoa
PuOmWPjTQ7x/4UOheSLHHxsm0q/jwfIOLbaOdAwPGg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZsGQcY+961oFBohVxjQVu2H8WgKVQ+3pYfRk/Ujv9e86hr5pI4AnFAOAiMPI
Z+b3Jxtz0FQlcEHnBQLleTyT7uGnN7YUucveCwXmnI3qQCAQcNqZxWQMR+ya
VecwhiiFhLWmotfeJDyonzP4z+9b8gyYeORp14r9dRoccaBCq+Z1+C4tvve7
9KTzj3+i8C11HRmstc8pzDZkgdhoznMHdmZSj3XgTsGEatC7rooo2IFs70tk
m2tVxXev9GObZSv8asR8kc8wVKUSRt6pM24BKxGNEQa/eZ47nqoafQW05X6i
Fx60wu7AWt3lRPkzzHvIHQXSV5GpjTI9dPdwGZ4gIA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GJiNQaCAlq0nPJ43BnPyJbMXrT7CJMyMLWl3lbh3Pxd7g35Xduou/DqXFgj/
8IzDyK+ne+z+j7z0w0Nt69qPgU5GEDfT/7+06+teWSYLaqF+dv7UchkaNUjH
bHH9w5pjuWS47TYr2YXvKgjmFcvUoqCjrKA8Dz34ojSwuBOqFa00giwnUeFw
vYPFU5W73B9XH/S5XBLCWmxl7kIuIzxnSNyB59Rs3MOPZDVX1baG6VFqJpHJ
+vKZmBRm6ibFGlDOJXpwNRjxeosttf/Ac8RdG4hPvqr79Nq9ps4etl0IuSG2
3I23mzVREeGstLpw9NmA8KNmRz5zcZVNgBwK5RNcng==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
f0keXQ0i2scRjffYOUE/FUx6tQd+EK0iGE7nyf3BVPUYwmaRjjxL8rsbYa/5
xyvPwjOyztYz1I+0mJRJHm86Amee/qK2hWjpRZUGcMBXsuP903TeiCnQiDkP
a1QCr5t5yv9fppeisalP58uZNBnEA/0xqz3QgbbLu9E+rF5G4dA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
M+ezqmHpQHROhgHAwpljdhuHwbC05A8n4fbTaX9v1RttmJeR1/UCnmoTEfK2
UYZzMEGNMCeDN2JHkmCossy0j14/2MtIwdFHw+QGoe2fTxTIlpoECQkGeNgc
b2vEJ6WpOrR8rZBB5LuGnIYwS+qq1eUlaHQxMNCx0u9frc0egubyIPq+3uWL
mhtas5Vfqx27h8IFkEr2RsYOuGzy3nxBJJc7f2fS8tdXhuLtUKgiRl6qVrRP
UIlqPQ5q3Q0thdX5ERPxc0XYMp3EUtohr0BkYdovk3PrAPQURi8AWoAYkjrd
/Cbrax5lhw4qeTmxIF/68rcYAGqgRuSGjsT2q8QNvts3Au/M84esO8/qoFft
DhJSj6eBN7I6MpEzJfF1KmMWglA5ILcSA/uI+hIFXexMHE5SiZwJB0Aowp/e
lmcw1JzVjLMme6PPanSb7vn8kGz7EEtSVUbP1bJ5AeOzIoR401h4eQRhtKRb
A/+bRFftA4ysvOdIqbLcnbGSp3oPMbe0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
etQhtv3yLE8x4P+//Ti2gKMpodlcWjqkzgvP8RChNuQ9ktRK4vOwhkTzIw8/
0DwMe2YV6th5QmS4rAf/+b7mUzikxoWDTpQLFlRwYB3HhSKhSZYO+7IoK2Q5
di9Aas6D2tv4ruwg5DJ+35AdMPduu3BMHPjn5e1r5ML/FnYMUYM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kZk29f6E47SfVzZNCcXarjwA8vZ8YWhaSzi/DFJzbv1AeE7CVDVbaXA74TC2
EzvBiroNC148EFWjEZ56mGQjsTitBf/cBhSc/kXCEyNJWf7QR7YNuyz32QDz
7jXsaFehofVV8LQFmH0txilt3RB/X7AoyNLn37g2sIrXU2ZRZfA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 106304)
`pragma protect data_block
pzEPErI2LwZvaOb0BR/BJHyRpzPZWZYCJ5fTCDS3g1cMgrDgj+It3kKSUqbn
YLnnCs5b8veSqv7SLBwLJBR0QoTrFGsWB0T3Kgsq9TGWERalKu2hbqWJa25v
FvFlVL4h9dzu6wm7z4FVSw55fUTiJhmql/oY8OHjq+gt0YGircSPWZ1thN2j
Luzku1lETOecps6vlOhNd6jmrFoxhevMWTy0J5rG7rc3ssUn7bIOr9AqOVI7
+rKRAovU1gcxjA/EkIc/41a3/ggb5t43YzCdwd155i7cF447fiU2IlO05C8J
s9/tZzp9gJgiG8LLFRCV3MK28IyrC3lnr3RQi9VRQO6mmWSi3waG6DOBCQG1
BUyyFvMFtddvshTjUgdO+9Afqm6CVDwUJoc/JPFndsZYdeT4bblMJv7HC8A2
jJ4C0a6SDXKonoq+zQZjWQgV4M3KQHzrWCB0FR31wgV+X/zyevVCazO5vdKS
fYVPcXVT9+bpe1d3xrtU5Oj27DHS4kzaJkTmGScAbg/v3E5ty7QnDNOPx+jF
j0OGPXHe9KmNLMvx6RTYRF83yEFCCX6RYlyg0mKFgkPNIy5NwJbnnK+WUrFS
4C7zSFvwf8XG+BfbgJfIv9g9umaLnuwh+gON4cRBK8pLgHUWPhJP0ysWkJWG
RFoWwgUWmqxLQdqP/JSo3ZfzjmuSvtfbhCb9krzDFOupRPXCE4nVP3RroYIC
aZ6+5iwy0Gs0r3gxHEh3FNxJ2CcL37v7FnZ6lDpfGi7qGknSTnImnzbArEWj
q25EF6KFIwVB9XidahxujaX541szPdsflmsZniPF+lnZgradGrZM/pt2Cz/T
tSqdMkPkHiO/BYSIV/sV5P2cxs4/zIQ14CM36lEZBm6LWYsyDWb1KYXThoYr
crrdykkZg/L5VadmN1QtZBQpmWt4lZp22gGFg5Q1/iBsAt2NPWWgUSZxEMip
NCRQV2bn0Ic0pyfCp/ywWLF4cf1YEQeHgTIYiWB5Rbxi7pK3JXBJ6buee9HT
p/7Me8bBIfkuh44iH6E2A0EovNNZ7C9BXSSCfGngmFGOJvhFG0/tEBSyhacQ
eKmdK/jB0spUQunko27D8SSZXuLDemErDrXLFUFitd9bZHM0ULfTH3pjilTn
71sDSJdskxCSW4SS/0HyaTjq1Bk9pT/e0oDSGKnIaJXqyMahhNgte70RlP0H
K9IVGlMJcm5zqX+P0WuRJPBJ0YYlNDshA2x/h1gC6uSk4KHANGB7g56mIVLI
xLyOE3bXB4IQo+BAkKO4MXFBKvyYJoHJ8jaAV97QF0VuHMm3RNjSfis7BtoP
uHc7IS6AgtLL887lAUBTM/NrBZEw2NVv8wFMH1dfvd0VkTEzo2AQax+Y1byJ
qNvWGnvJswSnUGP6hEzhCjfrTgRj7rME1ZoOFgM7sY1qNHZeuPgDZhOrkmiK
Konj6xVGuxva+rjzSZNv+1wcXUAvLbOlgKgcv+AAJ2Ls3vkWWIUttVSrUPLi
JO139k4tf6btJq1w2dCcNhS1hN66OEzYZDYvmIUbKCChFsg4XJRXwk9li1jd
ywVj7xpos8F/+J8gUqb5d+IsIhglp8nM/lTY6YIJf/8Q9xFgVnbWaId2Zh4F
ApXiy35zABkyre4PeTSb01C3HqFbDmd2HusLTr5sSnVqOrRnmnHZbCNdJOnW
Sr7bWGgAJtwt7xtNIkdIzWaZ2ZkjJVx6c41/i5ERNYMWNUUGEW3fsT9Ivucu
IDApUBmcEs1OUWl5iMbYaMJHoMQpI463+OujcW7ZlApdwg7xVnYe72IMTsLk
4l9pcItRcqhvG/ODcQn060o+Ckr4m8qk2UBLiaT8+eNKSetpNZmS+YUfle4+
BvyOuDFCHCXzW4nZOwioQPB9FG6NLxld80BjE1V/n3ureYwjAXvY48JLPXwz
eDH/BhhA2EevjxttklQSEC4qk/zcflFWEn3Vtx/WLVeUfO5acLL5xROuNRid
GyD4e/9RsZRC8E/iOr2/YuzKgJelb5DuCP/0AB6AIHoIPrl/zROFm/4wSHxY
Wl6qUk32eHnbpusQO2Rtoy3YXPf/qIGmWJEfNynyqxF911oryzhVTszzHFUo
fi+xDtY8TL2cuCLembCspu5zSy5PINzXjGtoQJUL2wPFDXct4bqz9KOULg26
ZAcco1j/yHpWTiQpZR/RXOBknjIipQjZ/WuQalJQDRvi+Z+0Vf412ddEQwZU
qxu5Cln/usNtkJdQzoWr1p8cpKLYzenEB/wJdRhMwGWVDWZieN+uEGUp2Sb2
4vNAJL8cc0ErXRIWlzq5pvKHjv0BBxdjdVZZ40H1j53bBc+pkD2hAWIj8lIQ
KGAfEWJVnoYDxQQANPeeD2DSgUk5IR1Mfw+7DG3DmgbvFhZF2zseiS7L3ymz
K8sxi6uM6JO1MGM0Bk9KlGxlH/NyQUWX0z5Mkd7Tr2RmlIYFQe1e2D0ptxvB
7AMKX9H6+kLfHl9IvIIvM2zYvQxgmD5gc3wZdxe0d+1+MvAIVA7fL2AjCziH
ZhFb3wBm7kSM4GZ+eMuAQ0c5WMtx1itnfesqYMbbD5F1lXj6RUhqfB6sCZYZ
XonkaFi7Fr0QC3Y8xHO1HnZaIXASEj7zYewGtp2cmPt7jchP1MVFGnZkr0ri
WMZg09bNRBhCqTn42EG89hkEU5G/O0HRWiUaJbwgBBZ/wG7EoB83orx/hOXE
IQmzzVBhFQIiQTCOQizJ02r3FgrSNMp9BvOPGytsNU236utDGpSgd7iIen0E
i9GXrucfhIRiN4hnKcKckhZoVW4RR3c/sRUIPChDxxxgV7VYa3NEu+S6vdsL
1RMfpPBAeh0DmBEGoB4+j71lDYSlKu6cnQM3sTlLT7Tq1KtnF+VVNDDhy9O0
dpaNgOmpt+aSNecmt3fezbU/UDWXE4op0O9yX8JdF0Qc/Ql/o5dtA0tJpD7H
wPSmCfuYPtBtJGc2hlLcTG3RIJ0Do55pec5oyA/79k2Kna3H0yHwQWmpw8hI
bPsV0LIkW/KRmSMyd23TltrQMCCayaSvHG63fj4dnLojw7wbOLpiielZvGAU
rEF5iAif5YUpoiORWx2MLz293JiNiaJHejyOSKJRn+0ZND2jLUOmDYBxSMh+
77/aHUuaBOgG614Fj47bddzpGsaF1frmlklsyxxK8Yzk1+AO+fvwq2mJHrL7
Iszf48QpwiYtb+huX0ctAI3D9AgixmMg2yO13pboN/tmhhR9KP70mS6jKxzo
nxIGewaeIeO8g5103nKKz1F8KabnqqI0cUsnHOKHz6MZaV5g7+PBthID7Y0j
fx7kvDZ+g1d9ywcd3+0zvuYnMAHVKWT2Oica50V2C3skEelYUoaAkWx3OTIa
gnaKDHHXnekxOX7S4h+RIMIGe8+1xaXKnujgHstifCNGt6Zcx20d+HaM6H2C
/pW3JQIFqGZIGDdMJydwb4I2qj5ObyXB4Xm9yJ1GabBQ6m9sj5vWhHElKjsW
AkToPhM8OfKbjJbMVdZIMmEtm1yrKa9AjRAxegOnvIm2KlkEgg2dD3/hmhdX
+uIcGmvc7Cmcgtt74+hzPEHq8Amqddnnri+joUgE78z3zfxddGhh4FCZXZw1
o192xZ+f+5MmhpC4R8kuEDFB1haHJoM0dvHeEEgbS9EPR9lsfcMoye2uXY23
dhnSx89g/nDEGEOpgyR+Rx/iuAK8GARnLOmWlL3UZgFHUttgtFU3eezjPUBW
89YKjW41pvOCQkoPwgm4gDHHSA156o0oqOWERAJ3Nkh2L4n9EHZsc39LtMeZ
/E4MBNlX5wYza0rfxQS8Hyib5Wn3CMKAwPIctO1/PBvYT0xh9kh7EXtZQBUm
ssfCdEkYMAe1LSEYQhZ832hO+dB08ooFtQ3U1UaC8CqP7beg1FzsmToKlrNF
pJUbaNLYRb40al/xnTaVZjO7AhOALAu5BFhF/QBz/uI9E7wikAS1BETGR2AJ
YOGTjzJAQP+vooTV2Z2IaGQ3EqHUiT3C3DA85AJDsgkZPoNITGjoYBlRPHN6
V+Fgb/Kwhc/q/5k7+VDHAyWmZxefIr6ZEMt2F4mJjE5bN65SpCyXRteUK2TI
yAqJ+pZ+NnBiYUrWY59jiMM+FkDWK1cEODS5F1MHQtOorZPGSht4YA0dvino
XQpjpLj8kHSFEwLrYvhZHzrL/SFULJVf6kn49YC9Fh+GmfmOMVy/ZcVWTyOv
ifhLQAIGmcOqS2uITvtLP4aPWljFssUl7eNo6C9/y/knfkhR194r8PaDOj7u
xbH7hoSrhkIeCNj6DFsr7yyxTq2zPhehQnQPz2djFX4PwhEL1JYxRKzl+6LF
cZADtpuTzp2lP1aGjpF82DGMMeW/qnhmBmxioenKPnZ9ekPI+VRPDRq0hD67
kQHqRFgdo6Q7V6ta6QTJaRBiKbmaCzTfAvmj88ZYJHzZXNOxbH9a217l9/AS
ceGclQzGiDPweoBFt3BPyjZoed0XztHH0Q+2kZ6yolYaGtq5Zy02HpIUEdcs
Bt1oV0BOj7VHS4qS2OuxOMTOSyQaLwU8tZfmWvifFMgcH7Au/OR6owzvqmLc
g3pX7nECCp5SlotUXmlS4a3ntF8p8/KLaxflnBmoBSVoUgsrDDZy+WOJ8nfd
y29tq2pf6EHrLVcGT6icGRSst4VbsRoTTzlzeTxKvWvVchjR7bGoDLf5ozDS
NqA4toGg178aAbx3xENJDZVhFETWvWyjMENV/iM5mapWDfUyfLs7pmANIGgo
KOpzhWKtd4pR7vUhSvAY6C5irCkzAsvFX50Um12jqK7mdDcU81ulhZbn+sWN
D8m/TFawkTZFoJYLgF3V+TRyKBtXDhwxuZ41DbZufF7wW/Kk3XsSgCz0UK62
xmyNsW8KqOe3ZRwV79we6OdGkVtMVHVy61Zdony8eirToSjRwTeOj5WbGQQV
iZd3N/EGAI3WmrxNSAmy4W1e3A3IvbQHlsXNU8VnB6pTNhqjQhrO3TrWM2rv
W/i/xlXoQoxZxeO70Qs/H7twauZ2+zLde5ezKMi0sv7zRp0lgCNKclAKKhUg
BEZKPWOwWDfxZK+AV0ekWK0mVxaIrBjC+ifyeNKhGDlndq5qGrvj38NV/xNN
/DfL5Rw7ux2bv3nu5TPUaVs3w9dmH3UHBFv/0Vg6lRxgYAaaoLV5kb2uwbDi
vZuGdHV2x573qgf8VU//eiP7Ln8Oe1/DZVhIL0fIB/H+DnZh0/ADvypfOwqE
zKiW+28mL/e6VnTRDbn93i/bhuHj9ZFHGPL4sTColRSiaDJCFP0OEmnZpZDF
Dy3syH+AwevpDkIFlWanFYdOnDKH2tkoV9h6CbBrOOhi588MemUJavI7xYUg
HaOrIpggRd8sJ25e/hba7OXMVKvWlRnTrM3+suRdAbrDvzSc0UGflJrYLnjF
LXYC7qaFgzHUOHCBqcoK7wreDQ5h7MoKwsFfwVm5TjGaFsFQ13eiRrNstl07
MeytFPmZVwFSYzVKwr2HwatngX5YjWNe44Wo1gFhxIr+j+czgGy2X8WegxXJ
1XYJNfrh5jbnJwmvNzvWoIo5u6jqFDvKg+3zgY/wLsXXwr9SPPIjT134fHVt
8nu66f6uV8pjoKJwMYKpOrFDFBiRGOtffQckwFmAMV3sOSx1kwSN9nBOAR9P
Du/6YIRhQ0cvgfU0bP70CTG2Tyq9KjcLD7VByfM6t2DH+7kckrdAZ8MCtnPF
HGLbN64n4+ujDqgL8QUnibJdKjfXAK38imhy4662v/jkMyudDF7HFY9lslAe
zf/u0oGQ5GZ4UPExVD9fnd2QmYQM9Edm4zR68tu8MBLIPecvHV5aNeMe4SO5
vQnBl10zKgRWHv1Wn+5jlwYXdbXn78U/E3+Z+5YPr88iyBqQYrc4V+zqNs3n
MG4Ki7JDVlYy1qWgblQnqKdsCYJyBcZ+VWytO22ehU8j7oArpRGIkIkxnKFF
FasyoXnXkLkKYyLz+owUhMOJ4h5v1lAcafJ2u+clEuSMkXzz6DsKyXjy8Ux3
MK58BOIS+WZVHmCXweSzmV5PeR2BvRkMesMz7fROH3Kt95FQSmEGfopoePMG
EThqQ0AuQqQBMqR5yW6eF7y0zO1+Lh8UlQebReXnFlktdyQcn+KnvwKGPVci
i23aqa4fa3Rlqt/oNxW7PWoY0AwshZXCWJfGBZoyTePYUxcwm2QIeM4vM4Hu
JLH+xQNIiNmsLGS7hdXU+vbV4HNyT2eL7PFkYuxhG2bxfScy20dkdhPncpMM
OiR8Dib/wMH/5pxg1DxDiPtdWSDvaxCIdePUn7ZIc1aaQxjvMemAzcjz08dQ
/ePSad/OvCS+1+XoctU1xiPtQ5sDZqAiSPEHLviK3y/rByaz7RKu42lXHiRG
YEmxn1acRFKvvq14ttp51OfBGI5mWcUUEI/Fip2mROf3Tc166kLl0oSFGqoM
c79nsDuCNfUS1J5Yg72r/d174tJHTvtWNjDdHZesy+fniVgv+haZ1ic6D10y
Y6lBgBVYT5ffQ48FDz/A2dVctpc2F4Zh+70zMeQpPcVESg0+5f30NQ5GedAs
NZDuNcPRkBus4drwHuaFKExWSAbt225s5sTvjnQmeJOBWi1KUMMZMbcM97tY
s5Ln4us2Kug39gNoNr9E++PyFNZ0EDh8uJjLOoDoYB8x1wYVt3w9p8TTpsB2
ALGcytjEx3qkV5uhnypyDcBtPI+SKuaQNtOOzyWA0DwfmgDSz6iWmlAysbdp
FM1Sxh4dP9Qc64O5XKz58UinQSu6xokCbUwHDfmFRk1WsUSgp0WBr+tLAm6+
0iEOEnhn9hoiejgwirdsbYoxo+0U9dJ6+DDY7b/EgpxmhVBTDg+KLUQTGCBV
3pk1T7bPnMsArIC9am8S091niNojnBCtzUEc1xcM1ucnKKXJeVKAq9k+znta
OK2s0p5YeS7L3nFFpNjiQe0rV0+q1qMv3lObVS6ozwHCwLWpT+RRXqVxWvq0
vSMLgmnKl9EXgbGr8cXoI2X+G4KDYjV6/4cQqZpJfTdZZ+pgc3qW0CBLm5My
5q5n5Cp2LhuYRzXNgWsFAas/F4zaPJShBm7p6jOqnoh+rvN2+naO+d/N3hEC
9xSWN3JWwfFy3dd0zCSiuU4e8IDJ/4xWpObVEt0hfcHidtQaB2CKQkF3RgAS
hkumwdqwlBmeqei6iBkukrOB166IICfCGJdDcuYPSseLf6Yl3i8a1T7WPdD1
WYo8JMWKmV/QDi3S6OBlDiXaRDwBfzB/qdBByxPQ0nfcYIrAWFBBXge3TX82
jEBBOsiP4t8ZGnHYYbIjsty+lDKJjfkDC4sq+D2e2bYvN3Fj39tTNvaaLRKD
5kvB6jiK3bjHqMqbI95I7xXKmRHqxZYvEXwswd2AchImgPt/yb8fZwOQytos
hNsaayuJQ8aYLUzq1d590LzSfGJJ6ctigtcKaNvO/NDaj/9O5BsIP6SOkLwk
gYjPLVxZJQyf5ZQOspyX2x/9kOPolL8RoVD+DVlBkuSRXDFLysIp9IufbSvC
BrY0hbtMOk4Z4rKHG/Eq7U7AlnqGJCGrvH7UU8yPDskiFOpEkLZHAKhrK/pQ
CkrBD4sDq0ZG9lcTWd32tvLX5G3KAsfM6c4ob+lev5YR/a9pW5hjGGZcQrbu
UabFJeyw++1r9wW0Z4YcuXAbPCz44ANcNp6ukA4ClYakLWVT+OoA6UMlH07U
yCFkz7B/it1jcXLq7LRfxLHk96xuBtk/911S8eNdKfRqrmpzltknX3EBFTTV
ThXTMpV2fNVus2otcQVRim3GjMy7DIV3TFmTyebSMkxdyp0tbltCEe4Oa3kG
R7u6IyWRpni4rxiEl8XFpb80/S+3KMQK2C6arl03y+sraLOJkcsdMRN1svSt
WtMiQp5/+1qKJmYqFeqLjy7h9B6GK+8XPw4n6qvvhuCR76CevUz6lTc8X2cm
4QpOqsyRmtaE8qY8+/yKbILOtwNL5HFAhHVv5wPGuiffxxj2XlsECIiHRE5P
7XfkSLtzc6HPtM5YAz6um5RhLTBmQAbRs54gLGucz5UG4LCYpSrpp8tBhKcd
gQYKlvjMCO40XZ7RD0p6vAxOST0FBc0Yi76YllKja+4c1hvOtj6yFBxoNugH
0OivPgixCZZISpQJUnMMnBICPZ7wTzAFY2X+LvwnHlTmpcrUBSO1sqq/NGFj
uoMJl1TUygXrYhU1DtpSiX04T/C3VDV6TXWHXVYAlTrHawUFJfc419728+Bh
gBZkBunSRXLdEgX1wAzTtic3FN4XPcC9gw4ew8tPcq9ovk9DQP4aHqRCfiBN
lEIsZH8sRNEJmPfuFWlBKmsEAadmH2fySCZv0qe+qpfpH6I1wkqXiXjB0uNY
7plGUgRV8OwdhxezpqNgK0BTTJKHKrsiRl+cNyjAt0ewllxtUeEU+17oOIJ2
ahUONhk17apwtkZz+Dp2OshwBuc2+Eg/3Bb1gxqbk4WRNwXp1ip3Vxafd5Zq
Q9YOPJaAfHpS/YO5BTABhOVrgmzqkodMN14AWlGxpT7f9xIoEwBDmhpOpqKB
06o99cbXZ3j6h75rKIlJYCNW5+srUZpXxuqeovBU/HQUWV24T82NpNGXKZdS
ABnAUPlNAAPPVghS61kOF1ovGIJQxLh40hcRmblZgXzf3xAruJ0Ord6eBU3f
X+ItYwGR242fM+klYRnQg8Gbe8Ad/xV7ZFYQ2p5RWbZLpFkg1H01aLwlzpT/
u3Le4CocLx9gvw49WdNMYQGh22EcUeRgvpvpt9Ico4cqjyM9msCbY75wcOSA
MUroll34pnHnVLATF1StI5mN/rDsOt7ppTnxZ9r1HIlXYfK7UyDdlk2LXiX2
/JMllpCFRQ0fhJa1Y6TqE4IBmBXxcxVHS/EzVTwpQqeldvo6BQi+rXJ5IDb0
6FoT72YgTjeGp/SSaA6TNaLKLt0S9tGQV5W/YpyNNqs0uJ4H1rej+b2KAx4F
E0bofrkiumNqCbREbkqAjGhRcPu4jgMt/rK6F8eF4Tu+t88oroAENZ5t5Qbq
1gtn3bTccIewW5iKUqDWWGTOn7VvGP+mSwKG+oq3BaccXK2bi78O4yXp7B7z
uhlG7tJdI2NkNpuUZmKg3AJ2l1fwDIJICgzLpYgfM+jhU9E9kCxyHwHzZyJR
Lf22a9Zu7EOhlKkFh5M1zmWdq8k0tBhs/ZUjDtgAF4c6xuT/iF37i02tS8Q3
MwhWE6Wo+k+9g7toLCkzwoQREFbRUWTfEXt2SuWlybI9BOz/cWNxWmz/u2GI
GprG/CzoXiwOr8gnvXziBWBzATwxJt2VupymN5wHbLJBrA1jNFPaThT/eF5A
DP9vixnOHjgc8mYALYbXIiI34vdFlPlJyCPcYRF8vY1ZG3wxKNARXL9DHr9t
vQqK33WXLP7ITAjwbevLmxQWU/KnovmdSeKtBwCCvnIRUZ+taNV0qeDwyMQU
l3iIP54E/LMzJCR805FpJhkoES6jXRqT6MNF/NTOZDjiS94qO8AZqmoOfwng
25XyXN3PjH8zsVg+tdM89gyunUYHYUxTuH9NtVr/D3XNd3XQtz3irq8Fay0+
omhBro2Ou9sulhlV7CzKroP7KoAUje1sbih7I6DNu9MZVgs+Wv+tuPE8cmrn
ICt5Vv/MggikcnjrJrWkmQRR52aAiiFrkAJc/Z3/+ZPvPeKTEEbdnbi/dIr3
JkXd5Z2n2pdt2YWvvrEZKoqkiOjZXTvwnbX5WVRKvCt2/6LeMrl2gAn2hefm
hpQuGz1hFIDT1TW7Hr4KxKI+5wZIlla79fDAh+p1GtcBgp7pnVMOlNbdVzu6
kU3Ft4VPlpyuhg9WSFT2Plvsw5rCFwuAer8W+5yoV2VQmcy4MpScm30Qo4r4
VyITKpcfBpLohlXnR15y4uThM8TfcxejEZFrvTFgK+uTGNftI6JPsNtkOMUx
iQjSU75NBAAM2BdTOKv7tHQED2YCQN2HItXmT12UqiWSrGtjq6e4xp19BeXq
eI+V2JazjyI9EGgzD3GQI7/K09/kmoI0++21gz6RFGN7TYZesuZr0/5m3g7e
gkpjmMrQqxPtwgQDQF2gQt/exBv0M0tIAI+d6NmUL1fl9xGu6auXuB32q8Ju
RATwP5nHSnvKkBkSjsk4uVu+24E0QnaWfe1xIdGBTGsnPMUCYYlqmR40RpZe
O+cBvWS5mAUgvDfhvlgJwMpPAtMhybnBJLJacbZcMAP7OECX9l6qrQdwlZ0y
sr4BDKOP7RoUnItxiDbv3nXscbAhb5Dr3FKvU2SQYFbKA9kJS79LnraYMk1C
qn+/BEwiAfhk5qNqffwden5Uw+vu/dsBnBzAs+jn50zHmBbM5Yg7mAzgT+Ou
MJWiRIB8gtVXSTHjWXzBc6X2YxBCXZs6eXSI7gVuJfL/vAwOeU3gJ+JBpPix
ouNNo4SCS8jxK7tTnLSSsBWgWpR8S7hIkdTo4oCYHdDGkLkP8NzmlL0xrWcS
9Ar3ow8DZx2LUU9m3sP8mSGe3TiTQaQg8fqeXb+cyZARIaJ6Y0eZcQAo3yBh
wkGd815Y9GNinwA9RSejNZs1r6h90soYQ44Dx/mrEKRHxw5CbLXs1cbSXYYG
JJjNConl53MeuGAuMLhEWcPdUe6HwX2LrWcppzSAkpE05d6TyHkDJNe8ktLa
Mh9/gVkNBd3yepFoxwVtCh517huMrUuYGV9UsI+XZDX3oWpLrFYfduAVcevY
9eynEeqXmuVZKW2G+DLqM1r9P3OBZ094G4d81wkIWdCBsVvylAJ65b3HCw6O
G4X1a/MJ1ae3H3USZ/lUN8au2F5Eg3VpkDOKb3kokwpGIaZnsNHoaIZ7BRzt
eJWspfhm2qpWBsSA81qQkMs/zH5myJjzOeoijmE+NDFtJYopj/2FfZNm2Hwi
2L9aFbVWErPi0e/Jo31gWTgC9ugtoFyiJoq49YexmJqUhBxwiJFKwCF8ZYxy
fY36+5cgMOxLxyPYiYZ6waML21RmZeKzUVrbDhKngCsKzp14ITcIvSieeCUw
7WnRSO6BzUpfxt6GTKH013HJfI98Zbeu7+gmdHOSkTz89njrN1mP5XMk2zTa
inNPVxDcp2zwbLJvZijnw3DBfCG172ga4vZFvXBeFbK6LVrRQUJ0aGsYclpg
+g+Om7EqIKmE3Lj+Sn8H+QRkxVKxu3KI9rBeThTUNmVvTanzR3ZeZ0K5W3r2
PN0Vt3SJQi0KicSmZlJ2l1Q7VIJjbqBTe5j1KalouW/E4bIEi6XXd+KaHuat
5SDfQI2iKAW9grGl8m0orsEx0/xLDxARfyNkHQGQdXr2LvmPaRqznQ8N0cFc
WHiKg12GV2IKIQlQHiZPPv+mz+CpI+UFSo4MSmco2SXPULcfeloWIwj1QxAp
7wBh+DCbh6KTtQH/CmueKA2d2ObHVv3KN4u3SHoXonTz+jVNY0YZ36wPrzhU
auJ7bNsGbAtn7m9kAgN26dIlZOF7ZTMTyc80IzIrDjiUB0x0RIsNej+sM//N
r0nAJ/KIl5HRJV8QBxC/D2JXDigk8whSVqUdc3E9z/gaUk0IPpzc3+UNh1pC
wq4kf8DeHHFaafjz3HKsuSVTWv+VelAxH5OxMkCGULvar+HS9l5wTYb+wrsG
ebm9l1ORxJX7LCdWeQEVDqXASsxGkv5omJ2kPwy/6nw10HnUUTvnNmRnhMyE
LzT9Bb5AzwUYYxOMWlsDimy21C8PNSwclM27F/6eiOfYTRKQ1WIaGF9yWgax
7dI29en6MvIBk64JHbKdZHY4DgYJaAR144hWSykAwrHYK1eMdo8vphhS8dFv
YxsU4egmfwqfDBWdXjuVm8V5aB1WnyJpVgVM743E5z1bdkKybI3Jne+U1JVX
ZXcNmHi5a1Fi036TW3uVHxsKQlu4feYD+OKdtjwq4zUzDvd2XyDN0SMDQHxc
mk2C5kygymECHR0XPeLQrOQddP6DhczeS7FnB1letv0Gubei1myGd4O92OYE
Wp1lTgn1RNqj29vaZvKT8o5EPxKFRyKm75oaZmXhIYOUK2kqm68lhI6Z0HpT
JFJbBM6dskn8MzV7U3RsJ5iXKxAfyroiZlVkA43s3Ka1jPSG6FfwgQiHiR8V
iRzn44EaUm7O0trzj1v2CT1u7iqBLadpa9bhykjhwWVsJYI7nodDEXvPZbCZ
Wxtc0vrkP6BDf9QZ57NB9+/wk0el+Fh9joibwCUDOos2zWBJKMhBk6Kjfkga
XZjR/dGVwYbwRtDvIEAzw9+moVhx/lFtJbIcHoj2jFyxi1/mHdQtmBQpQtQ4
OZfqVdrFlcNYCReecjBCLTKHgpkui2S0vvnFW/0Fw/7DV0NN98JEJ6lgLcbS
9XGgHv8m7BLY8vQV/MwEwdTcZ45zr4z3E8sOtMWxgXcpaLkUpVJgCJEAWqU0
L8DY5PCtSCJZRgTms6oF4u5h8dc5lFDIk9MtaKJyg4WotllaA/BLjLXrwJC1
+N/uAtEak1yk0uS792goNwmyv7y+lTDKvtl/EWbFLDcZsKjQwych19DdhYsQ
afan8wQVFl8Ibzzybn0xk2eDF8/RJBzwdzawm6Fc+SPGaIqS/8gxUCRphMVv
C1uF/NbPEyNOG0LQfD2GjnCdyJi2lky5MsE2o26LHelx0lr8U4kRBspsOwNe
8AXbPqzJqhu06u7eT/8JdQFafJ45eTaZ9eCCg3ftLDUKXOcG+/TMsvWKxAVI
80r4l0U+X0mBI3YDB3vHH4DkkWuoLMVNMoIFJ/Cj459NH9GWhK18ICB29JLh
h10yqtZ0Fxsv9DJ0W2g3IdynzObjiNlDE5SRekVw00B7VDP0/yGZIqtiEDpb
rkN7GKcPEqSZqNo8BEBoE3nxeOXYCv7cPY+qbfLl/ZSGSCxkMFHnfpu1/x95
L0WadPWOFdF1J901q5ygkfceY4gU39g+45vS+X+TxafAsHJU+XVY95TEAaSt
wwfByiVMOAgIcc+B1kvEdrmQsqojUrSguVjUn8K7Uk5qn3iyQgkc7RDv8fka
/71L3mzvPGBymPRyBSb4tfFfRuvyCHIm3pzeO0iUQE3KY5qcgYb8TaSIDjn0
hIz77A+R5WCzERcnPjk/yYHHpHN2fYoyxcDQblznxioDUFRpPG+bjTO8peh0
FWoi0BIanChCmotj1mTgmncC1cn5MhlmO/fILgZUWc54dSLEgsC7pknqzLym
PiD7DupVrHRUQU++9MGh7ZeEIbBfV3URnel/GL+rDD2fTdC0G1fXutqsr9Qe
0kU8Lfwf0+ZZfj1U8mRyXCIRuuAWj77ZfuxvVCxYUULaCq+k/rdk2gB80K0b
ytbF35O4CXffvR04h2ehmQBHT1AlEohyayK/4KNfnD6pHtsr/kmsdn+02Km7
GnfbcrcDaIHD1uM+AIHN3DApvauaHUTp5mxzz8b4bLspsZc7I3VKvjpn12OZ
gYCZK227bLMI6Eh0lkVHFDYQoyu43w4QfD1uySojhCSR0mLYmWdnyktAXFJ7
BS3/YRRQvTKlh4KEM1jlMqj5yK/kC/aWls54+K3j7wftMIexYrj3h6iQDr2w
uDOebIrzGhEIYPI8rPIlv8ZwEnOMSg3FuqR5k9gcAZ8h0uD67pACRDXR+EKr
8UpAs4Coom8KZSgDi1/4g+1z1BGFB/GvSR/NYvrX+AHLxcFS15M19WprC0cI
5gbDwmbk1ybcknjiop0ZFuAX5tcxuhWkdktYRwmsotMZXrCvARXpWUCzHkjj
shhmVWzvjb+Zc6pFSWs3yOH2AAEOcII7Q3TZZBoBsJnqjnc7pDTFFv/3/OpY
dRmKT7ZdZNwW6MgsWO0hHkO7ZX8SOBVG51Ik9v/3wgiBVSndUMDgMXWltifp
TRH9ZYyyTK3wnvWDAndLD31O7Mfw+hoTEwkY9sjQaIiuvAhviFty2zOfMV3l
meoSWVoHaQ0Cmv6oPkCxrUbTbORu00JFg9Ci1uJxWnEfItF8NKg4Slsv88/5
/jhHQBteTYbxF42hezu/tBz/sW1F4Q+hzhnuQRsOAZuvDIbXjuHkMOzP1Lt9
oGAgkSuLrOj3RlVVXRMMGNxS+z7XuIx/QqkN4TvRyZrkmkM4ijP8TTH/LkTg
Gib6vwrSP7mu27lE4AzfmjHacjgDjeFp/2L/C1yRNgMaAWjtfkM5Y9/+e115
oLZtF4HSZjNRo42NuX6folpmf8yk2kGzVpizPPzPPAQeC50rhKTg6K+YAAku
AARbgXK0q+5u+GpZ5FKfekpyy5Zz3uJX+/xD73DpiTEl6NU6rtE1bMY3GkD+
v15vTF8Q01EgEIfmn+dsObu06Gzuzi6K6oi1rGZSfRZ+7af/jkiiHR/TIVbo
D/54SJ8lPT8MBw8aaU+Q1ObBad4nN0MNqDbNUxKuYGuUTAsgzxATNkPQviLt
ReM5C1bxZ3SbjBb/ujAGZNGsFF1H2XuJPiHlBqUzZ7gybGB7aRanNG3AbQaj
z99A6UeHYdoRnOZIvy/BiUzeISotTWhP2ONQhjsMXSWqJJVoGQJF0gVyzHMU
j1hSMi/101TovqhBV8r3lTpmX3DIqW8hunKLnkifIi7JOiKoUP3PuK0v2FhP
88wuDfNWchgaL9F6tmP/BuImqPCfKcCZ9enzjZk8y8M475HA33VfwOXaisd9
RnpZ5qYdF5vOFA6YHblIsLM/HCa2IdCqukpTXc2xV+GTNh+UPlhXyCBOb8QP
qjJuzU2grwI/Uu5/+0B6io547h3Y3AYh/Z6URsH3bPYOGoEC9tOn6aiYhYja
Vf+OqVj77IMU5FbHJtTATjqPNE3r7xUBgBMWkobG/fa3jPhM+hVRmxui1xPP
/62dJk6n490myaY14oTGXEIgAz1pz225Ppw8mPdVNp8up0+i2u+HZlEHtHoB
jpCQSrcIghT+68wjN82dNfOuo9lh9HnQrw3VCMCIjYV/OYTAroQ0DXmGrwG7
5mWETXuaOAmYC9mFeQKE3pZH7lFH3FgXM2IRUwDS8Vete9+jJxbo5kpmZp/W
un2xXXTWGYFpSUKNt4uxU80PN/zLH+jcFr3TedkxSnzJs1up4Ns9m1rm2RWU
KQRAOeyRJVQTQ4cIABOoYOINLCNP35XGWehGIZRwFPiq/tDCbMbMKj1Jaa1A
uWd1EVTf+njdAK40yxbv41C3IYWTlhyoKsXrikSUvYqNuyXnWRc7WLVWq+/i
utMQ8LPcJil7qJqhvYR+lbcVcOP5vhCugTM7MEWgEmNBWSQdhIiGqpvcLaEG
PRY0iff7zO8TWEavb4XidpsR/dg7t3+BP3Ct04Lp0EzHVIHIks5FQoUXksT5
1SKez69Jd0jxzIhQCAQpbocFnGv8XupfO6v+rvt8yhNh9rNW9NXymspRW/rW
Y3ZbPTpYT/Cfw1ZNMWbkkNXOR9L7dxDgNgQny1bpSTk0zvRyauzMe33k2ksV
VkmP3h5S+ibzJJ51VruXwyQPv/9jPeK9vYrwCnWiY9H6tgyXatMenXcqWCMm
1xFJ0VPfOu1dIDiOuXiObL23imroehtEVQw1OCL0jH3roLMeVAG/Ljl7e3Ru
4dhyTz6LRYu5N3hje8YRAxqRqxT59WrnlQWtlmLeBePIbEJ/gaFJ9hBf2fI2
G68e8jbH+alX2pSN5QjUz6pIWgNTsDMwZOT7bGWXWiOT5WhT+Jaa2r0/kCPR
i6L+tqJ3cTIlhdA8sI4irae/EmY4m58psF9oiMY1YfKN2dBZc7EhoUGdW95Y
wvBt19qkWcCre0EtObj8DarioO9q2kmwRFiOL3gF+3z1bg2M4lwGFeiziDU8
EZZuqYu6QP7xc52M/BdlR/VxT3THteUDfRfy8TJ1ewwLe+7BriBftJ48L0EJ
RUqKe1YsG5ApxlYXdLKdnHJjPeUbXGirlnQ9NNjlk5N2LC17ghfpE/wxSBgF
GimGgaowBvHoR56LZlCb2FKbulO0TKBk6oUpQH4+WuwlizOsT6cNPNCvx/Oe
WEp2pkK4+dXjrvia3MTPrDOEh5ETi1FTWZt7Wsg/NZ+1A74m1DiR47kqpVLR
NIBmMT2hAFL6FuX0qjdYi7R/0jw9XjttMDZGGxm4sWP9PHNuYGx0e333LY/c
Rfi2tG0Dob6mVhVAt1du/FanC1vGzm1eM/FlzMXe3PaEmmSoNmppCDctEDzT
o49JFOS63o1lvc19N72qPc2ZcL2eVLnHZxt6n6paFl3Uh0IhXaNNlg2PDPyD
C9DRMsRI0RMAwi5o8qdsC0UOo9HRrnTRXOBjPmt3Q1CEVKiDzguoUOBN5xVv
UnNT8aQBOKFohWsImTjJacZ6Bemb0suWqD+po1HRkHGFVLuqmBCCCBXBoAUH
RJGOOfPB3ciG1Wq+oSjD0Vz1udxrTYTAVTREwLSOs76sravUKzKxLxEtv1B1
77MZKuAxapsAiEavU86ZgmGXs4Sdg6+z6PDJGtBdnPDVjquEzUvcgcBhdDdC
VpRMLbHsAapz2Yg+Ese57rJS//NaDkrmOhfRhKdtE88A1PHO4MV5g2CSKf6a
MSZx38cU02ynmQla7M9foiRxeN4RLmx5tZ9DPExtJp11RBOcl62kZLLxFK7Y
WIN39TygmMwAPNFi7lP85Gln6+P0P8WqdrQTqO6PMvlII4z5jW/fv/UMW2Xa
7beLWW0wpzp9peAI2QYtrDBCghrfcbEnH/TY3Ns1LNqke2VMWlUDI335ImXm
5rM06nBGfx5KNFvrIaAyxRTtiF2Wxl7DQFjD8exaPsBvN7lJiOGPQcRegNYK
OsIWxFm8Vt40jK8YYsKsyDKMVIU9383tt3xAFwcScZwTLglNK1yHdVVsW0gy
lW0WhNQ7Q6/l7Hs8W10eyU5Ygyu7+rNbUJVBXrPauHYMsHz3ZrJrt6usGItQ
c3X5Nndw6neSSwbs5tBmw/drwD/oVvf/TSau7KqCVZL2ck5yf9NhyHqoZNXq
HrJjeR5PY/c36+AH+g1VA1uNzaP8w5VwGofXg7PNM8Fa/9Otr1jZVAh6hj/n
hQ5wNk0WboYUqT7/in0UNpq5DDvXXiSafHhT9vGuzkQyI8x1Lm9pX8R6tegG
Yr6vLKAx22qzvy1ZbJML+CSP9rYKLQD97gk5mBx43RF0Do/Ohfva5x+KQetC
aKQfm8wxVbHWrDd4EiIAN4qOd/sDCDdmsNyob1vWmzepSrRkaQtohAHvXL+3
HFqD3jUDUEmGSCC5AxyAkMOb20SB45CDdEp9I/MSKRlmnMsthgo6V2gaxq8i
JFFHPn49/4aaLQ3C/nOzqgAvqe1Y9BuiJZ16EZNoNNoKyB/lgSvpedFfUDIv
t2RK9Cm5CqmgYZezQsN3VSZxdcsxGVJDA/cF4cuX1giEn9OVTmYCyAzweMDj
//+Z2TgjoIxIVOtVzlTW6t/OKHK2nHvX9LloMOLSzYhUHLLL5rWtTRCA3so7
ZG94jhoCAk/Xwo1cpUPUAZ7ikA+7AViKhe8cNupFxD1BAmXALwVBt4tHoJz+
0lKazzGamvC9S6s5yuMKDqvrH/Q4yWckQPNV1W9Cdu0vcBa7P6J9XWLAZLgF
ZAegzjadJ5NPWkgPqZVG+iD8Os4k2D7K4LQgrzWR0qksQUwJYsiENvLeY6hU
VIGyoJShV3Qq1Iyx4svX7F1qOwN00hzliIrvcqT3NYdDs933cNMJKsm5mE/f
v7bBionhL4/MhTOkm+6kJ32L91tVbBxM+IwT4jIV5omcOxJFOSeoEtzyNon2
NoYZQKYoMvjFe/4SZ1GiftQo9mEXY7+A3bYs7Iv6nxnP70UDl3L/aVRWd7MA
Tj4PBRbaavoFLCy7OgGMgP/KAur0+CKu3pPCbkoMOM14LQuM61ZpnGEx0njc
nAogYu7rZRSVL30oOB6L7ikSujbwmLFDqoY+oVaSmqyHt0Rb9D6+8KRgXVzS
/9TtCXoQzaaGEXKu9a70aHOp6kd5LQ+CU8zxZglrleqpYpKQbSel6hof3MXa
q4ajcqtB/3oEzDBL6U3eLow69uDEqzGbZvINF7YRX8JazZ8zKvOEl33yUeL2
fn2yAtaOL3bKVGsdToZjVuuLmjDWpMvvvamkRsqOzWdH1e2I0bA9wx5EKrlG
VQAhmDxeHeUjU8GU7cPw1V6sQ3wDoOR24v87/uwxZmBT4vyhxDZl5lAbzkgO
GCNy5bFEtbsDz8x/jHUNMZ36lCT5/URKyr7PKdSBRiDQlG9MFch1AO6px8FA
Wa5Nxbd7S6ndz6ZKZDUVDhZTfnkiZjXe3c6JbuCp6vInXjgsU15MHNo//dQf
Kasvvo2uLsa16MomgxfJgmN93JqmAfSRWCT0QCNV1K1yBwirKo+92ffkrmut
qw8JQkxSfzyHktUiM7roOHNp8kSs3CCak/fpt6UxSC/+B4TKplFL5LaPW5gC
AfPRc3NnAB4odhz2wKkXADFBflJ2O2BU6E2eZVZvOd7uyOIW4Tdv22+goAVc
85ozsvxWocezjQDoKcQ5kYLSxH0xWtBBn1MYyR/Ifglt3r2F5mT6PIj27Ulr
Y8Vq7y6P7e1gnZVgB8vZhyIMavzGX0MmGx+t2OX133hWGEpLj3UzsMWaArE/
9b1/7HQtGOOOitXa2NfVaDb1sHJkL2ftvXO7ppvlcnpfLZ57nBDcb7XFzV6i
0P0WIm7YMJxOIi9ALX3dv7PXPXlLdhDPOCgpz1aTnkx0h7ezdKjRkhVQkpHs
AuThJVnZVemft0w/jUo0u6tn9jj72AfjVY9+THse7kilKhaO6tO91jG39mnp
TRCxEPK2SrT7iRPmKrirCEm5+iNM8IONBRl0gCkNAR9pnBV4phEqjpQilw2V
c3OHoi15dCqZpq15J/WHTEaElprt4yCjhAimRGo8tQJWppYR0h6BPyhQZ0BU
Btp+K9nqqoH6K9EkmcGr9eeN8HhsIl4IbfiJGOonrOEUz98XiyPHQhhZzpMh
BEI+mAezykmA4CBq1KVWNRqAkdvTXvOKwgbsBdpNUBP0hYN5/C0G03ZEcX+6
n5jbCJgiHjyRDN1UQAGtggsmt9e6WEQ4mvAO/o8IatvrJtUUe8N11X2JbWhg
iKHhTSyEHldJ3oZywlIP69p4TowpEz4jB/4WHtM2qrze+66rHPMyYFBTOfXL
3jfPCUQPRpEpctg+X1qXW4+THh/omOUSVNzJOhf+OrubIKBdkrfu04YWZj9m
ntEp7Q5TommWLDZ15AKAZIoWTovfuebKYv0JUguMogbbMuLMhEj9FmFMRwYR
xme4+/GUMJurC3xcjAuomk0XCg0BKte6s/h06DtRFCEjerhCZ5A1G9OAnqg5
XMfAIbfTdZBEAGNkb0Ie5AJejL0oqr3ohV47Wrq2EufSaQXMPgCnVaZkhGLz
C5fiGHqTDmCeDcbHMCvyMDJgZC5yel5EqJZJNpJ8BCt2rJy+Sv20h1YnNvT9
rS+fiSOMgl4ZWrxTPRNMoG51HEoc16ZbTbTvfdqc8G9zxASYkf9puE+Ts1ii
F2oU0a0z8IxCpK/dedU99kjz8l50xBL7O0H0KXeY2MJmkefx7WGqipTUPn+B
dQUVwiPctDi7egIqz3POBgQaYwtohEh3Y8Q0NQMN1k4i7SgVm3gzgTTMV63b
OQuLoqb48BL6LElCycI6e8H3Z9UO0C8hzzrMChTHn2PaXt6ij2yxZbuNBklh
ySPcBrGnwsXEAWIpiRsKjfgK87C/MwtROxh9Lq9XxZHKUBZFAzdCD3yaKuVN
5R3B/ob7l5Lo/qQwQ5oSLsOW/cdNCO4kWQnElPvVDrKtJ34AYOm7/QyZrdUl
vTJng6zLNWTfNGaFs3A4EJIsolxqlPvoiu/rD8vuOPcFRb1+y3FceiI/zqVl
AqDg+/Mc5A35fpv6IdU2RQpQgKvpbIpcEGfmwfVABJeuG9Km3fyvoFpKSBsp
tlH40j1ISlMawRGmFfnDUpPM0pjsn5AF5YPtIf1MS1dv2zw3yHJizD79n/Rn
pVj4VVm7bOMV4GPszJHJtOvxjNlqdgak9UmebfaZH//GFmG4h7ttwf0opmXu
eCpzxgaPxsa/mTt9qCRpnUK88d2aMNF1DLzaCYHTcM0xJnmEhJpVW/+CgRk4
ZprJXqi9gXH5CuEoJUYglPzwDE1e5jdL3n0WCfd91j7TiGDFLbrz0/gfeImu
TCHZbnkh2pz5t/6ds3kFwETFL0Vi12FHtKygDBpQtv6CkXW1b/xz0avQc2Ut
x2x07fONa2zWv1NXlNM/lRcZGlDg+yS68GA/91a3Y3PCbr4RzbZSSmIu5TM0
Xv7MiSkk9LUwqh80lgn5ch82uVsEUpEC7TerOuGxCQUnguh26xLgfd9HetWF
qmUckszJtD2z0XX2vV1UCqcTCpqIsU93IxBs11uA8R+B+1ktLpNjF0e8Dv1N
SoWS7Prc/K8cEdBS5VTZZWemEZeBXMQuwdZwt4wBP6mldaWUiUPjxjxotop8
eHTkvv78a7SzdrAHYt3KFgHN2pZuOv5PpPMwP7pD52tBynU/OARck501XBNK
0gTPP3wnF6aGkX69FnUBKXD1SPks+rl4cXn6P35Ie2KB4j25sITt3NTF7MEx
RFuc6/IbPldSbKRX7Egbe7wx+q3d40Poz0LDJXLDEp9ZlzvPM9g13yhACNcD
rTprkZsXcjnonrLwuR+EqFLGwfSLnwbXToRzF9Bhw+tgTvpzP0VwkKUTJenW
4lXDdkAB39rWiqb1Ih1NSL9bOZeGFQi0DFiuX+jjWJpEFFfr3HzeKOAmTILd
h4MU+sSaRwhDkYLoOoUjx660nAzSHi9I+XnShQwK4x6nz2niw5lA42DKrPE0
uVAIQtlcMugLFp8lkG4OLHxNmIjHNuuWOaoy+SZZ2zOe554a6IGVFjpsEYpq
IXtxZQVkJ5QjSNqlnKGbuF2HEtpAJzJWyfwNHDdWB2jQCSzDorwLn76LbaPi
K85Txwn8FVjACuHIJqma+NIwkGSbfQpuW9v/a4Hz++OF6X1rKJYhrvt6S+6e
7aAKuskw1aE+diQkdkCJ250xbqX4TW1gxLflrbysvROqL/xkq28f75wQ8PRX
bP4WWgnI1WIoDO2ebz7Qby9EcQS7ZccnY6J+Tyu7JlFA0gPCHxqDTHBbTUw5
JhNq5D0EBoRa/3hTqfyCN1EUIBNbwL1HcqR97iJykmFytz1bOkiszyAEWw6H
9MKT7pBJ65ql2pQqquHDspmHHyCSdr/3E6klYJOGFnNbCzYpIktkdhDV8Fl4
2o9KIb0aVThRXUcrX3poVbz3e4CnP5AN1+TKLn7vQDoiyAfbrHm/0/qM/rw1
DW8dtnKcE9AU5wTz86bVKwXChK2JyalUP7m7BkHY2qdHT2tJO3oXq2jvROSm
FpDi9gTsBiEmouiwYSVvvuXn80+sWctimAmjsxII4cCXVFMczm8n+mb72rpH
BDeUWFl0rjDKS4uXVg1LB9oMQCyihGxt1rDxj7UoK7ZPYsLB71PLNKgLP7NK
8Hdsl2FSTNPLSBF+KRpS97ihOuEM+d6f0fCFPoqk+r3GXZVIpt8jSsHoUHdG
o/2b3TNsgZYi+xvgZ8JsB1Dj8/eFUac8zMW1TGreAcpMrPY12qlaQjJ2gezq
Y0WQ752abc7e84aWCf9o61htjRWW1OsQKCcCq6pSIrVwGwrgxc5ARDuCcKiM
FyZV+kI7UqCRJjflIQynhidAW0UQ99GVvMAVThJKJH5H4naVVwu4e3cxLk1T
nVRvQceiiXL/oPXh2HeBsppz69sVF7qriOwI02Wxxc5JyWmNMaSs2SyW04u8
el4ywGRKvljbnFNOqQoMy7h9q3ftEQUEJZRsZZROhJHHyYRLxYGH7v0XD0KL
i5TS3+4CJBL8gyD2tKoLesM7U7iyD9yWarMcO1qm61sTVk4dazQYfrMzd68p
b+iqa1oPYPeKq+Xz1BLl5unikf3hBYnY5E2gcvFTEePjcUFjDMnxTJ4mA4/z
L+MDwNdRAkRDYQhPJP4FDNzPXHvcBW7jDIXQDyxJpHR3fEtWycAAAqylMzw5
/sFkqj0UU9l3lyb0xZr+cXlxn+GDsj7NdUsxsq5cLPE2J7nIJJgzIh/cXZfn
Uwb0f8R7UGoOspAV6gCj+sZ7uH77xJcUecG8PVJtd7hMlSNBuHAIXWAA6tEQ
JBA9zGdqavCKOaRZ/vliq1Jy1VJZyq2xYSQLyEUBnqbfE8xHwgYa0/JqhXKa
wnPkLoNhBRudp5RxES55KnYg11zZeiOor/ML8gGtJw48tKsEfejZWPGagUW6
/Uxl7+8baSuUcc2mCtWeifac6Y0TEbYEfA4/Eg/vC5x3Hjfr1A3XaBCIDqek
PrE21Sp1z+i17k5u93XOA/PVeTOG+XQ0eN+xpQrz8WFfkhJ8e4/V37d+xEkA
1TCIXllGNQT8VLCoU3KmhF5o1IQJGQexrVxAminxPK246A3p2ORQgNif8WlY
7INFMTcsLXzzEvEKFlBeUtQENYkIi1l0rO5LgCESA4ZqRyoi5Lp5e76+BH2Q
lQ4Bz/fTb7QcFZjNip9NCaCo9+a+YhhkQ7eqjfGXMISC1vnBi9iCcq2B5WQH
Gmsz++/Ij/Kgf6+eHGTpcgAA2ijkJwjRgQtiqKWyUKPlhggwTVY5Yc+aeZ7t
AWwdSWYWYwOLsS27B3JUcMuTThkPdpFWx+rTHP8FiDz1h6XWzUOgCZodhBr1
OeI9KSS/gZOSqC3khgNHMXYRvhlxaUpOn9KUPVOuolLfcIo762RhlZOM3al6
1D18vY68HXB6Ym3FQKLoAQ9+RLorZ6jCtTVP5aT1u2hyUkKGqyrRyfjmcgqY
uyUhmkmpKsn4GwzdPuKxvVe+hQBg9f5Tmb//PokiKtoqgcqxUO7Y7++if2b8
4OozLwDw3kuu78aQsSaZnvVKN/WITNM5X+vMGSTJVjILiS6hXJRl2Krdh8N6
P1/AybUUP/6UdfgNpOGJlH8GBcT233pPMkKuTS9l4ruB/q62JxLMAY37ux0l
1Xcp9wzDecvc+vuonDA80GRiffW5UkK/wToKdbfFcp3YexGcTVDYsSqOOXgl
Llf702aumpQL3C5Ss+pJvJE0T0zV/4qQdN6/ZU5tqqXDMvezpbSITjRUPMKa
qwpZb+LH7wwP9AWGgTwCWZerJs8XBBP35HqX+5oE2KvJiTv1vLM1V937y7Fj
s+06BeQT0Tb6H+UTVrdDFu4t1oph/glGSCW47o0ygv3MNf3fanO68TETiLZd
63dEElNouOMle33uwVx0rg1x6orqaVaidhtfp3ohiqSJPP7Cp1LNL7AOQvV/
ER1fa3l5HKBx6DI4Ah+J5KC0o+I/CovvPIopkTWij5YwP9Z6dOSHr3F28tTX
KeK1QKVYwOB5y6Jh1fmuyghVwR9WitehBWmLKCvoWbP6ii8RDdKX7/Xkvxu6
ZGwVj4cxD2h7CLoFO2qRVkeWAS3Tm7f1nYUEPSdX2CVtzXFT85yqd+XvcGGs
hUSUxNNZ3dfF13fqqJWzRZv/4lYQStb0R/Wbq9F8fmtRgtXZ0IfRSWtFFksI
XnbdeUNLAeT08Qat89db6/s7kOZrv7SvmWEsKiSNx7pZR+8p2cpq5RqyjRxC
h1cj31bSSbr2Q//tsAVamaC1NW9eepab1OjIYdXiKZsFi67i3M8Cu2s3Fxfm
7zAD2nBwNLmdF2UMazkJ+cRAe6HXeewjm5TouTJvHolbyfee/KvXqDasVia3
6m80dlZDAopPMBOzE6EAMxR/ktTonLB+rHFigSWV+IXrWftUdaZirE9sSxWi
EbVPp4/R4jSYgkgBqA0eXxPc3XIQjtzDqpfJdhecSYrKdtZ3rDkPZ9jqyv8Y
IRSs5ZA0l//78w6poxA/GN3br1pwXOdyFvugNpF6KibYKT28ENCC9AS/LG39
/TCOqb1oChDxko2znBt8ynsDtGXXnHQnO9avxranEJWMdGyiGbhqfaHEaUIy
gX9nMSCj9QoT2HTNFEhGuMlqPZ+tYfZTn2Cf4zlD9ey5LhnQydjqiGe8nJVy
j+aZ6jskDg4s+VCuF2r93PY17eLrL7UXmYrKL0iXthWtWlb2Qksa8oX1glFT
y5yzE0TkObmJ2dwtumndLHuEEnIsu/2jzXY4DX2+p7+biN/3O392ciwExhFb
gDuulSulpqSWTuW4/rDHZnu6cJ6KwGkMiiNq/Y2RkwX8CTGjgpXnq0BcoIGE
XSyZgg+Hm+tFKGILfZVj5tUtNXIHp9srrfndv2LwkEOi7/U4eIdAZxvkEJ9v
NhXXk2CUngVX6tZ0seGED47TXJgSx2GMnarYS6RukQ7VmZ1aKo43iXxDJmJW
2jiwSbxLrnxf9zP+Lj4gHwCkARjurnWVPjnbX1mV9XGZWrtyFfevZQO1OXd7
lNagVPJl9EeR9GpneqIgVYP9g0nZ99cngqLnGT5nyM4ugQ4KnsNMTsmkR8N1
ZTGkpfNhiHmSn37qXiXqO6dBYzDVB2rlq/pXwdpi5vfZXYgNHACQpSqsVsaM
NtYAIjrTPqLiEQE/R1/8oUsjoMlSbH8Y+a1vhCrs/o851FnhqrQAN07VHExl
UxhAQMsgtl6qScGSW6MWcHbSR5XG16KLQwDMuNwMAqX7J/VwOpKG9N7yhaZO
Rd/QrXLImt6Sf0/obtgfvPt/yYuKvSegv5FOtcBuBJOvnrmwnbAepZdfJ42J
qrc0Baaob5/ykSAMDW58IFGUaoV5qd81uUga4lU5YIYrUJ+1O2tETTJA4eNb
dXGVu4qnbseEPYwsRyrXW+/6fqbwDhkHcSQQVflNB6xWXKYT7pZZMzkDL3Ca
ZIyFzl/rVKMCBcplh654cncenZZ5GhqWZDt4QGIC6CwkhCy5t3vdkOOwLqXl
0WLrN0q2svQy9Ycbi1a4rmSBIt61n2p94Fep/bUR6lBABwAX3cu4bjyOc20C
+3QOrK7J93WskOXBUYz4xFncrSWBSqirD+lU9uNlg0WBPHFFjjwKuplD74A7
oPvxC6HYOz0pbyQVNSj3pIfaukBwQvPldWg0uCwghVlwaNWBlf6y+lM2sJm9
X91axl8qCd8tEgNjOfFUKdxG4I2/2mFGOXvjSGZvWvg4+hrK3if0TUGI1zmc
vW4YQbY+0sl0CjTVbMTm27q0rpXi6XdAiJ6B1ljF3OTRCpXBWTsT+/LK7vkr
bKQ17FVoD2PRi8n/V334sTihG30MmO/ytWFtp+mgcvHQeyr8iZdz2L+qOvYS
hue5orGtu3qzrPjqK2XRt5RYHLMJhe4nOZGtaJ/Jk/j5n3ue+HycdUnCY3Dq
XXESpzx+lxWxJ8S7HVQY62YoSWXYOb8Uo5Y6UnbXDAslr1//d3ZCschXV6bc
pNx4/I8HOFDJqWr/bBunLYFwRlyn4JGhXI4lvAVUiTrXZe8TpnEPcp3hGXyi
VLS5Jzj6wPA6dFF5BEAUDaVe1H4RkRLG1jLg6EuZ71bsnjgW442BcB0cpyi8
bkOpppAqelK0cJ/8YYBy/9R+TVrjcujULyK49VQQtKxTuwoOc3pwDaBDJ2dM
KtgouDZfU1s/Cdv6YiW3BBtbEAkdysHvtkAIkh6GBo3cU9yz4lJYMaMDnC/J
1QCyrYR++YJzmbaWiHJC4zBwG6W3VUDhQuLWg2FIRKthmcOIGmDOhW1u735D
IYgb3aYghX86Vts5nCDyM490nDahXSWvv/49Zq/TLeKh2ziVbp3CSo2BIqmH
JQApXsURg1jlLsWqfYXgRwGleHjCRiM0Ef0QHUcJaxkCYrsck00TT+W28ssE
dU/YfN9kQGMFLCvslHPgd1fjCe2rMQzRX8uYLaZPoL1rCGW6zduBgUVJGdjn
6RCmpejukiJx9aW22b7zrgA8nlC7cijDxXr5LuGexWmyoMTcbg9Co/V8b4Kx
2LIc9QdMFEd4AThjSyYtHuFBXZ2T0gI5WytlWI/bwVksQgstGJuKk0lIu0rA
GvrFxAPXlDRWUzkIzAyYuLCfP6vXHLwNxgm0CFDLfMtBu/uNZHwYPvUBPyQz
iC9Fg51KzxaH4fXDMVQ6oVSjD6fBan8z8Jbp9mM4eVZJyPo5L6bRj0iTpFTx
2EC1EAlp5ynCcv1mbX1OuTCDeoUkh37gaOw8u3efQ5SHcEi6a/u4N36aHLwL
azqI3IdkxNSJcK4mYVUmyO0u4jBBdX0uHaCwJiTxjFzt0DMF7czn9J0p/38o
+CIKhTofRDxCTuqmHVz4CQYoUZrS+tdkEtYOnCV9ugu+SvrwovNx7pP8pCCi
L7PyDj8DAaxmVOzjQg9rg3wr9cFxYgYuv7il85NHF2d02lYq96gmyfXPzTNP
2J5+gyGyn+hQYr4ivFpjGxiG8Sol7RnYv7hKH8rQCQDZmUEHto9th8b6bHN2
MlXTa6emGglIbez20Ued9XDgAYdbrnGDM6pze5J5iHUeemf5hN+7Y6TeVH3I
kTmLmIKsyHYEdOB4dJOVi5ToduNcBXqpXERO66yceNNrzwSeWibIzHAtbl9o
7Wam91414hAjDtEHU5yqvGg8I/Ulv382fXtG15qY/7LNQsABJnRuGn6qskE/
R+g+nYRCgOHfFHY05FLEmlmmvyYYfCU8i3vnqdZe0bQILCRTR05OYWLSeR0O
czPtuUk1SVYM205GFpPKNuZo+jsfioHDjUY6I30NzAo7dp2cSjzLTJjxTRxE
L4g+GHrfYvdjhysM2e3n6WWf1rytqThs8ljkuIiR54lUlgIYfacE5hfTigdy
cektnFEvKEqig6nc0l8eN6II47jB2ZxbfPPgRdO1MDSWjcDsOFcPS7LX2Kh6
O8TV9I7w3iQifOeV3ND0no+sOrAd/3azG7fr6kNa+A/Y9Rezig7YnkBypGxV
FSfGR6dc8mCsPCWMshoL6BLjE1EQ957daubRoKlmDDSgp9EGfS2IDbpdzQJM
DLiTuL9BtO/R7Ml1zsRFG6QQXBREGBZHdEBrK5uojD3IGjEVXKWV4oocIzDq
EvRXJySX8cNet2Fsg9r4O5ucLyP0UW36pcqizyGTs5eNIRGdGMj0HmdYgm3J
lINLhsvD2Bmi8vW/uqetRlaENI0c6iZ19dDxjOnMNy9McxcEOPiU5hlXz7Zt
i8JFoDF5UOpBNwMEzceueTGwucJu7gcRdoOUjR4DWnRgofZRG1UorwTlXt82
zpb6pcTFkRAGy82DnELUE5tf81nFcCxgL1Hs4MUvgTuT/0uMfkrEdI6hABSy
nVkU1fJ/zkE7txYC8XX2p45U8GRZFosGvfC9ISD1IIP21NMdcaVkhiMktxhD
lhHMDBWghkVsp2oPV5b5JJuGtkLoF7RUSCn96qJbFwpAiRTIkretf0PMatfU
W+Xy0LxJK4vGqttLOcDE/3vHqEs5iH/FV9B8K3hJFGO+VSqdS5y1WKVVcIIH
eQs3bdAxRNb5lws50Es9R/iIJq1n3fz79EikBsMrf/ziLAFg4h4ZcoCl+9ES
3zMO6v6D9n8v6SyrFLzgdbZlqlHxPfUKx00wiOa8Sfbm9GDqSFwPjfHNxZLx
lR8mFGQeYz34aiiyjtL/hpd3EbeuD+J7TivF8g0pJpCj1zs0SHLNpXxBmjxc
jekynvXPAroCBoMdb2kPfJWQ7fQzwwjIxqCItzOZKEPkORU+UTpiPvb6PtHj
y7j2nKhfMQxnbP3mc5i4H31ASLzydj4qD8HkHA8AG7jZ7BmemQYwJaAazEXp
koTl2MyWSVKJcA9AQqpACPhNKrQ6B6GhV4ZruTmM8wpPFOs8eEN5oRqK/Bct
gCLiNkfD3NVrU1GQTUE0ImJMYHSRt7yabkKD2D35/AiwqFcKkaww2yvBE5t7
8QuS3653gkKj7VrYy5szOnzjxwYe9Oqj63DSbrBIVnnId01msB0hAdx7O6qm
6x5YjJAoV6+M94pYon6cZXrlYuH7g/cK/bNGuejJ9/p++2Qr9MFKJRr86U4q
lwmI/b9xdr9lxKq3pr2tyQG3HtzUT5jGGJ4cyyFUudjZoSrz6R7ncfw+QYGG
lehwBZTJe0VefPGvqVs+AJgYmCOSE4ZMN+0MZMgazOLSZJYgoKXJHETA/erf
gk2lrv7HQ5HYggorVF/z1kgMCJ/A+++gi/sNwgDb44zseSgnlmvj+JRwcaHS
7JKyUTnIPhkOi6K1F/2u31vYHa9kOj4dq2EHlReXUVYJ8km/LT0Wh/b8yL3I
Qc/O+JbSl2/afeOo1/Q4EhSgCa81oKwHJb7MGp6E6kvy6yBJKmdiGGIuql6W
xDRD/pGOODCDttHcueE34+Ri9oWTnwl2tT9CenY3J88kC4FkvjHjWMCMWOA6
nUJquSDmFem9eIJPJj0+OSDWVo4h5m0qKjiSC9snQHWNgspZYJw9XWQ9TQK7
lQcBibs+Mq1BUqG3psdePlqtagx0LPdKhpNbg5C7l4SHnICkeE6Ox43W+Kfh
0lglbkOMUZ2BGRWpQjgOulT/PCMhZRksuk0h0B4aDCu5eG2b3epbt5+AODUz
RbBkn5TBt6nxaQrdNAZTCXP02XjKgJGidL7lH/K4UIrjLWUqTnnXEB8iooeb
PGX59bZ2DRLmecma/CYtfE8C4TJuuJE7YST0FvDGosboWYx8QNvLWGLIVGkB
KLr7eoopyfpBMSN9AkC5Ca7fg56v2BGUHb7l3cM1JIvX3uVf+O8ez81wELDR
MktLEDfKRwqe4bxZSz+j3Q3kwZwbCYvK/kUn7xUrlXKumCmvTQyam3c4p5xN
gp5/1/KNeLngFHVZRi59OLh4wasQHh8Zr02+ExHp+d113lAvWVTeHc1eKa6b
bLveval3q0VyJe+1S9FzgXtZrDDx1hQlRQuCHgpDVddxE45B6BJkUvLec2rD
h261pN5xsQtET5/Lh8gltqB9W5EQ09zFxB+0wBFG9YjO4y2Sq6I97OScXs4d
oJ8t4egaCVVavnIy0o4D9gz35a2YnLIMXC8wsnLG3pPFWG3FBSVjFkdeZNEG
ENIpsXu8dNGpbD64AKkbgzEaGOMiDilJwIURa4dlnCssjc6Kg+QiDRdbj8Pe
z51D4ffpThWkFGn4QZvUR5i+jC8BzrbCBRIE/HxDluCUjnNIDpQP5cxPkAy1
68XFu9LR62fT7VLHW3I9rozwcK6O91QZ8kSobjRpjWffDTkgfVwNjnE4Fzpk
ekyKMoEHP1uV0WkYNIGMHb9QjBFEqf/EpVsK7PGdZ19rhFWTiXRtzvpeLp8/
OFqz7FT4bXBuFi5Vq9r4UwCQ0kv0qmiOtUr712Mt9zV6n9wt8njfnO4bvq4p
F2NscLxF1MPDzD43XeOH8nUY8tQNQR90xLkZaynINbZXLFP46zkyd5tSGjvK
HqsCIvcsYsCa6oI7kho68/z8L6nCYnTNH2X5Jxx6lvkD+9h6ML9eWutmvoU5
9//hq/d26rZiB6Xmg9duPskkmKSbH6c50g1jiSblX6+t3I001hVaNjI8eEOI
OEMEP614LOREW4ftEQ8awL5dUQHpZQ5kTcr4L/i7MvtBgP3nMQlytcx8wzNa
ofxVL8xdVLA76mw7tXLyOU7/uIUxTPaIIrN5QSsawqMGy1Dv8FTvmmftf2oE
lkiavDzGX7a1LQSb4qvebOa2qfPPcrgbacNWq5PHU/fTlK787NiVMyco6xfl
liS+m2pSBAwfK3pdZcG33mjfLdTT8fcug1eIoh+yocLSVzha14btZH4bST8G
24DQGsdTShJgSys3bkgDV7Hls0Mql/ri5OJlLepdPP/1FL0ztkpXxYzO03XO
dyhOhnb79T8k4M9qxPClcjJmREo8QzTjLkhsn/OJG3n3kHhCxQCsPE4jAWeQ
ljcHEMr8WRsKTwPboUBcLevZduUr+DA/mEaEc9HzKxkIcVJe0fZGESBxT687
oAe4tYEZ4gKw9rn3MMk5+isdNNXh26kYNEqzDHeQo2bATXJ3a7yne2vamN0o
ke3P1p7JDPgtQMggUAV+wGXtveWLOkr8/nvzuZiwuboxJ2ZWgZdsueyv8Hm7
Bs4+eg7ppKEDrY1Sg9QIUl8hwrowJFe/WmrjJEghJUiPFkZzwoX0KwsQEK7T
QScdRq8nA/BEfQNe5NTRO6eiWvyr9Vq/bajRvCKofA6p6lmnHjhEOPr2QB4R
yJ5JFvqQeDFVH7mk4Ma3RsWcUat+wlKxvgJQVNlsXsuQA3r0g+oi/FcsMTj7
GsuzHU7PAh3UUnkMaUyiV9kzTUF4x0F2KnL5ejMkzMLEZeH6nk6qbLYmggO6
B5jUmObpafzQIJuh1otEAhy81fhV6x8BiYRQJzg7HhHuzWW4JGX6+vzmvss3
Fc6+G3Ijxmq/0+7fZqiQdvB501FX1Am4KozTtSeLRAYrhm3db2gMPOJRXYMV
zyK25f3H3nYDv8GlSR/YA+e9QIGZ5O2T6UgIQbEbRnvU5f1JLawoX0MMeGkY
h3OH2ZNrnvhXBgPLKecdaG30IDWCw2mRDN89QlzAXiuuNmeilOukBViv2hyh
cMlXKusWEb8fDrOKS1q/YO+X5LmltCT5vVydgcjcJ4uxs0Ofd85Wv9Y642hJ
xh+G+/xccibHGNJNbEgE1l7qXp3kwhkWDhFtrqB3aO8SzznbAfef68PCS4p9
nnAAkt1iVSAwZKqv8jtQBAMCt5LrKBpSNtHVGS6fYpyxol8Mvo5SCkzIrVmQ
lWy5Fj/qUU3o7Y8uW9FX50469Jyx20CRnsTi264RYM0i5LZd/B96RLPouHfp
F2zG5dSmh8lcxsgstLj7ALwo248EzKX++jasNlL8kRi72LM9uNqK7BNGRcHt
0vOKsC5B1d8ILG5/2UOj8K4I9GIN7+gNoi8VY0tCdzeYl54UnbIwQ4havybz
jJEmxw5doVKEUxBpfjlTJ3Ps0aU6gem9M8frimcwZjJJEe7ABEnmBWyS4KXn
YD4gTTivlUEaEwOzXLsrO4IRECc4IDDjWYGM8QciwS393r+z5cY2uJBPMRAT
MzEUMKa9U/kvInJ6pqqW8gciS+2aWqltBMuexTOjo/ujRm81XN2EYrlWtVl1
dsC8HYHdpZq1AvamAsd7MlCJsNNXQtvP+0dw6J74c2mr6YTEuq7Fe+/v/xyZ
/TXvgbS5NoD/Js0eYjpX+qVhnTNZOOCWqN8jHigL4lLWRsywCMG6/FPS8kaI
kgG13iIBD+RmhDAtEqxVe+AiScib9O71WYa8IT6vd4OFQC4R5KAcCKlbFhXo
QndxC8z8gX/PTw642nzStXQ6/h2aM4xEc3qYlpeib6JkNpnIZmP8dpQM14XG
/QYihu+rY6U8Y2HxNPMw0tRRgecgyj/Dj8ee71bnkz82pCx/wpVHAzCXg3O3
QeWpXWH4QESb7qIy2ObzM+sKbo+gEGE3HJt1RozU5v/bsOxXM0MxXhgwKXZs
U3xBc0Gpf3VV76sRw5lfu45v2ryVUEwTcdvduBYsO+NeSVcB77Hmw3tSuP7+
gX5c3hO4/JevS8ns1fYpemsKk/nIJ3XwioGVhGrZzWRRXbU2OfKyOcB1BkjR
VmMourrtaKbKNYNMJ7dCSKwhs9KmAu1BZjIHYaEd3h14bQjxHk8nLnCMYpAh
lCgNKq6TD/okrsHWHj64IvX5+R0zeXVq5n6f9FMWu8NeO2xiBAryCs9sH42J
7gMZELWtcB6+3sPjupugkqXZw7frDo6H9Ubqw0flixxnXgTYuMsWvkVbl1/z
tTz+ScatOJq/qaE8sL8onf9e0qmRtUfYpW3x/PLP1fsfuPYD9dWQFbgJnatr
B8mOkVDdHa7O3Yoc1rUfzKryvLwXfwFgDWjfWWSSZBFyoTqRVcs5yjLZB26n
obkGWQhc/LuQff+dmkh0pibRj+tcU6bzCItAkfv6Uln1/fyPxtCyNqBvvv3z
hsJXkRt8apy5nqH2aMwpMpM/1wp/nDk18yeyASNZiftma4DzTia1iuUvXjgi
ikSQT0sezb8nTuXiky7kiRF0wX3Vk/i5CdjlyxBh6ff3ux4XA5hyesGv0Yny
HqrMMHjCVg4HcIRyVlLoi0P3YIwOP8+5aizKJcMGN92h7gMKumWW+9L35iwo
jVtbyiwlg2Y5Xk8Eytd4kNlsO9oOgZK1RY31GIENnAvhvYkHYBXO5T9h5Y3q
zW2Zsnwrkxq1mALTn/3dC7Kpym4usVvke3cwlw1xtrIf0aJ+vfUPrbkXdAvx
2cNfU/0SAS+zXHiDNMKa4lGJZW7V2bVRqY+7RRoRJ6kOzdbXHwHRMtjkHqHH
mhEZk4N+zrSGe9xyXaA4Ji28yLdTAliDR0BzPJ3dATHGFrkIaUD/Ahub675y
3asX2xABbMAvfU7CWCk0pLoewFegnPgz/AhTBG8Ac3ApZWCcnNmIZObSmKHn
pdw61xRLzca2TJNwJLTLtzYh8QjHcPX1UryrpbMj5SqWo2yFC7znskj1vAPw
WK4AoNCRRXbhFsiXZDB+SKkzrXYM0bShhJzdDQvYYqORz1Er7mLiW/Nn07Ai
1PgND3RJHV18A0VuCWGz6I1sBqCkLvxqii6IcJR5fYWukpJjvWUV8uorr6hb
95MTbbFToB0ulIcwjTAJw/2nFzebaxkzVRwgZhE3vPNviF5WmEWEYdHTwPC9
9yWHwlHQks1HjheM4GvNm7BkNtKI1u251ehk/whUzFRnjCUa8zi4EPIdSM5W
y1dUtKlnz1vthzs2NMXDAXXgqpVyhVGya9KHlwfH9Lp3UvK2gkaB6J/XpOew
yDgvU0tASqxAK1whFcMCHs1p3ohoSFNfgrK6nHW3gWHR3Xz9I0wpKV3ibEyY
XwUssYVljwW9BiHL0be2OTAyTGigjlvGanvhpQc3NU8bkmQuDEDslhK8mhbg
j7gAsEkGdzTwjiXU/7EGb/18lWoBL6ipyPNJDLvolfvBNplrLQAJfCsRSQUF
oG2AGrymHCpGfkdrp4086e0dg1hdQL/0lriI+3Bvb2FsRk08kFr+NTcRRn7F
3VyktGmpn1ZUcBc62f0yiGNY9C88r2/bhl6DU0V7V2EncTuZxXtbjoZJN1vF
xX0x3rN+VoFCRs7/PYuCpr2okZXhEJKUdbMSS8VPbMsfovdMzMuNs89Mfjyk
oTpZdWjbol2VMPsY1GI3WDyys01pHgiQrTD0pzbxF+tVYCymr3sTbI7bGJ+U
vocj/AmIIa9mqIpAtg9N1rPiIt2vza5ss5hvTE0RWpRUfZMnQb/56wF689QB
sveqCr8TLE3CBhp625ETqvYRDtKKuD9fHadIiR3PCJVPcZbz1AvtophxTTHN
//wHcd+/eFZ15LqYcWHWo9X/88GwzhwClhInBCZ7f/meN5w1Sskw9wyW0HCC
E120IWTkJsNAmDPSxFvQGYtjY+S3kO8xBraNs712DK2Chp+M2zar+0jGyfA+
/dbgmrlqFIwQPOWn4YOUtLTakpRIi7VO24QzfSVxgjYcgYU2aqt1/BUL6poe
I2WfZKz2CHuciyWg4JEBPdbWdPvo2E1cpFSeOZ1tkLHgdDpgXZw7SB2zJjgU
1FHMkekG98DNhhyI4ekX0lDgoh9SQrFjSb9/46oq3TokfbUfLh7h/Qu89j1d
aS/bkU/WUDPbXnP4HXdKRz2NXRGKQhyUN6bVr4uwka2OB/Tnpl6GWiikwDrb
ovrIm8fFvwe1DvM1Q+aX9zhxCfcgRVSsUFRgBV24Jon9c4f5r69OvIc+rOcc
MghvX5jR7ffKiKpsnnT9K9TTB26nbZkThONPwc0aHnnfyqqO71k0nCLWhQ2o
HFDLgjtBfvGawF04qOFO6VSpRjtFCL0FkBNzazwaq5K7RNOP5HHMdsgOtDGa
hIQctc2uP+T5i16+PiHnRwtrnadwj410XDlSbB1VZzRFDb+Lz/uC/5NLYD/k
WDUjjk8SDsIceShdZuYvELvOoCl3sRU5PVZmgegWZILLfctn6HpSF3G16YPl
mfaF/5BKXxyUnfs4FOGGMvPZYVVqyaA5nDc1WO2+vQjTxklM55voyowrUrTF
+8QCeYmh0QCu0jEnL8vUrvjrJNQZsu7JGQCZNyPA+/1hbY8/caFWvri3Wyo3
xCpwa905AVkOiDg5w5YFyKqXwOROikRDaM21Uh435B6htKjrgQM3KW09CDkx
H2rscPG51jkkfYoHnJ/FuKqrhL9x+/dS9FaqMih0Xy2KNz62BKkNI2YuBFQ6
gEIM8eG+fKbJk9uqPTsgcoRLVjzj3A5rB8Dcg+WoYoEHPQJjhdXTNb9RzFHc
3D7Zey/iCt/sz3nljaOtMbnupqC3rfF7FppY/kdqoZpzpm4bLebkET9AT+KE
eMOhsYqtk7qCf0aLxXE/Zx4HVcZV4n8vraQfiBwUB3OgOvWbRYnYGS6z/w8v
g+9AXAHd736ijuKGNDUXWEcgmR1qGLo0hnVoxFD4/NMC2HLyS3ZiyL1uFy+N
MAcS5jM0o+wl0w5dh5CB6UqoxjPXIvfVb3ybjOdPvOjGnlbde0brbMbVHGwq
Gogxwbjv2qCPY8pehBR0Ozq3gttiuDS9k0fwXuMxVWOOHYBYHMiGbOCl76U9
+6Yjdp6IfBdlsQNO7Gz9jTOQDNQb6e9UhqoTIzNcy+UygJoT1czWWswycyU2
67Umvhqul7k+4mOTvIFsg53PDtnrqW8H3Ty4g23FbvUzYaptdfhIvniBmv/i
tsoMDYWKgpB845AA5qfG8LyJrhEcQOaw5Iht2rZCrE1qL9qcwf10Go+SExoi
InaoXaLyoopgHE9F+qHOggBgLk9NbXYwDOm+agi2JFb5reGFkAaDfOCbFKgS
of69cuGAwfqpTT00dSv1afrrQ2kvaTkBRa/w7ONjji2VB2X70+2KHVakMxm2
9XwUee33rxTs8k465dKBCtefdXDSFGiV2Rq162RcXgoey0hUhP3JxsCfdqeY
Rebpe6dX9F2ijtINrfMIND9QLY83+iomCkwmZlxZQOgJ7aFcq6awiciyBaaZ
fWhB3SW7AUftkFOvj5iRhgMdwXehwsvXVksbD53Qyg6+rBytKzOKBT7jAnq9
RPlh7GC6NZh8HX2Ewv7NKlF06QKvm3mSlJ96wMDOBY8BJvEGtp09UfXR2Sy2
rdIU2UydqQaK7gg9an+a7CeULAHjR0XunNkjY+NI6Z7ofYaFy0GyEUJqHSul
0EeRLnRFTGgPG8mwVEgN+ecXFZHPt74TFWH/oFdeefCgFhr2zUNeSOfWX56R
yCY44fMLqQRgLyl2ETM89v7+hE0qcXsySmcs8gBpe9ItxRlcMx83EEUWSNlg
+IT2zHBVc14MyomtiH+/4g3mjzCNVHkaAzeUXw+Hw/pZshQq0gKyTCsVUuu1
83DWrV7L6XMaJfcu74nMQW1+WO7yoaWxqIHIjVfDRsmDimhA91D3BpT9e+07
km+Bxf2mrZWxQB10YB8dfsYKAWC7mV63sezl40SXUZ8FyRpee9Y7nmhxPVW6
bxMgScdfZ12FDGJNxj+s737JVr5T6LWPaJm5+pAbxKCe+T+ZeZ3PWQKgDwW9
lMISklxMhqhaTALE6SZLs+d9AsC3hFniMvwFqFzt0qlvNINVrBbrfLgPYGs3
a5zltmlXXwGbDuMBnOYSARGAkHocK+g8Z/7A1o8fRikEQfBDK37kL0MiBIiS
EHK9Ysb54+lTkB6W3m49jycl44NMpzS9Z8xFWrjf+FIjXVafu48wc3cfgpQC
nKmHofy8wOZJPryRMx7MLkuE4hX9etb3bYXtYsd8ROfaNQ+y4BY2txbC5b98
MwCztwp637RYM0eA5MfXmLpIhlxsaEdv5d7vxcGBygAIpbzutwDpAZLnhefb
D1hmevVB/tAsHvjSyUx0uFoC5yoYdzQYqPhg4PJ1lqBdyl0acIu2Ar0c2Zst
xA3huFLSB1xiAJgVg8NW11/KVzlsSmvmsnt+eVwB7HdzK80GOF+bkv9hA72z
yKarhhf15NTvt2aK3He/VzJvHbsCAsIs5CawiCRC4IBMT75PO7+V+RC4gxUy
RYVptGa/L9+5U2UZIYdal1rJ0cqc28cQuDYyXeq+COrMhkLoBOwuzeBhZIfL
uUWopTob/teNdCurIvJMQqk1Nie8s41waPMuzohTGe6BYKogSIyWaVDEbqrp
aKRywFr3FSmOTSvQ/BRKFjh0OclmOUuH8CiSPJ/0kXu4IHGY2hkoyJCfrvjE
zSuElfsPhGEONAKcZodgF/k1HvIx7ncucfZkCVtYnGC85tApm94D/5t2O4kR
wF4w1ZSAGAYrkOHuJThdOYQyocP7isvthGauo5b9k54dlJtpCCJ5C0FIaNls
H1HWfDdm6BGeYZyNhgTVDYqY175p5tYslQJkzZQMu2i31C4mDXyDoxmDlop0
qLqRAEGuOQCwL+Os3b2Cq3BxcHDyMkepH8Ar7eZ347U12PuWoj7/ECjhQXRx
2z2Goa+HIGwYiMttyNUvE68741XJ/JAN6xROi7S0f6TS0ckVo2YfGQfKGC+E
YapwYmp2iE5wSBlJHOXs+nD4oocuFqrqTeSfRyLJJvgLJW7aoK1tFPLyi6bh
1SzqS5XaoDuiABDSuXeb0JvBPIjOZdmIBsT3jjlngj268iLbrCax0WpUckp1
bErq4A5KwE1JWZuFqv7V6AtI8bK56kF0apLfRrTbrkmx89CYgku0ABRVR6RT
iFD+d58sYzwiqcJsjm8GK/LX3AiRoKxCh0aooRAdmnFVp3wU9ta5HhRnrrLT
yvM5QXxjJXDv0TZ8ODApby1uES3PqU3t9lnF5eaGbZw7h0XkSnnv0rwa5iqB
RKaxwttHf+B8G7iYZ9W7BZpI7wzy9LcFApl/60ZGG181z3iUs7tC0BUQ3AWv
lOkyRxG6KpUCttSAo7ssmyDTn6mh1UmGMWjcD2Yv81ulWoHCL7j+rjTVIrKN
emR9AqCgL8RGJEllz6Diq5xbHSPRxzZmzRrxTp0KNtF3+j6PKaq5SD5W/TtC
uWJ/tH0I5+bGvBIyBdWMTeLbAO7bOr/vPcY/5xxf0A3C7jS0fKqb5l6oyL3j
0x8lsuNkw7MYA65cpIV6wHkWJulBG9/B1Nn/+ObfQ1oyyIxQe2qaXpE/dnSc
KX5sXDyq0a8jfuUAW3qfNvqLbQIzTRi118iT4Ni/LY98lyTBFdtaCayoxrsk
G+idNs27r+zWps3dFVbsjgNK93BCV+ArWdB1Br1s4BuxO1UYNVcXYZWc4V+W
560CegmCKrOCvXvQdHABb1dxp8YslNDMkAfAiU0ANVK2hMgjfDJH7TeefTVV
qXPo4xcyk3PqCo7G7x6Xxw+h7r6VY8CZtH5lcSAmzz3nRPFf0Txe9DLraWHY
RpJA7gZ0pARkLjdR50olf4nH4mVg2fUIwfgzk1xZcbXKaJiRqaeDVA5KldT5
Sad6kDH3tcIOkLCCBHZ3QxwDxFhdlXX+9fuwn6WNCZ2/nJiVE7wh/xbvLpho
Ft/Ys1A750EMTPLfTEgE3S8/O1SIXghB8dLOubFBWvNw6l90UeDF2H8n3BCO
IeTX2/I+/vgs5fZ2WozgknS+9nyYIAafmNM1Y1rKUW+vT7nuoTVNojQ5OZbV
aHQQzBCo8llD8myQEpCNoJ/1QTDJCCq9zC80U9IAwS7vWNiYUiVKCppcm4wh
bfupNW8rfJpCgOQx7d/qfND8ED6tnslYOGhpCo3tzDeqf1GH/wEsd/ThBGyo
EnnrQOyC9JXA5ZD/b7yGEGRdLwte1FOJfV63CKdFbd8T8JX09UQlgKC+IAJs
9a3Z/aKeow2nUfYYB7qWVKXhXUsBfnmQBEZY9ono24NtbW64EBLSHAYb0c4G
FqFBDKkVUzs/s0nZ727O+42EJttNi6mssLYRLeTybSGbrvLrRLV84JR+vHX9
NWlNUGE2nvcKufqDmMFy/dih60npH0lX6KKEZLkel4BcUS7Z/m+vyNfSgtRb
qUPQ0VB4krhuiDyBNt4Rba2m+sVAF/GT7LvcuvdRG13ADub1lhA1uWYkgQOq
50QKNUdKvBw1GR2aZpHt14aUiQlx5uvdVro2BT4KP0DZb2vT3hQLSxGWrfvi
3dzHkGy6V3x+p+QSsCJ+V+3eVjvGnR4R93vqAL7oGw7viNYy4QmweCoVTh2v
hHz4t8zme5LRubh4yMcR4e2Yq+F1F5OVAYbJxNqAg16URNx8x6UooVvYpfpe
VwXRDwjWhod9JcwqmmdH08TZKF+LRAIgoS4TczfQdhJO7hnP+IgsDy0KkZBu
qPZCjfBl8v4tPLbjUxwx74yYtltJYFbQn9NA1hDh0UQSLSIa039kbfpD3Eku
jrxPj5CXC5FU5NCT/sBYPMFMe3q8KxIpFqxuT7Q76jPI7LUgGVjsqA/SPCh6
DrJzGHJZdFaYhqiCFuY5FlcWUJes8rBL7c/lBgO4YPQhl+9MslURVYM4pQhn
NO7OC83C1cRnWC//E4Qc/hqBKH5xWZLXycbvwq+SK4hPO4Ro1U74p/GlCJSy
LSGMQ7TCgSnY89K7zYLd1aGc4s+CuDjXCDaXzqNONHzC47g0l2xwf4yhlR7w
dKJpPqkwVa8teJFMlq/aYhMXpZARnyKiWoiSz4OAuQAkOohlbw+tnc1gaLWi
5TkTzQpAaIhjCng1VvfRQpgDY2ISeN5he1Fr7F1IlRkIRFkE7JgGp3Ktikv1
P1qSWfRSGjVkHoOzeEDumkRylNqED5wcNQXPbfS9QDVP8eICNZsJrued8byy
TxVy6FxbfKm02zqU7hqiEtMbLHIWQkOK8jt1Cbj/nC0+JBTX4L9Dzm3Nvq2L
I3bF5nNyBG+sskQnKF1IK7HkTx1TcKWXiG17Lbzjt9lwYKDW7ZQSc0PGZcSI
nKMQ70klfcX8pUvKqVTejEnlGMQoDzpoPx4yVjXSs9lS56pugo645p9/CP6R
4rqvsVBaNzV2Yqz/PyVb65dgnqB2BMtuIxDyFWJ7CiHUM260PqwzOejBjAfd
IjijqbtPZvl+w5PtA3cjXrXo8TkSdJHnsl088MskByXIY5AVP0q+SkMVpbJ5
qf2z0pRDr5lbcW/vuaIaGjsFvDRQuDKSb6wxpob+48AkRvyxgHDNjl+86iHc
ixYkLs+9Ou31I09TJSCSooI03ROjQ1kcUn/Ylcsvo54RtP9UcktMtRjmsqpN
2/LIEXwMzD/DLDfl89eJw/59AIRUtMdI4jdY0aLDbfk3mwPy40pKX7PDyE3K
isqKK5ubWr4/Ju4rqKwryb86zzvfcKq/72aUCmkYZNAdxi+K6Tp6Npd1kXCa
DqqepMJLv4Yuy6aJ87+MHxFi/oM9S6V5PSuocRrEE2QxjMqOcgw5ESZx/+FZ
PsxTkmtUiGkkZMlleU5T4Uwl9o1xPYzlAUD9KVIlA4ZTIlJ3wuUhOpwq5VO8
7O9s/tTQfkAv4XL153fMBgyvUtNHING13gnkrHMlZ4lmE8NVj97SbbVa3CZD
azfkYLM8l/twF1f0dGsjNpw4gNF6gttxNRvtEaGZa3RwmqgcafP6fPvACfxv
NQfiFeiVipH9Fn0wxW8VG3DYOW2q6tzY/ZeitVc/ss08chhQIYiRw4hOOuCi
skvoRFxhaSNvreEvn29M+Zhtv/7S0fCHhuhug7jS3TbCFdnlG/dyMTjRk6MK
fMk2+CIquKuCnh4/tx1YK8E7LNNDXWT3Bt/slxBAyHlRHai/NMwjIl1LrT67
H73fIwRfyGr5xhoOhN7h9xnQrZPEZpJMaxYFJMVhnGYc4iHLBygc/y7UTlNu
3I6hnWxcLQoj9zYnybpVzmkg36HakmGFOgrX3mTCEkUxapLSi9F+XOKLmU3q
IFebRSmVH/SLSmnLt9WWbyHzl8ijQ6PsYyhlQbYcme9McuYNYckgy6tvZyAw
Du0b7BH/e++laHHOri+Gd3Uged1xg+zjiplf+TBuWrphRpuUP7RJah/Tz5+i
A6YxwcneXuNZ9R7PNThUNBH/yYdMslIjFMwl/dItwJh0Nwy11mPnRWsfYvR2
2wCdyI+Nk9m1Y0Mrn9NS1JEp+fSkP5IBs6dvdVHq6ax+1ChG+74Bh3gV6oEC
8ESyag6pPQ8S1IbNoHyuZ4EfLgDTnjywDz1kWsvZ7nSPMscL1zvKITz/skcd
fnIemtqm6Ln+gbQfGJTnzrnEKfILdQ0r2qMxHM8OBFu9gynG5+auGlUeAzUq
5srfrfjFAcx2QSsZfRkcQcpVxCwMu/0cEscIoWr43ztomV3hUZeqEaMrgyKS
0jAcyfB1M5Ags5n4rC07nuzW+va3SAwwHkQRsDO4TJxXmDoMrdaCjn2RTZ/k
P63VsB5y+gNFcsucVCv9cmjFpGS33BF3rFAWH1e1oG1KEpyGEC4GYwSyntld
/YCIJavKuEHsK2/Ev2YR4jd2I7LPEukslthIBVrLOx9ljlMhxAxjVIJ0X90v
eTTbXYihFMljF2EODms5IstNAz5EdnvkguHz7YMAnkA7eKz4kxDegYhSC7Fd
oNPWPuGf46O2sUN1UY7QaCPKYkxMzYKhnwPtaDjG+KxTTP8nr5N+4ySah+0b
6NeVZhVZhklZXIwP7lYFRC/1xRKH7BA++/gkDeK2Os7J0JWtmo+VUgmgTaLL
4oG+lx2fOoYoPDpTxhyzMGE5IParP5C6w7qye5idAawEz8fV1czNsGuV+cs/
Z5X+H7si8NU2VsbJkA4mI0mIr4u7lPwEIt9Wrbb9A3g9MyzejzKEAIh0veOX
dmpOVPHxDUXKdtUZSecnI9TBmdiSkZmqg3ysVCdiDTAXozerKtzQ+JX6BMnn
/TeoHHWxHvuL1gLFnMzwHIDM+AkMRA2RBehVXRpDROLvXKZM6SBv+SEpKJW0
U1kXjAcoUPX2PaOMv6afAhw6/D+mC+2UEb9W9gpYh+TWOPhu729qyCD3qA/z
BHSgk0uGAyrD8BjZIZYjiWKJ/ufVD85ZrJS6oA93Ri53QuM+ysUd4c3AmdEb
mUyRudpyPPVvED4tn89YGA9tGF8Rtu62sPqNeVFm11CCNpI0SXwFCy4ddAeK
DDMVqMJxzSDqv8U4Zp2S93uFBxXPAMtR7rzGzesL97KAFWcA/NG6DgQcfnjk
uqCHsyJysVXDqAB8ZS9DrAYFGmFSKhjEXpplYrdzkQlSAre7bwTwY7j/XZKV
MXCo2CL+pMZdepC+exjxuUYjUaZXNfgi+N5SVY2f/Svb1JvFd+wEdXoYXaiz
f70CyULuw/yvi16qi7CpP4yCk1vhxF2zA6g0/EYSybSLAhqCPldCiqIpyXfD
uavEjdA/+P8EkRQ+/slDUcEP+4CM3obystx3OtsjW/ICYcZSy7UIiZKgiTtN
g7EOqN0gb91zMkdrJ6YprshcQcZhqBmaZGe4oYo4DHu4s1b96T4vmbBFgNkA
Zske9h4sheV+LV9+K1M3aymqI+jro34S3J2naWe5y13ormTKmA88eH6+o7hQ
MYSvS1aAV0fv+k8hurLYutxSP2F6PJFleaG9M+ATvC7ve8/KDHfaD2v25Fiz
F3lGWRyMNtEv+p7qZxmXcWe+rXje/j6G91rzjgf5Dal3Xy2DFzrB0ucLSR1+
RBdoqe1PDZiKjaLtBv8NnH73Steq+rQbyLXRJzY8HHmZMUGIOMg6k4gDmD1N
2o7MWQqVgCALYptUOw8L2OimBpIVjvnQzi1b3ffjFesbsUqrm7UH6AN+dzF+
c+Cbs9uAitaNX2/B+5xFX1iDBKTIv9SZojaRMmb5z3OghTnukoYy1bwGfsLl
qgeCCQW1Oq8+JVidf6yHSi4GxSkDLVZlUbriEOyPd9qOxLAF0h/t5kD5utmd
XUbCLRcv0b5XVr0uKve8WR/4I4xTLhb/5/QC82umtMEcPLVWSnux/orLzoPs
8u0mo6rsUGXPzlGs1wF+Tq1jwByrOW7dySdUMFljMJOLL7kCnlFN1KL57h5w
1Idyae/EzvgJgGrBtQiwnsyibWnlk+eL0LZHHXSQjIUhAE28aQrxMP3QEGbl
7+B5921TK+CsKzuVPKbQV7Fnxj1cvI+hEI06NwoAptcU0orYHTD4j7vVT6Go
o0cWZWxfVXwhbD366oL5tMFTtAaLKRMKjgglG8roBNjYUjOfL2vGJrzHtJni
yayvUpX4VEYfXpFbsldu7jQrB0E7+JlUQNCt8eNGVQWSGDMdlx94S48suTCq
cDHxK0u9bcMvhMMrDAwoRi15L06QoBTmXqtG0cod9BjQDP9wyJddxcugGoMw
piqDAVL50IArpkGEUnYAhtMSAVDb8sYqBvl+DZVMcoJ8qPrdzRIe0j5xC45L
rBRLBgZGPzqAkxPWvye1kldiJ2j1taP3IFdOcyMJVshgcr+JCC9DT3YXftEk
SL9cQxvzwUS7XMx5gc6A1k0iExlwBa+xCn+Q4F2CuE7fJk1rfuJLNcLyUkQX
IDs2YGaMlax9LKyld8rpc6rQUPRaPTYwWAI2QJrcBoeF/UKwGgURs47wHD4X
R+ICsjcOILmn3RXx9LD31ltumPZLtjHzL9MsIOqhUWOQ/B+PEIvfs00GEJku
mbf0hwFsK1SJX1EKrrFw3GlzV0RpQhp0ROOHUqGaPe0fx1KXObi7wntsXPyo
RG4s4GYDlAOuFJWibg16S1sDj1mB9tjW/Ny4jSOCnyJp5+rXxNTxdGqth33e
YEJSuPz5ni6OiLqkcgNWvb9n+w8pSH12aa1c76/s0WOJPzVEz1/zkCPvb/xH
4hqYED06304C5/2MGC6sr6KyfEBkYzFJ4VlP49sxM5wltUVhGDVXxOA0zgfz
LdFjKyOfQdm+h/6EWLO9CyDLZyn1Z8LZ4pMFIQTuG52TdyOUxsYIwIPcXzHw
euP02Yz4LerpzhfqiW0AwdSKZHUu6SSUGcRZHJAVWYaDbMGudbzB5UUr+Wpv
55J2WUlr0fg9I/W3Wjb0tOeFbZyQ7O/X25aiOS7Bq0Q42k8FUdaoDWqzqf13
MZ9hooCwSjDqum9Er7w0CXbgC7vldQNew8NJTGrgn1yB4pMs6dmmbtYC8hlB
wEmyIexpBKJRP8W119HIyHIa7QzYQNtjzhD/uKwzM0tLcaG237IUMskOEBv6
L+otLz+uxIVQucdaKzX2Rtn2niyp6RXYH2jKiXlpUrQiQW8qq4m7XxnEsGy3
zjsDgO9wiz16fzGCy/Dl2VVn/nas+DaenQf0OezEOJRuojavWyXCqh1YX6iZ
xWN4QbjuMrTGvHTelGoDdz97k6tbfWzQOLv/2K8ZDAVX+5n73AcWuO4zLoRB
P5uAnAaxTt5113qdvAUaJmmXd7MGoAgQ4Oj+SpxeqsHz0PGPwx6P4NsdpnTm
o/01w+P8qSLL7gF0RnNTrCb3lkXu9aqP3OtO6LUJZE4XFSDDqvCJhN+AhcqB
Ek7viZ56UdAT4H5RzcGPWI8g/3FVQ40fQ1t0xSXxue1Ll8V5H0Hr+8xPWpaC
A9cbIiAmpaJ79OazuwV8e8FJWmAeUgz/Ywy2a1ssEu+4c+tiwgoe2A091N/p
/JBVjXeK3B/YiV/T5lDAxSs6joATkBjwEBxG30T9Llmhuqg4Q1Oyh/jJmwq5
prsoLg6dGQlfEuDkAanVqrpa2ehBsV1iw7px8VjbIikkdb6QAb6iwgIVU+Xy
5zrs6TOot/vMTPeBLRST9EXWdlSWHHMPkCpJ+N4hp85kdty2dzxLhJzA7ePE
MJ/o/foYw5rXbiOtZpcNRIq//2uVbQpQDLVk3CXa2mMToROzC+WyXXpmwCcx
tSmGJ+/oBXyAvqRzDXdCnC4BfumSjVhILwyjPP2oxS6P1Z2Ix9o0LlSNzpvS
fM34zeV0LWQrnPqSey6XzFoaUE8/F0sf7SnZ0r4K33EXXE0pXPqjyGE2xT0D
RRtnq17j4VSUME1cShdd4nSSEeAW4FyTMNxopZfEyP/tU003agE48M7XlDcX
17F9NTYhLT5Xq3AU/V+oXavjIHdF8pQNzbXQ1K3VvRyub2Zf2YKMgc8UnMTl
cRwCz46JFSrh+ZGLD7hx747lovadF+eae1/D1Jk5h9DULuVgYfrFOdrJA6Ph
7VcsU6ja572PFkv4NqxelzdM+OYMeG78OjK3U8zzYA8jHSuXdpIaJT6dvMfe
QgJDw8bo2ngD7wDGYjkvYaykF5c1we1E4G/wbSPHxIsBLKDJhvCSsQwacvOq
e0lWLS/3Di4FZFHtS3mPKUIrM22pwqm7+ICZQh13FwZfkq1CshzJE6mE1Il1
9tekLyEBt6tUCOjK8k4bUxWch0ZtssJtAGZTkGg+J+lgw3ER8hMKiHr3K3B+
VeQNcvX36Dyy0S7qF4FlTbCo5tFXmpVmN7D0SCVNYRmC+Q4bDidi8kj1Wam0
SSSWiqdRcMi8H+mJPzdnByszqdhMnosN/6q6WDX48cRPwCeS12vLKF68If6W
O6ZGXRA5wd5txxeNvg0SyQbduAyOoVJoxgNpm9xTVZkHWfnkY/4ZEKRn9wqx
aXb2NyWFYPlDUNRD453x7JrEO03xOmU9rB33l5Le5TpaVq1+an3Y6sWjC9Sq
ud4e4YDftqHXLBuX2TbEkiCz+RzuM1ZPDWnZExcYXXAnexgkuaO96AuSTEkD
vXnK7QsnWQE4UxgdBKKJGNIQyTUasmP7fit7dzzyp9ypH8NXEmwiAb/1tMsq
8ptvgDwuIFVrys2WCN9KJ2v/sO2IizPCBMPEtI/PwiR1sfs4fjF1OnHj376n
H/yop3x22y+KGKaWOxJyIu8xj+etxKu7AAWHkrlRtnrUJ9upwrP5cxan6i1Z
BEMX10MSRQcol1OBwccuVFT+oe3l0XqP1s7cq+wO7xEdUk33NZM2LbvJijpZ
5+0pFFvoxnipooWjJgEcc79OsTYhw4L9AOxEfWVJTV4nEiimD/ac8854YKyy
/lD02wW68siak8SNqY4Tph749CxPsTg8e1x7gIxSWnRVmsLY57FbEipKfmID
T8hKmq3eNSSxN5fUUx8pyEDSncuX2HUiVgDQ8drE33d4N27D+49IgYSQOq8O
K5nqbRHY+X0SwsbanRvm9xKe2IwQksrO8EABzisjpFMHRhX/yfrTtFBGxo/S
WAUdVOB/BP/yxAJL8xWk+wlYS9KuhbbmAq7uahn82tZ9/pvUGTspAeU81SQ2
nOuKbdHMTW1dyrwBbL3ZSbmFpv5Zre9BvVO8TNRLGl+eXMDVB35DaPeUvzQt
ShC/7s90RHF+mNAUtS8Ohb9Gxoc9IsEZ/gsTMJZGikfp7CwvXdRPFQT+KQfD
xYT0BZwXnJ0BkhWehBZXMmCL8EjUTFm/tY740yyJ9j5kxTyCg5zE8L2odsnc
CuYpvCp9IYCdaJioojhf01xSBtK/ODCBcgZHeZ35ou96bSt+D2FUakVhhgMl
2Y2txhi4NB0PVPvoLk38FgavCliM3uqQKSjBV31qLbl2g4MqCDN6e7AlE1zN
5zY9O6N9upqJSOMVW0J/Hm23Iw5HMnQi2ts81Hi1fQ1pdaS7l8p/uF5SjUo6
KqLNri9GbBIa9reBLAh3OfODok4hxtqCSpkGCF6S/2yZ5BgewQ3XNHVHdvF3
y5dFGJFpvXRBAIHwLkfNI8PBdI04TB/6dftWcFhvlcLLstO816DbMSicN1Bg
+QEzJK+/n7Lu8sn/JNhBn66zPulNCHeJaNTNkAWOqemgqoDVniCLUP0dq7+P
4TyXqBoyNwOj00nVqLN4NOddGuTRNGNWb04Bq+Qm7z9X5tk3PID4Hm9xa0Cu
6UuaPB9LXXqHPSYn1XyyC6v3pB1EbVnLiWr+38QmgMoiLV8uV1IBtvK9jRtA
YJz3Z1dYhg3KSIEIluO/EJCkpvA4XhdmwlZoaPFXfEap8HATgAAT6Le22+0r
Q2nIj102LhCxn0w/5/ZLPHCj0AD5JqOg4W86I4/6f8YCUJaVhggAOzIaUjpd
qXRTwjqiGoQKp5ib1gnsZA98TJYZstZXTtpuSXbxnnlg4K/QroiXOWhK+sxj
f41KC5Uj9ff4KQndvXigEXnVDgIsYSGBUwdrLl9XaiOrsZ81WHRThF5XApY+
ejKHf6A5/7uTIt5MJ1q53ykAEdubjhTIulWnYEwGTw4q/kjlPRRiUICvHWLR
VceyCKNdKDcAo8f4CkyuJBIPuNvVHbRcLpAJ9JDbRSVJdCsOxGsgH4HiL1S5
qccsQYyHSq2wWYWNeYXePBy4Rmw+ozG/BVDgtVllJqbweeCrRbw5Ot4Kr25c
YbP5UyERf/GZa4faARUnuqR+LC1eu1n6YCD6cQlTGgoYha1EnbonuraSgW+y
nr3Ynzq0cHa4pXa1oFkY2HTPzgCa+kdofXEn88rgBUOZcV5+h2gj2IVhIwSQ
VOT6lJRvKP8skqUNYWRwCKcvTlwUR0EVvVPd1wAGYusIdrxF3fXX99NghdSa
N9Try19C2Q+NYjVvCGqe9xUe301tKVSat21KvVmJcDOgLLYWb4qEtMuCbKi6
HzaiJjWsQBeQ75fHqILORAPXvtT7G56BA79d1T8p7fNMKm6em2iuCeWiWaJy
HH2lePPNSwx3upDvsmeiLndjOBQrmnap1+uQcZMEihXw52rEtVwmnvItfK4k
94UMBLbfv34VThox2Y/PFJt/ovLCx5+cW7tvatfsx8JtBLKAkInmsyQUvUs5
Aw3KLddsnhJTl1Q1qb0dgf57FJGVgH1TmrztPDXb6EJUKrRJZh6GlkhsQgCD
JLnld8a80hbc0TaOfgXJVaU2Gx+u0LtFniTtAd1H2hpx5Ksm5maPczNYh0me
SfyxMKBWxveyy14t8kdvICJQ+zcEb3V8+nbe6yjVtLWKtM1W1tNSkpWTwe3y
8T5OL4zqAJPC8DCtT2NwSicqEQAvpGqMsgieMj5hJIvsxeeB+Fq+/ywFPLrC
E/ukPV0r0Iac0tlb9F/662btAJEcCDBRo8ypSo6GhMZHZKxRicQBDNUMEyXV
8X3u2dIiykImMYrjmrb6Lm/EJMcPvpUieqh4oVoN9iXgD72sMQpIP9Jp2EVE
gvwD7jz6WN8ydOa+HULUjUn4L0ZLhZ01rLouFM1ECrb5q01EQpltZz+BFxL8
IC7am8xbTqH665ABnDWHeFt+WgcOMX0pAIflKkv+SXGM4S/ZIgkCG1NXsjcW
bZ2XYyw5oNBJQyVOwerVgFPANzksJjHA2Shcm2QpRiaLWbZIpBD9gI60mAjl
wb6QhXtF6Vp3IsLsKxskXQeJn3GMc0y+O4zyyMuwPT60Jb+wItyKzpWjDU75
EdWSqkXmDJ3U7rZxHnqJjOksiHXzK0M7EVPsQP4xSd9q0pMMB0Eln6Gi5hXj
D3oI3kEH8TaXxbuxa/3B8Btsm6y1PjmG8AngWIVIltmIe2fDVOr4r7K8yhAT
mH6dXP0M0TW0hkTijn/Y/4w53PwXDxOP4uqdZTOZCmsZUrITpGQe3Fy6gvZH
a/rdwDqzvQZA+d+Ew/LWJ7/ItH2hr8ieWsWdaHPNNMRRYcmtkDjho7LurrRn
wbLoU1vYaZS77x3Y9A5JJPSV39T66+98/pcWLit4s/gB+D2BrDAWBisZRsrC
1/Tuhksx1mCBdK9G8A15gWFXCHOWloz21lrU0Ckid1B2thQT2TDu3LU9gzxx
BIsXCrgDCjhqbwerjkqN7qY7DelC/8zwdBDcBglrN34klJXUOqhdoncv0h8o
owNF5VETLOgZT8mXjNpx1H5TEjM9DJ+kZiGYpEfVjE9DMn0uiG2W46h+5ijb
k38vS2i3eANueftGrxfOZZlxG/YU3Aj/8+Q+pLk0vlH+8FjVkVbETY5svzBi
UeFFYh20apWxhgBZnDRvGWqk627TbHxmFqC+Y0SumkZl406P3eCM+TzbdwBa
wEBPkXG5BqPKyJtsFm702d+pB8Lr2jKzeyYPWXLdoW8/YBJSORYaWBVYYonF
4+lmBZVEtvj0728RX7PgB8Dz6MRsFqVha9LtaERd4jFU/S16dHyCNS5Wdud5
WEM6NqEtL3g98rc3++v3qsnXgrMIRb66ebM7EPVqttA3LF4tClFyH06nMRpU
Y+CP5Sc4XS1z+XDAalWnByieoXDBAFoRNXdc5gzmhiMdK65cJe5qlMUrHwWJ
XLJ7oWPS2wyX+JjayjFxHas5QrUEOfgn4Z1PCRmr8+2OODr1+pS5/U/u+soW
VObUtV+S5kZsVfSwiIZZUlOOI3/47Rfg/3L2KMbryvaU6cVBfCpsg8vtEEc0
YjOBwvATlbb7Mp+Di10ZKwXpW4jiyvxp/NSKQ/gxDLnBE2QCcdTXqiyuwJvx
9MJJWRXQXhWoDYaMPczQmYAeV+o5SGZTrB+LeWtQcNaD6qLj3KUWZ2zP9USF
C/vTW5gh30GLCFHtOHE3U8pk5etIdDYfUeicX3q22DFJvWoHGthmPljUAe3R
mg0v3Orlqt6wncRjm1gcAXbsMbxhMVuy7tnH27nWsw7paksbw20p/v1T/g7C
/1d+oyrizj5/nZOz2AsBCnXqnLEDXvYW6l6mBCXVqgfdc2pUfZ+4kcgodZD3
PnyqauMilQo4CYZmaCLLe5YZ/9kdqeCaCaPVMY1XM4PhuAcGeyWRNQIaj4NG
LR7P59MLCKHCDN8s5Stl03+K8VXCzi/Xg7rVitGHiRMYHyj9cjc8IiS45930
cQu5zndou0aznjWtu/cHXgauCV9P2m/zfTH7s3iMtnP9sNU49DU9WwRHwwWd
iBjdW2RDm5nln7GbXcxYVvxGE8SNG8TyHRb3rCq+V86l/KkPQFxrmlRXyDj/
ws8qvUPB2QXcmXunZYVDBBAPdeL1AKpaSBlR7KfxFk+0uEl7mbCCP2deZF35
NoMzfn8d1+DCZ1TQK01S7Br9SL0N+nlOOUQSpVeMMPARMeCeCPWUYXuS06ne
BLs0uRjZLuRZOYgn9W8KW5k1Yj1AOIGnbwJa9LKJGqDTJR6GR2m1IK6FI9JS
zltM0SsiunJLIO8rvajstPxxZxVLileiY6uiVPt89JzkLWpPbf4ll5F18onN
6hjKgN86GGF6Uaabiyfk2d1xtf6DozsPYlQ+SoMM9YbtSjoekT0mx29n5KfK
3q/BaEK9VxJcIIlagyAxt7deR8ZyaIg1ttEcOW06V8ldrXQYN3KcQ9KhwPuh
/vXWxxG/LbVzgftIp+bjVY2R36l0f+/vSyU0EmDcDHdWMWXEE9PBwrzANdlQ
9yEoJCKHIt6dlbwCG58RfmORBifyKP4kQDm0wNHeqxutujO47wOwtN6YCpyJ
n5YQ4IQCbSALm3B8X3B0PYdmPcKk7u1T4C1AN19WcxFurJ6slEfX324PuW9h
hpQE7FEgUS5ZzJXUWB0lbfDgpiW0+56HRGvi7PP5ApztlWGlXQGD5mxoUE0x
maoW86SNwRJXMPOygMmBGn/Uib5Y8k4TSHnstEtaM58l4Q7s+8CxE4JpmQUG
MSZVwxZp3kCwq6D3JoBMV6vxetvAbQQNaa9BYvKx3P3WVOkr5zlJt2zvo/tp
K11zI//JviL7raSQmJKpSekysEEbJcOYaQv33hjjZ7vgUs5z1GzIcN8QyKJf
W40vJlbFk7k4v5iAe8HzZC2Oo1fEw83cRxSJG0ta1JBSdPHlL8Jfrury7Qii
PZf+STRjWk8UFls3mftLNOWkVoJU+Y5azUbQuCoo3m3WO7Ubb84hINGbmLRA
146MyfVBj3HS6FpfsMc/TMve0SnPi+LbBFVzMZjHYnTyje2G+e3hHqqxFfn5
tFDlbFJkh3Zm1wDvyzR0fRU1wiRpa3Q+dVhqTEbssYLu7Y/BFphdrd0xQHHr
3pGchSFbWTkiKgyq/7gbR0p4Zawm7O7p6MT3Ibrk5rc55naJhZKKWqxT17DF
D/X4ZFdWLj2TpFafqKkYZKbvt0GRTtMtjleCWeuivSlTkTtzoVow69FPPczp
X1tFIlARPF7zfivbYp7pni3ue+w+gJ8R8Qt/XM2UeED0ZeHDhCcEU9Rql8pB
dCz89bE+IsFDK6PTMIyeIRlZE3DGTQjfZvX1c9R7yQ62OW74YCr+4nkQcsgX
1P0dgWc0NGteRa9NkZMY0E6oxu5KppFx0j8a1kZqHevhkf3ihOaYVvfzUFmF
vPdPfLY+S1wvY8gI54AYO4U5wfHC9z4eHD1amwKvK5rRfIINXp2VmTLDmSN6
Y+sYEJ3lnaCVvTVCirJpv86f2BwR1ux7CNDVrm60E3p/RXjfn60w0dqOuxLO
nYSP1yOzi7DStq89c/DCelqongJBy/pP0de59GwwfNlw2gkO7g5s+dR2gWtf
kj/inGIFBLkY3dCrzLoi/L7Ne6AA+ho9lGtVeAY6ZnhwG1Kc20Bdbbxh8EUz
A7JqrZr929TZOUKYIOEWZUK+eOn+slfGgVLcPWMu1mtL1EjRt8L4xGS1hPy6
c9cDvG1Ai2AGf4bmsv1GZvllJQUQpR3b3rIVGWInHH8b+z3rIn7hsvO+k0De
eFeNN9V7JTOQVm3GWQ1VS1COF/GSlPa8gbDHsX1aWEa9GUiBD8xxbPLAXYt8
dPejMPNh6utCrVnPDvlwjhEpQQ4rPytsK1CU9offdlvM/Qrfv96HNv2CfGU/
qDA7fk1kyRwuDkxwgGDIO0VOf8hrVp26sfeAplhkukBoov5Yg6TRaUgVg65U
B60hoMuTxMZJwLQ/s7dLQW7d0NjCEwS2B8UtPYRU5cP6GdxJb83o9dFwR3LK
7AK1ujHho7Nk3Lic4LLmrQf1uMfXjSyjocnr70mo4IS32rjpGiE29Eh6YjJo
GBMOgc8TyS2Doe6SezMhkG1+vGf1LoKxz3M62EYgie6FtDt3BTXBUY2L/c1+
K3V63iM5z22HGKgVwTlz5TstEorE6m+Efmt4DA6voMrdZtjbwzAARmzpC6aN
exd/r0IxlYOP7L38NiUZvKErP4Na49VcflhqJcsK/qDJBhiWPD3qePNS2pB7
NP8aW1lhNpAYz1Py3atlvbzqjt1ZTXzNeRbyHmGB4pr3uMOLbNCdaXpD3suF
zc+NjwlAIbJdMRdH1AwU84N52UwMkkwyWaOyWNcSmgY5bvhG4dVTzwkqACev
SB3cxdyUH6Ac4g41F4bKbmlitQzwS0PInbvIkXlIAIhm0uReArxh+AiLlRsZ
kNcInbxrog7RnFTivnpy7Q9TeMH8y4HQxIVAGEy1uNATM53pLwS5M37PTvZA
uU19VJ0jyluHw3xtjqKTYsRm8Z925fxi9fPlAJhC4keKXtI0PyT5OFw/IFtz
UoqV94ctxaiQ737jxOGL/G5ef8cfD7KG4bm0EHbzsjchxXb+fPjwlw67PMHG
+FNZjD6Xr2O7Ao2mEs7Lcx7Eyc8mwEszLMWAOqCmxn+OwkkavktESgpVU053
EwgZ/Lb1leNk9fxVFhKlMuDAFOZBJmRd0/c8Z6vpUjS7C7m1HXjvOvUFzVI6
PNmhVj05IKZNkd81RJ3yod5fjveSVVMuBb5Zcyq+1i3MoMyRgS1ZjhbNa5Ni
XhT8qaE7WRBywXKnArWqZS0UOUBDN8Z2rpHF9Kvv8NMjuC/bST1CqIVofjjI
ReC7yt27U9is+Mso15S1Izs1NEvtGSQeXNmSF2PNywKAYY1t9FdsXzYibwt/
UZMlIo1SoZbLMRkEl2XWKOSLUI8qeH8Tuauq94I5Xcrz9+xivEQIKKUG9Vud
alQkHsrYZvwQtQa+27FRC717rrQnMsfvYLl5MJssDR6OHynGIsbzIPY8e0dY
ve+KGK/TiNPsVM29ef0llJu0LxHajnoNyhOBdLCXtRhiCrdIDdZEhaw5vZwF
8dTeJsWFDbI8z9f0zN/zMXNYWxS3Kld+GwtcCpv/uL28BEQNVkHQY+k3J3Ys
8POF51+5A341ZdHLQ6ZE7+zYXbgE6w3nJlXlY4OtFCuzf4XZ3hC68iJLp4XQ
4tIyoKfv9XzSSIwZ5gQHHudDd4GXMsph0bhXmkcQWWnVFVvTTsfeNJLeHs5X
OBWkD+JxRS7pRQtqWuBj5KVdljSXromsCAkKUZTIociE3l6K3urjlO1oe0/J
TIROBes++Ta0z+GzCU4kFY0i2RzewqXA8aUeujKXZyauiFuK4BGMYayxQnpy
1qHpDr+WfECOdo2Uuj0e4TS47Rl1XmGOnCCUCsyCoQA+I4Yd8noESCH8mKgN
J/7pe6mBJOEneGlqMBqC//GWhlqj6/jto9NEXtQA/I2l5bqSJerMMkNlykI0
MTdAlJTphTSnFD8ocUEwcAWIUMJZjj4K8/kMhwbLebCJMG9ycbsIPmSQazLg
oxb6PTTp9bQRUOYmrf378Ya9+JhDA+c9nS10usGz7sY1dfoPfVXhObx3pOfV
PiWyVORKZJWnvf9C9una5j8veFhNnUuZ24FXjB62VrCnAhQXQ4lg/MQQFaLn
P4WKBXmrPo2gsrj05LX2LrjtjrOOqoVA5bb1X3886qZs1jd0mYCYAGIsWMf/
jf8szab6m+0GrDeXnm1GFjj11FqTmOcDLUXCh/0YQU9L8uP/+2h6GfUDCi23
95bjn4WK8RC5ntsgfPN805cs6EOpCXwmr2K53lUvcnysZMF+NDtJn4XYi44Q
XUS1PjLjamaxsRc57lulhnUKiGhX94Zclq4SwVHFmYp8vv1OHfITcArQ4HNL
pjk/Nizk4IVWF8zG5HngvKomYqK7mTmhZ63CKhZi637KgK6Nfa6rvSCPGOUt
8U2LZ8EkIqEPAfQ8pC1Q+CwcLeGr6e+5O5PaFgVaRWdVwQwPpe8Qz55vWYLe
5vMTRgOAPLHpjoo9d4LwORSeEBO7zZX8lXikWyue04sSFfCAVSTbxf1ycyYx
OYdLYDCe00K4u30AgqYonFkdQRIoH/S6Yhi3bd+oO5wVYIcR21QeGhMTLqpy
OKvvMyFTNKHZRxIF/mpEtbPLB1HPv4bcAoJPWGsRoMdlFQU7dJgzLCbW53AW
VTmBzuC1b58E5pAH69mE9Gh044tHk7dXBPhiaxAI4fwrOdVIQkgPPFC2cMms
YrzQx4NT0HUIcrXTHBgjoocJIHydWOnR5vdHGWg+pBrfjKzII3oXeFnAQ5pr
oDiK1ZHZMjwzjZ3IcbN8qKGMiVUL4uCSknwcjHBKO6GiTivWLyVlc3vBKA93
Lnk/0hv8IlB4kRigVPTJEBUfid+tmAvjLPY6lHIyaCdsZKCpZqireOdKxwtD
5o4LOsUWc6iAFcEEKIguidD9affi9C+eS0yXJz7U9AkzVUdarqVKMkNtX5Xi
sIFqYUzUqg3xlCno52PGm+HnrN8Z4yTV83suM7QSnSYSP9lMiIzlMU/B0W60
8E97bXxUyLhDsUjaSYlqZCibNiQQYfAyIdC1vwbqxhJjA+o8q93Aa6WTblR0
Ar8dOGhRp9OhleZIWJb4Yi3J9pqCrc41xHFPDhXsg7P6c5+pCM0WEimT27qv
I6ULZPKsgklrD1PQ53aiIcGpBbM05dPAqkLDl63BLJu64Zsp8FUt29Eigb6+
6s2y2HtdBZ2FFwYCYia4URjwtxcpmnzMhHnncL+AUKxNN02JLz6JjMAhckhu
+6+rYiwwGjWlsEJkXtDg/U+xoxdKFbeCZA+e0rZYQzx1RisUe/Q3YZQ243Fo
t6i5+4MV2yAnRMtpKod5lQM0UwyE0xrZW31elONh1sUELnk4bN2ij8i/rjJN
nCo/XPDvYX19bPqR7XMYDHgnZ3yTt+41olO07133AI2p8/DTQw+QofwgQ7pM
EvxrjwvoeldKNat3rzavu67wFUxWpatRAC1vLbKs0KfCOMufG6lzTvPB2kp0
nJY58L/FEJc5Y2r8K+ZbK8iGxkseiAr0lDRDEnJto6aJ5I7MHzRyhpw4T/Lx
82YUP+yUMxS8hZbsaAZt/nbxwaDW5W4IZg8Q1NOWYqgIul9L1OfzdKwmEoxn
QFqZrvuxWlLMNZXWsvX5whX50wN3G6TM1cHhCHh/0kQnln56w1dwdW2J/V+a
9slsvqB/c9YXy7XzeT8yOdA501L5qDvI4Iqebi7kzfyFKON3RzAPX+LOVdU0
7QRzVePaprNNInxWL3dv30tIlCs+cAh36o5yG8xgkMza22/DM+0QAXNwVU9l
YXDoU29PRt8KZU6kDdYdHz2J8cjRwcoO4hPQg1s0HqTgiH8F/hzbWytUxqNO
cfLk3n78DqQtpIRC1XyN3h9bc0hLc6oM365JqXz3CBIRgRZx0i3opEI1Wh8Q
ChElP9gMAADrR2huQgJeBggY4vBxA2uvLITJZCdEuWBCfRyUypgAKNmKxGxu
gQk+41++9NQaMj//+i5WDJbTqZo4GhoXOExjVHBdlEcU2MXG24xEkGVrl3Qk
XN9HuFmq1un/IwohAMXhH0DbWbR5xCXHf41/poJBtyHnwK1k3JPFvc7HGIQ7
gw4/wyY0bWjcJWaUDduPj6hWLCispc+wHs6lo/qMcyZtelZuzBRY068Plvir
KJ4rDK3JqqJGPxenWzis7opqJMtE6wT2pAmi+ILd5gti46SbT1w8kqx0GED0
ev/VHjnG8F6ZO1GXyhzJdTUxDMk3zj5fCXf/OJzqk2FnB3pmaa8hYgCPkz6z
Zp6Tz5dkWWWfVH5LUmVbgZT//CBSCVAkWkZf3jcLI/LA15ELXaIudBYO5xC0
W21z+ah0RQJHLtuVQqIsIBz74RyWV8cR884ALTZZE65YpQpAmzqs2iNlNRPg
zZ3r1Ycc5wE82sZOYuQDbDPggDHKPbZ9RTD8qfdSCWCYa1s91tDu6EfMoafl
1SUtYQn6d+1LqUh4CqaVAjr/ITInjmdF8rsYHhMoO1nT18Mz/e33YqDZq9y1
e5nY/p2s++DFYLzIqGfogL7/27BVykLcjJREFLdZhToAl863WlEUphsU63Te
luUlGFUBAxUoH6rqOicns/NPyMFuCBP0ZERqFPn8KVTS7H4gDDHhOYn8Xpxm
lmD47/4oO9VbVJyIx8SqqFnzs/e356ETDx4Ei0fjIB4l89gEwaV6GzfIQsFe
rGBbaPCzUWqtd3TW5goZoPVfTD10beuO2uECvfmfPA77TZYYmGcvsF6/sTXk
AaeArQUpLW9smOw/08CApym3m35ZIcM9j+Ah3IF0BWqyAB48acluo7548IR6
uxrjY9EV5xdfLgLJ2nLGSPvXli/s1ya3iu+4sqbl5JNdgkCffNmanTjgxeBz
YCrBfLm1/Mp66b67DtNndYZYMgkr4H4PyVAYwsXOkK181vyZ1ZzovpWtffG1
LJcG3aMaxzYSYrHhoiwMyUgaoGSw1cFcy56WOgf0gaZewmgdTPlZxyUT65t/
w8g8ovmKCfNxTl/IrMhg4rS+MbQwSrnxkK52vDMVvf4Ncv16GNTSbGOKdIs3
h3YtC+C1rvCU2ov8TObkyay9Ljt+/uMRh8urXGLubPcaEYNZjwVNot8Rc6Tb
XVcIVRH43WcwLYk5lcPiEN+H2ietOwpV3vSO6gT57qdpOE/RtaZ77inelxZ3
vLWEpu07MV3ziYqfIN5JDmqDDL/+7o7mmvm1GjXsdYI6fA80oLLtCVXIDRAE
WpnbFPQTq9w3vTRQgyqZiICkuRDYfNTE9y42gAjXyZHRavO4SqIN43ER4AsO
p8V6uNNreAI5y+rKKvatBWn23l8bedLBEWMjVmijLB2Mpg0WZNpxBuXfltO/
4C4KnPajcz9ayj1QW3xATPB+U17sIRzYEDjhs+NMqgaY6P41F1x5m0pCv8mw
Ga+MW+5nYfE7qZ1eRFmb2ZhMVEAbk81rklP6Vu3LQexpg8Ac+lsWvxL5vzrz
VjGMt+mI+/E884eyr5+SOlfRma5YgcdDFRaQXNSY9kWDV8m6wy6IXZvFAg9X
gd0YxUtra8am/e7J04ZXgTQAD8J2mNz1LokX29zr9+fEGCtJlp0lPi6zbVIZ
gJ9QR6+KStaPS+n+Y2pzHsWlNXbx0jKTfM9L0tdkl33lNxSCEx5SjoBzTzBG
teqCWz+uwqn8Gp56g8rH7fgdLUgjrgIAfDPKST6ygG9RGK9GTQut5MWlmSlE
k83BtHyZZL9kDZp8KS7gMXhkBBDi9HW/HW/Rt2+5GIPGPwizfhYKmDyiKjoJ
HNoHOBkmHR8Dm5tadcYKezf63P8SMkFk0tls0Q3sTTkN92Qt3LqoTwzpetv1
dtZLkqdtsX9l/DFCGtF3/1PRmojR0kmfk6HPK66ssLuwkk6IU3PdoUFu4L5g
N1P/14rETBP3W9Yz16+Zu9Q3a57VzjLi0SZoBVqeREpJqP67kmQjR/KIMrM3
Mj2CGVmP4PzN1nR+nt2WRfaeZo6YDHiagLPEKEfDkAlBUwfjlH2OBePj8+u9
MmWthtNCLBwe8Bh4yAO1yoGQCneL+/I4uLO3trAnxRY+nTe4iIS/ylhSkak4
TROrbtyJnE+RJ/3g1+5BzQwax3CIzKoT1UUtems/8KypEowy8MpWb9kj95KT
XPZEuTi6+5xEYDMXRBYF8BzpXo02ax7fIQ59sP+++axifRrht1aU2L5hqa01
S9oWXlN9Fs8XVu0o+Trjv+XFAhk9uj803bZFsWaOSnCukUk1/TSOnWpy7Sl+
w8Tun0X/5SyWWcAP2XKi0Tyahdfdi4eXcJXYhLq6q7Ax3s3BpaItaLiSAC6g
nxM+jUaHHwSymz2kCoJEPN0RmvfxNkyVZuLDvomEP9RCWsK5Faka/o2153P4
VTrx8NECHbEp9cXynjkN2geD9PaoEzGlltEazMt2WFAEANnYDbm/zxJqr/cj
tRnhi+ArEuTx46waxdRqxxiQSoNBLCbQr++kx/hBEkjIaEBAlqrgUx9Cwlyd
1Qr73D3lDAiJnDrktgghQ/8ovCXrHHa7cPfk6qgDuDxfXzY8clFhmbsjZWI8
sSDm8qKVfEqxWPvjV7jdx8zJ+Glmp0aCULcj28yK1JYTwJ8riLO674GIu4uf
qzh1yU0o06IhZDt+iARqMHuNxG8RVZohX3vTHHEZKiwC/iKYWFvK3hZG5fta
VAcP9HlKVs8/jbcICPlHZQgAfREwO7HRwO70clOvCBI1vu7sVt3kXK7eCZ5w
BTkZpgUJSRUa4tbQ06OTY5jWdafmvHCRfePt097W7WDiqwsm7vmy9o1TMQmw
F+37aIeklWmwobZuMkdMXeLFrul/qlFp9pAKqxfaREB5SwOryFYpPLUHWH/4
QmqJJhYtSrWWEW9bytGfDXaleNE5T8sZ1PfrKUvfxqHti1vtTvZTJkIaND7y
rYDhinE8DHfpng0P5S7EBpMm8R1dIUb1qPF+K58ALAgWYEeQ8sOurqNDeTB0
TfYhFRi9U+KqDCkITvK21sAMcrk2ZmMLN8jniqGqWJVFtVJ3TTmdBplpt7Sx
d0RcnaJGIoqXhV+eOpnbWVVAfJcI5kdbUJyp62SDzt5YWRoEKKK/QcJcTQmB
SfDXQqquZWroe2cfW/1oXGFVUW39zgCayeYDpufGjfNSpgeJHj363cGWxsh/
aht+ttSwW68tBN4oKblYh3j8O2YmxebZ+vxDes2wYtObAaVayA+2lj9bjQAY
kZV2RnUoQiLDNJ45h8UYf5ZnZP3vVf4a9GsxAiO4GEYgrykRb1pgiBZIdK/7
1/KC6HOfqS9vZaiaaGa2SCv4lZmRIeE2l99+62MnKyIFjsaI2aLILoKnHvfP
/zwBuYNpIneuykmcX3u+6T+wyHCW+gEgrTwVW61S7VYFZxHJ8kBAPziXJqtJ
KC2gTFLPHYjhwubLBUZpjChzhqTOzyTgqyL4N8uEbubpgYx1wA5qRShU3P2o
DYXY5giFnKV4CXvhEzz/miBqHdjfE+SsXPjYdwNs2HQR3pc69mUDEOy5waky
urIO+qrax2ajtDDoOXQAJV+c2dCi9atSXNFP3lwKCRqjtFwEDb6E0sy8iduU
wgjwRnwnv2JqGzeUv+0Q4b/X9sC3lFAuloc34v3c/akvlK9N7eCSkPFIjlbL
WxzzD8IBInxmGaDRhD16gPIqAlldGLmpvhAuRQQFdOeI7G+tCCkIWyDCvDRi
l/yg7ykYAGl+fu13BMOtFmC5hduZrEJVyzaU65ampFEunH/+ogx3IjN9V6oU
EGhxJFbmAnINR9kVyrFkUNDcNOtYk3YwGOi880XsVMFY8K4GhLaL1DivbWKn
tuWVSyuHfzm4A05FK641lGRjrbzDiRqFMwiCaU36NPWHRM8BEA70/zUPWs1h
liUaqW1qA2LlCCb04N+++JqOgDyLTXe90MatJXt0ZIElCprex4tMwqRoHEyC
hH4Ykm8DBt1niJ286JrqYT3m6Ps65Pufq6srXHgm95xHyqHViqRMiMkX7voB
AsOSEicRVKM2exGBPMzOh6pbGdaE9wruAAvjkIfg0hiuVXD2xavndv+rwNQd
pcCIExx1Yr4kE6OrZx/Y9N9CjpfPbU40uujsNnTvgjisqHiCFqR2znVF+g5M
dXQWrAEGbUUHejYvyJ8/UDFpNnMFa8f+6UudzfkfVd+ID6GBh4jKWQO+EI5p
298w00aIevRCC6yKPo3sknmbt5toVkr4KqeanHrH06eEcAU390nN23lS2gU8
y3BgX3FP3mLCkaolV2VDr6lsREiawfSeOsUMCb6KsIl21WoQd+9P3pjneiuL
evPOjgqvz5vxU9wTaoe5e6qKkP4uaiXT1kwDOHJAJODTD0YzRdce16OZXPLg
e44wHLjcdkC3rVkgGfe3mx+9dEpjpOz6yEhLE+eAuA1XKHPXMy40TIblATMu
k6VrlgCEnpVllKfKhIKbquo5hsP3d87Alpilmb+7StVTBezMdxDDIhXyLhxw
BCUrj5RwpvUhGgL4ePscHiGEjU/fiPsX3bL/67ik44T1xNwrwurD8Go9hNKc
OZY0WUqoq5jkxWNihFgHOg3ng71mZa+R/dQ1Yryu5RT83heehPxvwUDUltfR
h/RTbAfjQUO3CAYPmmx4gaQa/GqvjdP5DNaUSO39iKs0mGsEkXh2uvC4tFWe
1H8/m91lxbB70dwXO/gV6p6hdGAeZXQSyKy4j6qizS6NDzr7VWvKwLZjqqlI
yDP18SwPcS+ecRBmJWJucrO6PisBbVMOe2/Re2X/Ei6sYGKNwMTImmYQ8de1
X/syr9dCI73ad4DkGH6NcXRzCBQ1jjl/yz/qbhrf7fUEXwYdFvGj3A0nLX5Z
JgT8DXnTamqfgwA1MvUhkBmNBogfcVFAiqTEY6mSHanTbjUiJdNdRzNf1kUW
2k+cAiGTr0YLJX6chewJpBEomPiCU4PEUnLRv81+tyBLfpQ3lnu1Rp4Tv3Wl
b+dTXbsoviyFzWoyZWdr/qwhkQDGuo2eXSM0+kOlSLa11dRMaC+AUvc16yOy
l8BcWT1nCtCzwyXQao17EXvFDiP2EL1DHSzRKD5JfGf78fDmNjVStELQgVU6
0seZdKDs5yXUmnjPMU5/9h2V93A55nDOLnxDdtDSkP0XSpIZL7POjsMwTM9r
CyPbew7ZI7+TLzgDRXZrIISiAPNBAUA+6dLLDnzFkUSV45u11KLTrbiL9ORs
I7PjwiwyQ34d7NFKqkkJOhUIdCPdyTfT0O3ylIyt0N/OeKjmlSrhaMPttNjy
ixTrIjEfsKoiULpABYwQ+H3mkVDeQWhvCKU/6Bp9ASqXY9/3x6cMoO1/L6s7
Xa/aXVFAV1lHN9S06bBMvrg4wnkvRgEPI9NAH94WueKkv7QuJLPC+ElwK9xm
j113OkssWtNUS9Kkk6h/TiEmUzKFj6qb5Vjjcpcu2t6q91EwCevK3ORhS9/4
kwWru+waLibMc2v/wzyrQ6kN+gOjND35nGUYVXvK2iLIof1w5jKF/XmmPNlk
JpmlwPByWxGyCwxIIeUs6+om5A8KS6nuhwdQ0oYiMnE3NuRySZ0+8It40ayX
SQlnMm7ayt7vSS221TojPHnsda6kPQnFQEuQ+Q+gBhSXK/bvhzlUSc8PK3+2
sAzxoRUA2cTweQ3AVcFsQ+JEPrDmZRRQIm8FMSx3acu3ZcwJzbRBVQQoK9H2
mp7t6ykcNrjb0uYp6Zt6AJ8jVMx5wHmqE3wNgoVNOJcdKn9or+FzujFCohuI
j6Dk8PXIIUEqJJr4jb5xqeOn6B7bftD+iGUOMg1z2aGfeY3kM28NxUgWlnVS
lZdlasowkt/kch5RBtV5UrKCjqk7kdrUT8wYEsN5KeRvr9VfmmFoUTu6/+w8
YtoL9BJ5MaVwy/+//tY2ApZrppSpc7ILNkGQuZ2vaOv97wom0Deu06aez41w
rHhCJF9+sSQISpxWnlUBwELpI9Bwu7FHoiR2ZYh08n+Urf7f917FuyhEzaAs
+/jBNJ0N5gxwQOQ9IBaaqLemUOrfnRdQ86ybIyjfVLIenmKw+7Llqb6GHM1E
GqYDBPG5275ZPnBzuPv2IhgX9Q2/gxFYfbGuMvTyFHOAXFG11h8+konem95B
SDOEv3KKuqbZBFrow+nIx7GQLbIcapXYanljwvQh3PaM47qH7IjXXyYmpNj1
D5GXTR4U5atrFWN9xx+fTkqFAV768HMXwyV1dn6gYbYeaS/pNxFv4JJ0X3xw
b9IkE6NOulxZvvS021kojPMg2Rg/D0TDTtdDDX4NSL+pwJxIL8rr5GNbnxXL
rL/cwKjqM2Es+3I0vZV/iUrYKy8YyifPw02Cg98t86llr/LOkUDshjt86WOK
p5rClT6zV2gu+Nd/X+Txjx4WLVbM5EL6vYUAx/pzk7R7dClVUSEzjog7dGsH
Mc23jE2V9JoyA1KC7W4Se9vPystT2TFWLgC0QhBXa79ivaUY0kXs3ZOvvLqs
ooWc8hxhDx74F4gEJSiVVO3TDEFBA2JeriiX1p5rTDJLgn/DCCABAW/IFqe/
l3zGLPdZwu4a/Lw91WBakH4sf+eBx9+8gIK1dBkEd9oG92LipnfWUM0BhbwN
oF4ROfd4LAKljohA8jQHCGBYsZOI4NPXnSaqPLeDUmsCnaJo7h19MvLEmzsF
NFa5jXZpmpj+J/Aj/io3yqWoIwiFDhCHce4TWZT1caSrLQGAP3DaGE9ua/lI
cDiqBYW3uC9zHiQ961TvibTHypjU3VmN1jZ1ME54iabcLtPYxN2tLPd3O2zn
rXdcb0rxnS//Ir05dB/923GEkPpqkMKDQUVyX7kwjlgXruSVdrRBXWDZxNxR
R04rGXcIvVXXJdbdQH/2tQQttPfSjV9DDE8z4UWYFsVAmOp7oVLENuuY+EyA
jXoCWxDLQ7uCWhJk+xb+D84yCjk0tuPW2qpl4V29e4Wkr2qkeEuJJLLhL8aQ
23YRg4zVhV6lwMQx3bgwdpOaDfBHX9NbzhlWsz+PeDM30H7vc18m6Vnjn2Uq
+7QbLaPqTy2GsEtEeawPBa/zZG8DJXjYXYzZOn0bMwrvvQDsMyE5iieHZVP3
CbHPKExh0sJFQtkJSsYw0E3iUTe5yVpoxsYXsaXz5dcIcSKEBm6Wl9n3YFGa
Owg6G5PSKa/r0EnEpy53iPKVFvwBRW7DL2ZJ4gJw0jn2yQBqHbOQpHHOS5FX
xS+WCKfI67tW89ic46wGhcYvZb4GfddVYO26UezaQrggJwXbtfnWYLeBnIru
3tWgCVjMX7QUo4qJXbP2iY8H2w6hEaddf+8LQ+cndfeYoqiLjorkVx6ClAaT
JDFzLtHvLkWFtE801wZhZaeyeB5XxRxdNcL1NYUlWxePa0481QhaHsr5QPPr
LHvn8GKpkoibfuotkLIibpAyh4Q4HrJxuOcWdUS1kmAM/btkYXwsAO/xowuL
T80YH5lfQA7YW4sBOYkQ3NmicbgPEdSTXa8sjpfse1PvRoSslmQCR8v7sMyY
N58EzHK5+x2H2afHJT/1PZO3eovspFxlcelffkWxT5J537rkKwll8b+tmyaE
xOTZibKYCDSTaksSA0y42apditmtBdgUH9mb0FF3h5TjeoVNT6dwfzwwQREJ
+69wdEM2sB8+dkMhGHzsQiW6El0YebuwwGcXizeAQnKviddfPeZn9+Vm2BDO
FLomelynK/JyRobqQZ/7pe6HAmtkBMs8rp2Cg50cOWNAnC+Ih1Eid9EQJ3TB
sLCZ5eamAPlaAcvyAjhOfoa4s8LeQsgf+fQoBZV+tvvcPK/enBn5bVmAJFvu
joFPW3ENZEYbQVueOavSelDh2stGFlKM2XN3ZQvDUl5tfR75jT75/yEBORgn
2Rwnug9JSD00GD+dagsWVDnbGh00jDhJNTcVXL0h13uy3M7sfZWrRQGhBtCU
1AR+2dBcuHOUyefgoXJRgyaSzFAsNLk1QPhrzpOqp6cSZlnFp5DkrlwwDEOr
S6o5oQnrKY2peckfrDHMR6dcaR37B7gui5T3Z5gVnf34kSSeFGKxcrueXla+
25eQ9P+O2jlUtIPjCGApWOshAXmALEjGpyD8bFQ5Qf+4sldZiCofmRTffjqH
dmCFUkT7Cpu4Rxq8dnYOF0p5Iunmm+gqut8Lm4Udp1FGYVAbsaJFpSF85Msr
X7oxwhRz01m5bjYy1daETRPraM0+zXx3srA0k0Zp8VuvHxOzI7saQcjyTHSD
OvmIhONPHsphm/5vxkUyNlqNWFh4gXr6Ez4deCKOyr+TQnZ+uXus+bYEpRjm
ilCHRBGJZIk1fE41gymhLnc+nrIpjYyoD9Zsr7/17/l1VbcgzGzsRQ/g1U/I
Cm0RkTId5rfBbQXc1JevbFxsChq5+zj+JUyfOAl7yDXSeJX3UUika53iP22y
BDx8diOYMoPts6W9be9IaOTRl22o7x+gYerlQJcGHQLRKEzbV9uojVfilweu
P/3ysPcuv9Fr+zqzmsewaeO+eMgy1wjpLdSaMQjdcpchMjWLjZOaqacRt9hj
MyhvrIY0edBX96V6VtM3wHXh7OEdLWuU4BMQE+faGW28+TiyhnUmEJ6SfymP
DFth8yffWesod6YQGcR2aufwirPsZbEQYACv/3iqCyWMz/Nqlf2zbsBvJAVD
Uy48P/dPSfGo1uCqo89MRr3HykZaX02jBgbeJNEGhOnAHvA0+Sblwx7IC+nM
sqTGvnB/GlZb4GLYqspp2m3nSkyi8x+y25h363OfN/a3sY+8AwrdZTkrUKlM
wTcBTyRCkc6VuhmJG6/GrutEPuYUjai0bvCkaGXjeZXMjxeefvW/j9dTxTMa
dpdmGYQqWMQB0+15dE+hSEMutwBMZMLJNqhDxWSRyriNg+rDpNVyZXoSiNys
8j8C6ikEOOHrbl5FPsNdnkqcLzZJZzLeM1QBtbvtJIGjLO4pjRP8LeqV1of7
DbELuBnYG92z/FYOsugGi5BJUNvHuLuopM9gGNaYF53rKFuq1cvQoRZCvl1y
OSogznS2uAT4wLOnghOMbReaVSqtYOvAvDEtOSKmUfFelksdMUyPjqkvZXv/
6Nv+4sQWZVYFdVEKcVmhjtq+mz7i3ROrf2lHTDfn7lwquUtNrGVjmkOWQ2Ot
xfJxoJF0ppQ03EGE5zpkULqmiCW9qwOU/1cpHwNSwxWidi4oIFjwoLEjDZf1
xB44xrxNMB2p+DQ5tbF+u6tFNiroB90sAmb2QUYGoSoMdxk1pHUoclRAxT+E
ujLMQlr/KJTeXn66PGZBhgUqk1RBHbzL3LmwRpjYSNvXT4CQKdd3yw5Qai4a
9UY3IJVj4UR9cKIPQjEt5rqTK8edrFljpS0ZQ8SpSRPOO5PNH/p276qNRQJr
TIl5mtQjOX7bujyKXtuZXSRniTnz+7LuFqAr2TJthKDK3XB74d3/XmEYSgiA
LTptdcebiPfp/Dy7v5sMe6GKCLeuBbQ/i/xwyxvQk+P1KANuwa1GsGjgTX5m
4qXtAZDBUrr3EBzYdODETaKXhhJ2uZ25eGETTrn5MkF9NxMbNYN8StB7KNb9
iC8Eh3mgUO9jcC4Nuy8PUbr+iW6kizcpKvBkoq0Yz+ObxuXE4PqNACw2hQBV
LK1BRGz32W+rvgDL+W9bDVxaORLn44Ypl7QM0MetIR2gsIMr00p4248kQenO
Gvb8D56Q4oKA0Vp0gpiPfU35WjI2m6mint24PMX30V3O/eg2FaLiHbDPKDOI
s4uTRV63FrD0D8x2l/SZjrIsa1kX4hh0HM/KQ1WLktJWFRAZSa3rcsgJZCXn
GKQI080BZEDKBg4XUw8YLePkP9NhYWc3zio3Mgx6KaWZOri4Jp50hp3zBvQe
bCLKX0336LqAuBWkA825EjlmqExc8rprD11D/YKQqKliMRcqclPQU4pJW9m9
4rO1mPsJXRKRMNWI4hx5VAGyn88wnYvXp3fBX0G5A+48+qevMf3TNxSwg7aG
XSWf1XPMRx2ty0FiK5WuVKU6USoopDfY03RBiXNlIsX5NVnRAV7jedYcwumz
RAI0z2FvwaNDDKzhyn9jPvr3rQR58cwhnkRolrzzGo3IAamhGGe/jW/1Z3rF
B55mBK6x96KhADh3qozhbPEG8WicIKF6B9z88K25dPkLigoJOn9ZgjRbwXR7
nhFSZNqviwlwXNUYudU6OPyli+8J3zEGNlOL075uVZu5oElki/vbR7+8e3V+
sw5tNRRq+iVrdBehNtGOul0F7z1L5Rvd+oi587UEuwyccD9nzz76k2Vy3+BL
nlL0XKpa3zwXqgwmY+y2uYTmCzIWmIeyrGR8UCtIXJG6eTGvPbqH0ja8OP4H
nog04BTNwwyH8mhxWF1Uf/bmfeDKqCrdicu1tU5OnQdob6voHPavSubHDrJw
QPnCNKNnVLZPX/EQAZ04O/q1TxtYJWSCI8KGBhI0XSsEvAg7aWR37LNvAEsE
gatlE0imzoJ/PSZTzV0N8DtRiZs2duNdNUCgG8JbuexjK+KZNwnYDpwd+SuO
XFuLOooat8ZtR1j9ry5ceuLTwl3d1P7VO8+n7gsc+gn4T0lxFLsHaXHNWIqG
aRUo1SUjZ6nfJ2EBhzvubXnzXeNBBHe+faCtJMSVmXAEn+gzz7a+X/iZK0Kz
Lq9s1sJ1xTu/m70pm/7lMB0Qv4b5cMOnFz0gN+dMPQu4zw6mb4fBDBwyMrrC
rb2NfssGMLkAR+fE6wMUXq7ug/ELZJo+SgaAzEKOJkUMGtpO58u209VGG7e8
NfslQVRjsv+RpD7XzokRaK5UNceVr1BiVDEbv4GyT09fCuyvBbPhX4scNGdV
ohCf0ZUbXqrvrS0kOZkgbxEqhev4ezFiNFxCLVqb8eVkXhfyeTNUYGHmaSIC
Ev+xG0Ia1PZU8k0h/D0SBqTDUoItWdEh1nZaaRp+GPehAhlodlF7O8thtr/u
mI7kAebUS+BAFLpBspc9JUpJMd75K9Xs2+VZArtMouBLGAJphPnRk1FsCWBn
R31ns99RoNHl13rDvK1yZG9Bhu6d9ceNJg54MB4Qrv1CvqjZB7I40clDYQkR
Uwu/0FsbFARf9/wAEAaq+EhkN0aQN/5RIvLwDgPkvIvojb33KKOpqHVQ8L4F
ELgiLQZOMbeeDt1h12FDmEH1SAwEvR/E1D856allo7hR197k4diLSPdARj8T
9qQWNgT2uN6WegEj0MSceB56d7pzgLbvFKyQqc3pgukci3RnzzhIYZdo7UHc
eOUn9dXUkyKxXGLDQhA4km2P0JIMxR2p5UAkTawrMfgPG5Cz6Td/5lUzxEVn
XGi+4dJljdG7bb7QjEXOzhqXFn+mYpSwX6jtOktWPqmXmYXshnwLAE2P27kc
Er0J4tlUGb6CczTv1lMnXbjDH93t7QfYPXs/DLqFF/aHBZ6ipOjjGXbfsEcB
OOA5wWr/mwEirFXUcokjg9aVVfCDLEdH+6CAirXUkFolySCXefBD6Htz6Rf0
ZcpbR4CpsW7ePkW1mQS3bqWpVQLbpMXoixSEmsUXkuI2YNpd3uA+LC10jaRr
BGnazaEISlUcEkzidSPwU6VsLe6X8cK6qMjwjRGYug/KvC6W4HtMEvMOsPhS
M0aVZwe/EYkdLbrRnoj1LFTT5y+zI+zWhSVK17fFr1LVvNRoDivrWA9YkBAu
ZnmR/03k51uzzKt+oiIhOsHpQdf3PFKx3TOPFDgWtxlkkc9K1C/XIghskKMB
vaLbJZJAjoJsJW1sAnaHdOGEeLMD+PHNAuOBTxTx13yGjd/6BO2WTT82UISg
8f/gfgMbyfSsKe8yJqX/2eK5sUT5Jc94/oes53YEVnGIufIDP8iGrxL5Tdns
9jWZsqORCLpOweU+Zf8sbWGJLQboda61xK8HKvwstadK1P4D4WS+0KOy1OxA
hF095BjnsVozFQT1I3XXPDKm+yLYTsThJz6+mxdY/1Kgi/vWGyD7W9qAsFuG
O7D97Fmlq3wv1lcMR2NiLRaYS1iFhjWh12jONrErk+gyo4P16wuGAyWWzEH4
e1234+6BD/2G4JSYVaVTqOlgp7X11cBhd/Hf1fJVciMYJuIvosLM5etLpBy/
einDZhklCzx+Ef0LVtAmqSn8W0GHvtb45s7NBhncraETMnuO6X5sPxTX6Q89
HuGeL5N7xl74zFh1KBYwCCpIEN8ar1n8Hmb+t8wyfe7g3jVy6LC7oKhB1YuF
Oq51tMyJLN6n0Gn785nbcDZdydnuKiFWo8hE4m1gPclY8yYsA7NCWWGYoaWy
hJHkswppeWnkznbhyjl7ngJrTbq6LUyv/JkQqwoTSCK59q8DfKyGZrsnUCPD
YOy5/pO1oEkTiANXOjnkf07SLRmSoGVwtcWgg7aC2VzEwu+Oin0N1L/n+xK7
c+QXf8WQ7dSofJFJuO7k+aYGo36bndE5baT4E0tTwFmjz67fmonoyURUWHCK
5zCHNWHvLQ0YVroS2cHEdek+J0wtRTEdb1DqMVrG38jNlGpZSMr0e3wMIZQG
/Fr1MqnkH5S6btb71N3vWxKS68GhrWKmUo4q9vw7ttaibAQX9d9OVQJvAsFL
kEUzpUU+pMNXaE8/HgsYJ/8v4cNVAV1x7L/Y0N1QkuGKtRhgZkpkDHouHUt9
rGIaIE7is8u8ccEW8eyiuqMAVamSVZwJZXsRrzqm0ouyfud7KPLk2rE/LZgX
VH3dorZqsI9bHzHp3u6n5Mfmecm+Q/xIKWs1IU/bZiz4MuE/NyfPKW2+z+wV
Bheqo4W0bKDCRQnQeurdFYyni5riO1ReiRpxgqONvZzMlhoig5k+SyFTuUZd
ZJ3D131Eb5B+CRYVbocWLCvCk1pP+3IhDl62JXAVsVktzYoYlz+gF0rLGChs
FA/4Kzybn8i/n9t/LCKHpHufg+7umoSAKMrERtrDxgeoOCYx1Yz78kV7hhEG
cKTFjvk89X2YwriHtGfRLqMzw86SpKo6ZGHt56NjqwWJXolMRy6JH11rCLT8
AboFpFUas8lZWciUn/cCn9Kb9uqRrGoCHwGLWrhsy8siiokevG9uFW3V/XLw
EWJwBj4HjlcPAx53bl53NhngUaTL0+zViFKMTO10fHv6ZjHbS6iM2l/BO3M5
u9s2h+CkAbZyRa0be0qmtFKgAjh7dEpGXUkMeDj2PSgkiI63vVL7fjRaT5tx
zDwBE5muBgmalYQU01kg7IhMPwsRaGZOWlVagXwXYoQVTo942+aGyvNX+mxL
3jpEFy9U+awASJyQyBJ8qDgrjlNRq9fiUwr2T7/vyr+KviU0b5IBt3RH+CDh
/MKdgNwbR9ZsYvJzS9gabdyngE6EN1pJsKM38iTkshoVIDbH6zEmllGR8flu
IkqO4Hfc/np9WqPvkEZPUwSZ1Uyp71zr5/FD1Ifq0C2gO/Lbe2IFZhbD1VFY
P/VxVXqiY5kOhtVdhA4cVWeHs1uGM5LnEo2xwXwhQbwZk8bk3lxLFM7jgR/e
BEvSwxeMD6OTnn9HuA8hU7SOP70f04MME7caQVh3zbQWofBfofHc2428HNe5
CI69FnFE+gaGerSnyVZ8FlCExoQToh+7/UYtrISadeX0uHF4U35LlnYIEPg2
5Ft6FKsC2wHzSBx4gwO0bIuQE77rxtQqMHRN2izTjNXhxTXnAUoEjo6eHs0v
yBs2bcDMBjX9riFwuazsHsxSnqy+2RuUpej6bslD/UpeCO/X/g/zIywZgI2r
6Um8XgL/74qWt7yVy7t/y7w4DMZTHADAEO0yE0RB10jkRq8/ulrb4rOiXZg4
qdCUkkW66rFdhFHFstDxNoBXMB1iJhX3kZA3NGAMebAsokr2TdNJvwPgXCn1
uYVSBYLt0/cVAoWlmYrOKkBowF6Y+xKgM3FQb2BXnk7WdkJOjOyve6SJQLVt
JNIpV7PnRozyUc/4b2k7AvfUCKAK/T9sIa7ueeT0YuVz2x0lYi7wBoAd2/H1
GhBL2LrwfxXwe70Qu1gfjZqENrGWvCg6ewtQL93GH6VZDrWTu7hkDScZlpNp
/PZDORjgBUPGx/iST1b2umJpGVhfiebLfiftuycdfSvPcNkbHIi+rCykUHnm
ErwountWUEEIiWIvVzfOyKZznV9bJ87ddxWrtS5mEPS+6ApgWqwT+LsQ9Y2E
aXCTlxxxWSU7zeOv6Q33bogYuLulBKJ5Gz5dq1TE/g/agm6yBCFnyrJQgCzR
geVHQ0f4W5O0VbgzzdtytDtVFsGXEuJ1MJ7aGjaBAXJg/IJ1wl277pe+NoJP
O4MwtqSRw/fDaMJQkdUGv3i8Lgm3WG5Ow7TrpQ8/HH1MBUMM3CFzzfF5IBNX
ziuhNjz/nIDVLFdrkYl4NesKmyaVQcQwGJ+cSX0y6c4EuA5vwWOU3DHRGhPp
ixwHOExi5WgmOSuSd7FCbEY7Q8/dc7K1ZqR9IxWYQk0YZrklNg8Juut2IRNH
u9tKMkY05ZpU8dnluzFch3MFLm3aj0kCWWnVOyVMDMDxDYeatwGu2HSKBZTs
T+PsO7IOkAvrwBHqjoNeK/GommF1d01XP+1ArEJtdOyi35DioWFeFCvHiWg7
SD6MOTw+E4hRAE+wytYhfjuezn7N71Bte0ZLROu+8RdB+cKaPGi0/GtGSuin
Mi4+huPhrV69xmWXuT1AOxeusX9ZQpkONjsC4R8nUU41CJ2sAdzUfL5CaJab
50v2IaJIPwxu/HpAdOmTXZ04fOsrV5Q0ojOETJabD1idnFTjM62bfDETx2uy
VM/zr61hrOydOoq/KRUCjypIgKU5vGzfEhFF+9HWZlpWApcMHuYO7odChSck
p8coJ/VHSQbXUrv4dOv7CtZhuyC/zP21KvAoAarP71gV4okVgi56IMqvnRY4
8WGkT3eQqKt4X+Psof2vqLNoAUasXqj8jYuixWsYVhSJKRm3D8o9VXwHZe5/
ITAyPYBia4L7uVtlGs45cYtI6ekDnIK6vvYo7ySyHfrxJH8CLNCI+gwzTR+u
xGXtrrNYdn0AcgzNMHO5U+yJ9pqfar6tsOEd0gaipmJpTMth7rGSTWvdv1gh
cdOKFTLmgv3lS9xGJOmYO/S1b1Ehyx2C2NATjw/RGHFFIL92Z7y863MYXGLt
kCkLQmjku4siOwhgnTcU5znHaRJCHA5NL0smLkYgAJU5B6wt1/0w8LTNNp+I
dDb+jf+JfwbIFYTThtBLfJbR/kvIFFf8YFeuVauq8svRodpQTnq0k5PpTC2Q
Vpl4Cx7bZs7n3dO9u08oBR3gD5jLVe0DzT4ru1X5X5cS0sYYEZoFNqKwTQYZ
c83flMP3NySYPdJuvpW6yWBsxSEUlngpUvs6mJycA2b/4zRPt3kgxzf26aUL
7wp55XUC1I3bZ4nmazFHZqEr/dCY40dXa8i321UZoRsxrIIYP711leFNJUtO
BaIedcHPXQXikCMaB+w3ffbnnGPltN3xqFC/naqYSq7nNCxO3vd28x0QYNlE
mDszDchSfgruymGLnQibomfvLr48QOWdnUC1iwz/hXLUUqbH3XkxfRZiB3ph
9a9JlkNUGLFnzX2UMaprWYGFE9WgpoZIKmFCCBBdQBRIHHmdRfb46p28jr1F
jvJvhlpPqwV0MrfSHLwV1exps53QFtL5Pc2yg1gsFeWPNKk+Rbt6tamv8drW
XuxG64PL72aaQi0CxwZzizgyZBQ8fM4Ndd/UKPRlo/qynkuFNHLAE4cd/qye
bOMeYATh2O+FKvL5YCPtG4sBkRjji8Kwh7CndDzGpxJ1+RfXabOfqKUIjkGS
PfafvraVSwEBmGUY7HLUDsCorRP5iVz09tq48bckA7SxAvHV97vdA4j8FyjI
QzQU+O5i58GY28reAL/tYXipCE1LCrreIRmVCeQ0XKedUtqsSeepWeXjISFc
kjrHb+3m3jpr+HNDH9mn8T77bdtvQJvp20h6DNRRdViZailGip3QFdki7jDn
rSgfu275Bg7d2UMBITjwsfOMlL0eX0nXchLFQwkvePKU/JFppchJONuNxLfv
3DlMxCgJK2eWoeB91OFxS05Q7SCrIU1UhZcfbibF/dzMuMVUYmVWObEIfmPI
4INKm8H3GuMYom2z+XiSMcq7xgH1pJw1uI763+tHEWS0mTiRCZoN+P8xWJL7
tlStUEzAqmw9Mx8SWfvrNhCk1ogCtZn+Q3JYogkFZGdPOLWxULgrVkmI1Dp/
U4mjsYjRRJrNd6W4b88Uli8sLXvdDYzX6hIB1dsPNNOJOM9+l6MJzLD6/X4D
JI3559rHF5xxTy9a/dLLlza1kTmDdJ3st1hvUz8qwSgI13noWSeYKOgBthdH
35WJmTv+EstxC3mb2fiiMwU/3imgq6LXqC4P9PCFYTUzWmzIWk1sbBNnuC8R
Eb5Bry0C7/8SURQpKEgFNfnev3U/Esldcj2LPtC7+Sq6tbsuOHgc7ku9e+mv
0j85WzK0do36WV7ij0zrSJJiZgnGJi7fMnBEcAqaTIaIN1Qg8gGecom0sJ8i
LK+z1EN4BLMgwK3wM9wqx7jhJVIMaFcAE58FnH/ycCew9zRJgkyjE0gAyrrt
SNx2F+XlTfiWTchi+yAUlfgvjoblWG6upiEl801EgFobYnrifFXph4X92jT4
hTugga9h9XO2X+lKQbggwd/Xw6077B574kpTMkgs2Wu7Jto2CP0fdOJlQO00
t6zIchCiIpB9EfjkDsDw3PVhsWLuMy3gJRZ/gJvG1d+ERWKINhsNAQiM1DHB
j37eabqud5A2FVbJNDFEm39JxnsMHEHol5gi8EE7AcH+SpkXAjIPLqQz0H2E
hZZLPjuYpKHgRzye61pzEH73EoDwZaTuJ88SY+4t9btHtSqyqLTJssBiA25F
eApftruA0kqbfDjU/q0Tm4LabeAjBvS2xvjox1Fr/P8Ekq0Jq4us1t2mkPGM
FlDfhxf7zT4TTp2EzCu9uyoVT9l0ZpldP/5Sf8Ww4kNxuJ4k6T0uYG0NediI
xj7tIYblTLEvAU7joJ2yCziMBLQIPnMTIvBhfOdmkPrxcBaULzr9c9XPuPwU
gtf5OffrVsgpk16mNjOe5tR5yzwBtAZ11/mjpvqg4VQcrxezak7sVmSHKsWo
IPxb+7XSIP/7dBqGYJjcH7KTFLp7lQ8GZ29mToyP/2Q7Oi0in2r9lgAT3/9c
LQHLpwlpTHjJEugLrQ1j3wXH0NX1I7Xsa7SwjbW6xa84IfYo/aYS0/QI600V
WiSUbdU8UklyfvUYZM6lQOM597UZlDuDnx+wB2mq5EbTWVykd98g9RDpHSYe
m9vojAYdU/ADrrwpXghg2ui96NsWrfuS+beA48hEvCljH0K36Np9aqvXUMYG
A1+gU7F5SRH0SskfaLpGFXRoeWhzKidIfhlNqi1gCr+iqYfsc6WS8z3lxtZV
/V3qyCug+h5zBZcU7y7ayAn8qjVX0LS8voYfsMDxscsx4ykqTSxK1IJJqGzg
5211rKHVxBo8+B6GT03PJQB9Uc6CzTJvZcfNirCOCC/hGwlBTANotaQbL80U
S/GpWMCFsJ4ysOHfulkgOSHCGyCqynhYwh+ce9PXaSb1/vzBFhqByUOltsVZ
Bjm+Q/5IfeUdkheGHdl7Hxb/Uu7CnMs6rZOEltIb/KFWuLdQCaZ8Fx+G36Ai
kE8wIi4jqoblRo/1XcoZXvlPY1X3KdCgHRCJbILhc/Kb+CHosSKS8CNfSwBs
vXjER30CrCPEBjdZHLYoYmyfXVn3E+eDF/gL4ImnRoFMooyfR1qGDsdnTKSP
OlFu2hkarP+VSKO1MRlrxPFtBitrHVFVu0CphkuDR+0okB+sphS7SSAafNHu
XTLC2kDLbEJUjxRWAsFMg+iN2pgm6FgV/aWkMFoZq3DtaY5iJdTA+yNUWnrz
tHm5e0GkwP6QcjyaItyHIn6q+jwC4U4sL4DHZ7iOupR5+hQNgw+Hu+QUfKZY
TmTVjO+97szLjTzAv6bXIcGM0IgeLEfx6cR/iSvAQ/6GoHJxxQKgzRxl1CDR
PV93sLfTArJATeLNzKz9whiAHJZBlVax2P1QdKGLrENmmwg5idFSFYvzwqQR
vBMabv60MCctyhbNVdt+KFbBFBlxhDY6rxQ1xAYgQayWYIaZXHKcs02tvjDo
m77zbbPHnq/VmFk33kpryKs9uWPIMmAGmzmajpCg6TbIm/GEfq7ZCKeSoHJJ
9g2POKcbvJhQR1nCcdqyxL4QrqCzOwlCqk32v4n69fPO2J7yboDt8yHnEauz
ujQ8SiseK/UsvuEz12/Z+N/iHqZv0z4IDKl79J6Slq2i0+vBTRSkyUyOQIFL
wFsOsGJ6wthKk9zUF1JrKN035TYnDprFqBjpBqFZtRWgNmvbQBJ66UeRmCek
p3PpzGFBJdYdA6Bu5HoSQ9lp7dxybXquKLxDMXS1ElBlTgFpQO13TbZgN2d2
KucmbPa1NDuDs5zO2v0/t1B7DfIUQwd2OkwEyB/tJqX9C7efYmZ6EisiNC6j
MIESlzLbn8BJXhtVoxkRRsO7cC/f+xGxvQF+P3updI73aXT/YsQLZ9NoExVa
r/l0rxhJVOaLQTQK0gke+AGq10TWE9/SWHZcFwFt+dNHc1Kpb+wxuzADD+XL
LgQ9Mn1xyVyChtWX8a2Z12b4q+bYJZeeYwZE2XmwZ9mHy9nthbghzaAZelB0
Yh+a5D6wknXXBafzf+ZuLeO7SZzYgXZxaLhWoLMuzZ8FUeTAE4z/LXId/lxO
CmjqDeiAoagl2MQB7JnRQ+EGpxsjL4jfo5JDD0W8GoKOztOIBUjrWrLlrHOs
sk+KjoGmQJB7EpMxLcqoUGasJUE7svydAYEMuE4DeXTw10GXPMXA7v4vtEnc
NlZl8K57168504j+TJumdTHCm1KjTNqoiQKDODWMjxGSkQ1yHnHVT2rT/mkv
YgEGFj1C/ZMXh8AXYmSPXohz+cLvocP/CSWAP4ecZXtpBNq8w1qMg6kxLk0b
N1pvJl+s0itsqPG48zuPXyaK84GR/I9hgJViYRMu0O6HDLoYcFeZTaEZYkW/
AgLDuJCM+AJaBhWh4p/eNSRzmplJZwDEDaOfaTUUidb2h0YAeq4QopM9kH7+
oKn/SQl+0bJaQg/1eWUNl6mwAXi28hoCjoI0m5ZP9b8afr7irZtARQw0Dd9p
XuID4THF+duLnLcdcyLoa3XbJ67OYIW9OOQ7a6VVB/rL8OOkpqHfG50t4Vjh
9oFeXy3eoeq4MA4iqh73PmPdMZm/vzM6/nURYP8/uJ0konxJ4pPOsFFjKFby
e+6/zKPdpctA6XkjlmGD/bmXLprlnDsMonPWjEOycH/tkk+tWuidCvh1r3RI
smN0gZwaY/M9Lpj1CR0LYxcOUcW7bYGDRunBKD8NVjVilwKp001E3b4a6ZnD
+c65NUBYZJlbiNRV3jLcKNRfcdc49JUCHjVizFG6VuAraM3O63swGVqwenbq
acaCKLLseUMvtT21+bhOwjCnOe/7JdPj0vQ7Z105SKmX4L24QXQ5ZM13ol7Y
T2UwHW3X3LV0kUAa/tX06KCS4hz1oXznQO8Bz7FxRDnAb10qSUPBfJ8Hi8vf
oDAweYr21MAhvpMmQCNQD1peyta1d9hjfVVDtVE1t0TAxt8O1WKe7itG37/J
n4oh4vYrefuiWyK6FFepkfdPbTe02HsHr6H9RECYcVsgRlhi3maF++F2VCLQ
KizJ3hIDP4eE1zcv92f3QqODptmXEFR2F6QvoyJsubZ0FhgTiacpvX/MSuE6
v+dYhk8UgSKbfjatHtdGkInbVcJLmYbRmeSqcbsqR6jQP+xOznr4jwi+ZE46
tfc+5XGdPHIzI4g0tJIJCnfbU1rcChhYdIqmUMdZ87Fp2fGrbDWGMJcqb2Qb
aiaobVdNZgsgdF4c4/ym/DoKd3zKAtDQS5lISWRNyHpadj0bobHzrClxuUeC
3iVJRU/vS7KgSL0DsvDDjDHBUpsW2ECK43VHzt4mdoQqikbvKyCDl9xcpvx5
slndLIVUn6nrvN4PHn06wDQZEYjQDff9f9iYW/IDH1q8gC91+Ld3idwnFmnh
CzK6lul4boXw8BleQwaUPsIirrUCdvXOC6RhaOUoFsagGQfQoB6+hoohFr9i
6jcjSIjjKyB1CI7OHyJUpf92+Nb2GC5I42K8WDUWNlzHAJsMBEKnzj1b4MMJ
ASC9tRIZDhrJdRZybo5qGHXK4Rf9jYXG+FkBk8NlB6U9PvBlnIBlLWdswkd6
RShDvbi9XC1THC3zxXus6HBH8al6g7Unl1a40983a39HSZgxykTLixc6qFIt
z3553GcxWtYbeWa6q9bUARirbUBMiAREgZcL3pPKnelLpEGVF5ivXtAiSZJZ
n1UR0f5eM8QSIJ/C8YtWS6Y3pjpWhGz3ryROhxF3vTDMYj4O4u6/2cmAXItA
/Zhdp61t0uVYoz7nA9644yNot0G1h2gIQ2Gbuh2MsirOJFDdfwjkfAUCmIGU
vHoxvX01P1htQ/Pz2U07OewmllTQJPhbXdsyXavY1TTJwSIewJWeGy/HcQGE
NbLmMtpr17lPUVOOazM+D/tfTIK8SIXEr4TmzvefT5QFJN+EafvgYLx1XGNO
TrAMSmrpOq1eO+cbt8mxLoyP+LFq5K2viiyGlq7IcuHJCErZ+684zMOT4T3m
3mWcX6ZUlMJSg+1UzWFJ89bhr2NoHUXae4K5YkXmFVQrowJMs1nWV1YfWrG7
XyFBLmivAfP4dvMuuVPBD/D0JiZu7P4l8AQQ4gJnQuWEoWHgbyD3B66WBZr3
xMdgWrhooFEqDACqnSBhL0DBipM9GeHPvfdzaTcgdzulqP1yJJvwaoJeO6DH
6kaDzIt8/hIcPDpVu5BncK5jzR5y4IVl/TVMSKzmnllK13qgN+ZMJda3dcYZ
jw6Vk3C4rxIv4KaMayy3udbygQXsF2GEcUhD0VGVLyqp8CfDWYAVx9SC5FO6
zKDwsBXEZVlDydc4R0r4cPnmIhUJJr1SWmkeEPM9aCartqn9GP6muyrwiSkM
u9sdL5D50/YzLSGlR0Mn95bfgP/1vfJJSq7bO4KA6aRhE7Br6tkymk7bciSF
xpPo/mqz3mrBELR6rm8hQpkrO8Y3zR5SkIsMc6Q5Ws7XQvPYIarzDSdphck5
K1/lWGp5Vw+GoFe5vSzNWEpCm5Cii87av5bsXP/LDbDvjNKcpO8e+KbsixO6
+sFMerC3Sh8JXGES31CNl8KmFmai2UEIByuFjP/wH5CHmfx8S/OxKq84TQzy
mO7hes5g4zUR7Myxug7IdWKl3XAbtWcAbzYox6WE6kbQSwWF69Oekc29e5rW
Mkwf5dF2EsmUHkzuc4P+KNt6qoKsuXV49zMUIM6ki5xEYb/WLlhf1RCuxYm+
mM22X6pKDm1O8my5V3O7HAvKieb1VhXhgbSvCRm25a7muNlnH3vJtAywUAGw
EE13QRF0USDAZ1sFaeviPK4lI4KLaRmB7kDVSYoAswgEzVwneMc3hUteffaP
z4x6rMmW2NRajR0KYqK+BiFvZon62g9W/vyEDNMmtRl12kIkuDR4Y3UMnNpa
C3xns+nnsQk6U8RmPTqKz+x8HXBSDazBKldQIGGsBv0rRUlYQ6xGYZBTXXaI
vGO00YVDtCi52jdOEgxO5Pp/k3FIbyzc1QxVytVEjQ3TwdGxFFNgJqnQxMQQ
r6ACN/QGZMw9u3BH1Om4vCXk468CL7IjZuzg/duzbMJ1M9QSQ9R22/PPERF8
DQtDHTHbAjbi3kNmwF6SLzSptkuHXYfmB/viafR9vsMTfab9WlolHQY3A0Fu
Ke3QZ9ncXtk7pJOVkCSv1ShKnK+14BKhLLKXXWrpyuzfnCBa/obRNwHm2I8v
QR0i9CEABjGNfSRpXWjOnKXSdxGptqasqYKtw6e4U+Jp/L9EWeG1PZOpzCFv
eXR3bUgL2o4yZLGdZDnQokKsjEzRYO1qskgHW87ae2OcYcduOyHg85alc6jp
UmisTV6gHP8o88wlgJ+wuRJNG31p98WR4poGIbrR0uPzC2KgS+avPFRPlMnd
EKKEtfK+GTAdUb90HxJO+M0cOZitNqw7FYCxIU7ek3CdKflLvWWEU5mPk8kV
sYvDqjdRmnzLoai0JSdM5bxsnxhvAdNbJePM3EXl19AVRldUHXFlpm7yaEaD
dd0Gquiha4s5W7LQPODITs1cb7dYBXvtANRJ8if0OeRdx3rfWf8kq4GBZRz1
twUptRZdKSI/SDxDmFyuWbAr3pGKTcpxQ8h+fj9e0KW48vO3+RNyLoMFyEfO
26L6jXtUyiMSZqLQx01+BK9kchLLmQQQZm3aAoYJdW6NJs6W2lZwoOry1mb7
pBaYmvMHO3gHJRPYZTfHRRPOXw0lQJInWUnJDcMmCSBfS124q/H8h9e6X4yv
wU9YkzoPftL9NrshXStxNBtwa8UWeubuS3FeFfNuIEsPBKPiPM4J0g4vHzZ+
3HaMK2v+n8zSnNtjsvS0x7vxcC2MosVulDg/faMsXp+L/HyePyRNGSassjCu
dv1PwpUeDvgQaObZNxvIjtIHKMu1fnajsmowAFKysCElK6VCd2a4Sd9Jq/VW
5ZG3ua7Wj1eHEW9J2TQAnNOZcSON2OwQq+XcDKxoCZsNswqAUkywcPJQaSZI
qWJcSYXm5iPGucpCQSCjoXzXfdPZ1rpPiG/a9iUy3LpKe5ZCT43voJY0NWTR
x1W/c76aqc08FZIWeY3RDHfVZnvZCeEIS5nOqGIbVRW3ztwZrFUv9OpT1BiF
lxv9PPa0zSQAaD+VfCWHlmHKNgPsNDYwZH/GePJUYXZkqm5GrdX2K5BBVIa3
9eA5ROdHK/vK6fC71HHcBBf7o6qQr10IqZL4Mx1we4OhYiFvb+q2B05HmG6d
XYtR9csr6GP8a3GhuDsWoN8P8jnGxT7zjSHg2xFLG/h51lhzackPveSgMxiN
aPVXea1XsctUqmnIiWzB0uP45D7fAuQh3ezQ11hMxT0CDXLyxRwVfdndc3hP
W6NoZ5IbPNHO76kIKQ91r9iE2TTQfCs6K6vmrDmMkdlD9Lvu/aoBdwnKnyfN
iCg13/wpYLcedkyZ9Mn101MRr83m826OCGg/2fUBpSpuD+y78J2XTEFMqUyl
IO6BEiJ2U4qV1tuhYpUQVXSG1f6AN6Kzc7rxRaJ4wZC+40wf0sffhtjAISEZ
PXtkM/ZIPCptWPOtkwb5ERxU7Uvi86ooFNlrKh51PLq5fuU09sqX10Em+7YZ
geBXa/SQiiKEZfey0Icgg3ts27ucfOMNWEC3x7A9qnXCdPnklKpSIbLq5Tk2
A8TIDrkWkbw5gxzfh4MNKvt76EJjbza3N5VvdRuKM/r1EMt1ysXz/R8KsX8D
rdtOCWolWNCsTk2xO8u5oUtXTGU0I9927oH4J19VIXzyP9FBf0xGELz35MtY
bgc725O9oUPCuTxwLiRUm5P+WmlCdc4orxoBgTM4NmQbp8SN7P9TUrkMsh94
C8MVYXeH9YMhDTaELFzsQSDTiAh3xhclJHv9DPfGR+tQ2Bv2v5lz8sUWI3qZ
6JA4EDbbO7q9orN+gsKkDdSEP375A50YGPjkDci2emowU28rflTec3Tb/COl
W+na/qglBIid7RkEnxmcYE7XWT4USoAYm2GoJKbzsc7Kewe4kLtKro9rkmxJ
Wl6l+qvWffu7tKrUPv2xHtVcdtzX98wD01HUN8QCoAyp9ajmgbQTtub0c0av
NC63FXOZTNxEb3/3JRPaOEog1C8t9IZEEJ0+r+7rsaXM+bqOXTOQlRyXPQOZ
gCrTsEeygj5FBTxb0q4vGJ8nguChc0onX5jK6sQPYL8ewWfGryTwHdle1GtE
7I5ld7dlpbKobFWDF1TLPBvgtWVqCCTO8R+VhETJYteeIuQ/Y/iFqxxkcW91
FDSxAdlGQYAMvaxYaShqa+Gb4LCyxpOX9t8NBE0Sx9W+sjxzjVx11prvAgrc
aJif7lyMzhnzpJZSpGCLaA9427DdC8Xa26rc0HdXydQJkK8YUt0/MGByjqes
0Dty/sOBEgIfSSSDfPJ6aO+rk0NckOY9ss+JSZctgxRWyciq2YZMYFSOSl3b
wCX1J2+jYdG/C+WdQ3UUNMNsin7YpGIr0T5bT9E0cSlSgXPqHFzPcu3s6xB2
0vCzXQIlc7TOr22pO70oinMGLIzujnTp5euheoEZNfbQHjPddojakNGlsCQz
mPY1V6excbR2smWwf81AgyuumrJovsR9157r50FhgKC8JNrdNPJkPVVDGhGt
YVx8wdveOuheeNV93BVSN09RA/q297AhHuIxipCsM3M2P/fNoGrnshzFmzGt
UidefYKHTu4DniNZMxRV+EIRrzZg3a+l7ThHlB5d1u2l8NexaXzfCfaCx/ZD
T+lSCRy38tZ1AbL0MJaH95WvBq2a1rsNXMFd/TNxxi+XNOa07W8NwGucc3tY
Tfep9Rccbza6edMlWGrp6BfIcK2Wtn8TDMraCXtzX6CpvBVS8cAjz4BEem/R
dmpVk+DEgW/YgXI8+rrBzVv6pJ3YBWgqOQx3+5V+WcfJYyBKN7Ndf+7YItlr
sw+0uvAi/G0W0nmm9Qt8o+QnQ07HtKlCXY2yQ/kyerVlij75dUMgSSk6J+61
7RAkLsHb8wHne5PaW/eSsoSjws/P+RIRY+hpY+cLSrVWMdEUltxmxocQ/N+7
knoL24XHLfR0KySFASxsT3A6bqNF0wCuiaLOy/NO6fyJ8N2n+qJ5PAl27go0
hTV28VDb20chcp0DPBRmbj90fDZX/d3W0dBzLe1Ps6GwGJKd3lpvyBaKrhqS
Kc4Y3lKy1JiqyKXfwSW8benA5PUIAkwA5TGUilxlUFi/OTHIAjA7sduws8uc
TuyQV8O6TkrB077v9OUsIkTkFRRWTkkelEpyiqqyP5uwJloWmYrYMHhbP5Fb
K6xBcCFlpR1npTFImwmVb0vNzOXC1AmkUmxXOKu0R7yan330Hif05aT/yJ8d
jrz4Vdio89ivO9Im0cIOs/Dv89uZK6gOffFg8nMy8nkdCjTiWiugBKas4aJ+
OFWs+f3JzfAchTAl0ogu/LzfTb2feZkRsiGimPLCIiT/C58i96GoauKXFTz/
FzXcUUrkV3VEYlVwTVmn5xLJLrY1ZEPy3Mu1rS2YnUgo0Yx4leI8eJ1uNyFd
hGiLD1yQzj4Ojy0BcB2NrIukVhlOvAmSGlPfFT8Ep0mqQhZJt9EGKlVP226g
gR+VjWKsavmyWrw2neDzDsDc7vgkhlVgEYnGCnsMoraVCRrKcm+XlrpPXPat
jWHbOj+B2Wgh8HYa/ndQcD7Dwv31w3xO/nxKe6IaWGgfVR6v22z6OoeF/99v
U0sFa0GzNKVX+BnEmol7stjxiPZFqsrw1AmQuOYEZEGWcxDeHgNJxaxACS+R
4DS7myCMv4SsAC0lp8GLl0jrbyPUjyKkuVYjrQO5d6LGaCfOXnVMH3JRjHzw
Wi2QKr2N9bAH/ArHj0g3wrzRKTCy2gZxjTPsAVIoA0XVu/1bjWWlqtKfw8g+
CHJyeQSRfru9hDLwReGc3/3RuyGN0+tQ+EBATEFiBEiUDFzUAh9NGn5WM41M
FmzGWNSKAjgMQpqrpun8556YHQDk4cYyWTLjfgJq29YUMpMsgaRogstMEPiZ
wTX2YNgehqL+G2NXq9w29NzjuhHhzOdwO4FOpwWetVGZxasSmVViYum29lbg
/QXc51aTvC/Ltu9xeJ+nqN/idKtyOkDH8O2c+5s+RFFHGkneqLRtUxjPR5fG
cHuGqgG3IdVpe8hxq4mm8cucyBlZ7h4MeuyBp+1y94aUDlGaNjVJfDaZpM8X
1wvsIvEQsYZaSUiqhiYXb5qlMQ9HidMSPS3pTnr/Ng1y4SmARiwKko2fnZ3Z
1mejZ5iSPTw02QR/r7uIRU/0hvuvwTqMW2IxMCuOTEjjr+jcoL3Neg107L8w
O15Q2TudLTYEuOz4E2l7RhNRdo0+ZwvKoP7Tfq+bqR7LIPEax/q9VbABGkET
Wj+LKNoqY+1cxeVJcYQ4VyPKDSlg8UBi6dUHRi5PGuZGdqZGGIlfbCl0co2k
NNBvyuwf/U0AcF8jgsmjwwPYnckgCD+LBVigi/86adI11aTJDkx6aTFInfL+
KOf2jIX987k+kHsB2OkAgLmJYZejs2kcqOnugXxv7iXceUdo18kGOEtG/8kf
juvMACzS3TDzzszOxgT/R1cLGF1L5PUiUo7MJ7OvRKIdxanXo1bovQQPEd5c
xA12gzZlm7tXkZ+EtmfnXqx2uqtYtiNT+TlDqLvbxLjtb/9vbpJ+CRn0jowG
HOQOgFjIzeLQZx1DHD09yGD6k+d2NYhipjArh1pM2fV52+yeGgjYv99aOAtk
4eHA0xUxsxwmrPK8H10LAWhTej3FMuwGSOyf/Ye+U7HU51TpHEy0K923BLFs
tg1wRklRQ5IHHRLzh0/marpwBlNr37o7FaLw0k2A0ni0VlgpCIQLWBAG/reI
VnvAyD6OHPcUFZt8+JKrXWH5KVObx43C5AzbzFjANzlb/dP/E5mV4jpbJw1w
AXbbcqSoh0zKeudVLQoJ89mxPr/in63f6++OLCcwaFexVqzv7NjhuQfy8ugQ
hHUL2K9Kk6i2UZKkcNFdfhoB3mvzksm7BHpWaKiuxgJoN+JigqV6hBx9vX86
XLUKS35DIrsXwy6tLhqcNMp8lDh4oxVWwusmOP2/S5oYsrjPR+C6WbYQXJIN
1HapeKiwnDYcAzlfd9+00P1lDcvFYQGqVDrU7ueZw4+CImy84FOlUFWCvDLV
ZmdpTHdCwMhXE+WYL1AaYpg6Or5zY1Qll/n7pQIo+96QyG7LDQEtn6L7Ge8N
g+bE0Fbsmqb7dMjlX8viYPBP8ByWIgrdAEIPveFktzIIOjyE9UYHtKiyl7EW
ze29UjQCdpKbnTgw2tTah1GEe5VbstLF2TBPA6NwRgaq5K/knv8yiqa7tu90
aFxM3A53R1Jlfrzh67Az1xZGLYH8Ebmjunp9ALYMukKloRa05ig98rPBpLS5
qWIsuBqCZOg6YDVUsFRZwncvHQ7EdX+or+Okd8tLsu1y65zw7N258DL1WYKy
1xrHiutWjHBdRvbMUXEjK4MXwj5jsBsXfV7s3/mk4LJdaePBinjnzpfryEds
vpjqUzDy6uezdzQ9ykk/LmrA+K/5P8pS1ye21BHzP3MsUYIWd3DLqTPDCnpB
t3ipaLXvT+v5KOP50C8SBbq0rs59WCXvuP45WOe4O62rCN7GUHRYybwoRp5s
U+B8R/LwhTc5NI7xx8vBkT64EuEvoNAmvIpctXUkLqCiELAloETP29X3oOtZ
atNfENoOSA2uR/DWMxB3TK3bru7zJARCJAtT0rfAmoLeyfOyUO5MJGCYHZQw
cdbeoKOg5GbQfmKkPdLmPTrI3KDDz1Q+LljsTUbUA9fvuT8G/SlAEoasRY/8
2vmjjGrcLiKeYN1Eyv/VHMi5IhvjiIkIE8yS59OHRWG0LDlov2enXHMNzhTU
IlIni78nZ90APWl84hi782tHgCNbzoYapY1+/by5HuscvGGe8Yt0FPzZRqjN
ax6gDFOrRT8Zx64JyuSl0/V6v2DmeSaGKp2o7c1LSodIKEoKf9D/LjzvZDPo
bWRbxkLuPGjOeDReMLkEiDTFxpko3V5jpws1f1BHjOR1Oo9GUiIOkyAvDhgJ
xcw0DQrh3ukGEAkOguspF2/1c/P9LWQwY/5PVB1KEQaF9DVL/yyIUQKN/eio
CKW2nrjibRm2O/8QkEIoriQnMRMskfl8PJVCvzLip5H9tONdYehuBVrE/Rbl
quC4maKcfNap4Sv3xnA4JvO+0pyssp0gQ1SxEIVlMgXHs7vGevhLVSFbA3Ek
y+WPAHLE2iHnWmqL/p+Gexgy7yBZSpIu0ORZlvVZPvA+DUJWe9gEzw/wbjrP
iRywUNYvXV8bBHyigpvzW/e220Yj9kDsQ+RZkrCCGarsS8myP/mDoL26P+R+
75N32ItuDwAAK0czbBajPHo38AVNLLBmtaIlshmIz4d2We3w6l1ov/gcYrg0
Yw9BJu+RaTa/dPlRiCT4Hghur1TgSc/F8VojnddyNKrwPYwqnhNC5xRSq7Rv
7XbJG3P1yY43YCzFobQ8Ve0IGv/OEcnqoCh0LNnMKHPwS3VT8+0tB4XU0792
BWWizgvaQQ0lMIW21C1H0w1MVHCbAWEXki76x/4zs2d9rymMXgnsgPLXpMdN
pMNoKsUnnFZUaIHmfNK9vJD3z4bhpODkl3l9MDroVrnM1/xEB6RjrMf02Adr
PtchMigURy84zFgt26/kBq50epv6wlZ/WYd61mgUoIcheR+EjEFRjuSBGBj9
LlEf1ZAChJCVucO94/2yBEOPI1x9mZU3Sj1pSPKeLr8cpG+L/piXSd1Qj5Bw
z3/vVPhlZKzPr2ddncDkqEVYWBKV5J/J/Yf1z5To7eXUwD53SaijRNRywmVW
mB3KEsQa8SDfemQ6bLDDmHClKLY8QPNeYwuVBNeTOgafpNDhX6w0ImTtGT58
oZsvRL5Mmi1tDDDtbuCp0lDxIPQgReS4aY7rMy3HSrPGrBdcKHNtwcW7IqPx
hetqRtPVMxEfYfBVrP/MzmEnvtCCDnTtbGf8AzZLLevLIYFcAHPaOtNx68Iw
R056aOtLZIo1ELHchDgmRlRomfhTbIWHDP7eKmFj7+pWwKTQeQBV/tb4ltl+
eDPi79Le4a4AYsc3U4t9HrCwrGwxpBiahoI46VVMx+F6Sz6iroLtn5c0T9g9
+4tNyxdNn4wcMWtZb1HfVREAJtoeSInelsTijlXqNRGc9gkJ5xo9+ucalBVA
YIMvK4jcS/reJ8diuif9YWkiR2500qf80uYm8rnK7x5OTDFRPGfntS29XHwV
VAPZkeLeUAN9Q9UxbCjUyaj3rhqVE3qvDLjOIEXJK25VvdBO5NPdj1CHU6eM
KtON34PV79rq+2YzdSvNn5Hdy02rg73HnIX5cG41cQEemQYyDMACwGw7ex2c
wcLetsMzYHZHvh/DeQO3k6wEdj02/a9Qv/ZQhAXcyWkgMFCKq6hUMzfXEdtE
zD9DRVPoeCceF48NGEOaN+c7HtKeRgNMh93niiwdeZnd9cgfCBm71raHVXyv
g4HuVwiBmrn52vQjZaGnKkZeiA0JyyqRinzA8YL3VheNErgQoEnVkmXUM6tn
5dYopyfHKssU1UJIV1FgcMOCqNMQk0Wqgf002FauQhy/IYzXoZQGSPkztoUI
1D/RA/xHfnoJjqhI/DEao237EgZVBVdjDQljR4jA2QbyYYtQuASo9UqyZbAS
3xWqBLeJYbRVZgHN+Si0A1vCge2hH/XXfwPjOFYPa4i6Ht4lyOhf9idLSV4H
I+3LY1kWqdURpV+IQa8FQJUo7xCt/trSypS4EzL/cUxysZumP8T0QCo6SrOv
Me/8OFYcXIH8SRcHPHxMEViBYjf1hJGOUmYw45CR9Zgt3jpEZf6hl2A/YBLX
VtJKCeGr4V3A/aIZO1X8e1aIVg5D2SdPZoGcrg6LiD03guQvB4meY4Ggd30w
PmvnWeX2uS4gejHl5p9ESWqKQRintTA1+Ao2c2u/djzbir05TS87VpvbLtFG
SPNag0qYdguprCg6REES9K2H+FDEhcJbGIU3t4as42KihNuElNJGQVCXrWm9
GBZaBzSXnsTwfsOmvKQWaIso57eJgd9QrRNeRgLG27H/dUPVE2Thc0ZeZRG3
rlYbFNpahge28WSLfCUt+bFuzKIvjAAkiKzhew0J4+1xYh25Te6Cy/WhIkTA
ZPRab3/nXLZK5K99cSNRcfyXEOkdMa2TggWLL8PzpjFkXQikMGI60ywZsvWY
Zg5orLPpo7EhF8Pk46Tw6+qIGt8UupwPrXY+gVD/q8FSEGgFzteQfItXzKy0
qD/nrL01CCwutRvU64LqGRu8S62wlM2WU/OW56pGHLL8V4UpDt8RSjJN0XLp
ToFKB0m1PU9p6CPBglqjvzozWubth2auFfwJL6lTqnOoSd7Kc+SnuJM8HDiw
S85j+bz9qPLDjLcfX4BajaxA99eMI+8YlxsdgMpeBz7LOEJ902jH/wPxFFbD
kr4NYJbKbeSakY0sASwUf+hOMHs2rV/YB9f25o6vx2CIeTc7xy9qzd2Z0xuH
t1FYQ4U0b6PbRUEU51d4EV4zkT2V8tOHyV+rxtNw7JHeeypXHlzGQ2hkHPnc
UwjvMjuSC1h4GF0+kX46QKBN+pBdHWJVFLRan0N80YIyNpn6YIvNXaor9eH9
NBhdllIV0W4Rlng9HymRr7tzzHboPwV5UvdPciVEs1747Nysf93PuMHudOde
PTbxa1Mzq28Y3YNzBsIOqYwQvmYy0fPNPa7gl7AdMqwHbOzM1iTq3kUk5ZR7
LpIgCRucl9vdcrLfqFmpLG3IXfxVyOU9Y1kHWDU/w07k8+f46pJpdkBq+mGL
vYi3NkEl4+y8KTm+I0NRGnq9DjFZ9yPMsVJGAUhppxYFvnCcXq1XxERhKwiz
2WyqC2YHJRlV2JPHOZA1nMXLgyPu5zfsT1h2ph/m6GkTxq9MUk3NHGZqmAaN
J6mOUmzNgfkPd7j7oCon98gMsj0at2DsHvCo1fNkRhEXHKf467oVhkInFPrM
G9Mlq36nfn7gr+tvpQgtYTxmj8oRmpiYo6Ts6DUuyzn19RlCzg9C/QIlHMuh
gPId5C/Y6OpbSH+UCepc+ibYR0kWoeLW8u2mxDNkBzYWejsLfGnugZoGpWTb
fS2JbUOazMuV/iE9YbTfwZinfX6Csa4X/W46Gw5LtPQVok9pBnUX7NWJsJNX
mSYA+VefewpJ+a9FOAjcPmhr/1m4wDA9B4Re7VyVBX9nTRjwWhcTtWDtgsBt
rGRz0zmAt1BPO9kcqCqTL2kwUKN06bgtai9DWpW3jJ2/qgBvoilF2dBg3QO6
e9pyP64aQjS/RxzVOKJt29XBE4JsRtk/I/BNpTUCwS2PnF8SMctv2WnYn5ZL
GSAVKk6sW9rXawV8I8jFndUS+qlQygQ0+yZd+Nc7d6kOBNFB4uCHnQBcBidU
ygMM+euJMQF1gVIdqCXu2YrFVPlr9+aQBMskR09cMs7hPW6aiWkCv5vNK8vS
rooxtILhu91Pzw3ZOqywMQJ1ORWKbA/bz6rgNf4rkpUYlobA3BocWDAS1sri
hCy0wIPq0n0jPw4jW4LQ8Z/1Wkz4c1+B5ws1zdf3teLHARq+rbSBLDoWLouv
8+WmovqLVu+CEMW5EnvOl5XrpKfU5ztcRtU0b2QQi2e2pMlI/f/bczNsV+ke
fF4zivMw7igvF4ti/kVfzYzXuMdYBVbCn7P7UZW825N/6As/yZD4IY1/TiYh
HLIv/Ltuo08ggGkxSkCXTh3jo3f8lRWc4GGEC5qiWH5WFUSMskEjnkMcGMuf
QdwShXH9OxDTzlB3DITXA2T1lLPcIeUaphjkxUH0Y1f3Jry7IrKA8qSPUjYB
ncp/F+wHCJ3yD5IH65iswZGdrJstt28a4BCD/gniynByEuyighLEADbmAOpu
9wav4p66b/Wz0FB89/WTvv/baU5cGZYqbD0227RbYvxipr/cjDPmQ0KnjwfE
WlAYlKltqMJPtRFOi6qokWVmMC5m+uHSWOAdTFuFUKa14fMkMZJ6egxCGGCs
HBW2LSlQCOyof6Dn4D8RyZ13uhf+gRffgS2lhYtzzImsZdXZQEdGp2/GvPTl
GWYb3NkioGcVV+xlgxM+ECAjbnvoramq8mOJUmOpH3s36HAbyvqiWTA9mtQz
MToKJ8gau82Y5sPHVgJsERSKMLLncddQyIxoMIVTetYAx2Aa8wLlrq77YmpS
mo6oTmvXUkIoF8z5Dpi8PMixCTNSnelZWt7bH7Y9o9pl3B6a2qPQoDR1b+nj
q30vmuBDfQhLE3lWfLwdT0UADcdl8Pym7PMgNvsOKE5yIe7MUB2hKoY6iXqt
j0iNccffhRluIz2AdWaxqUykw8nVxVSrSU0LSBuv2tXOXfCI3cyyAGhWIu6b
awJU0a154DbX7P5f+8M/mPrSBxyMGLLxtXXBrdo/qK1gzNp++jT3GI35ac/W
6iKirULVKLoIttRgnJZ8JjWYxXKNQYr6tGiUiKf2gD0sBBSx0S1deFUVVbVH
XlitY5ADGHgXur+GIe937JGGNCTtooS0/ILa7HG7KGAufHTvnRylTBmT78rT
uX5zKQQkr13D/wS1kyq2mIpCJ44AcajhLrd7WXptokoHUfwPPVJDN+5VpLu9
6/EcM17+GCh7uJvWDH0tVHisZSsPnnT6FMuWMmhRnkXAtwXlfRcceDnFa3dP
BQn//00oUbF0VBgXPnt/WJX5RhklA91pC9ZLCp8LFl3W1VOZZHtaBDW5PCAK
x4DkHZG9qRigigAn3uXkq6/amB+4atM5iYT5I5MFVVLyAry4EEnhEd6TXLjU
iAcdVstKoUApVqJUdxTTZpEXMJlyVsw3zUvAEgl9O5+J0iOjaGKbw33iLmXJ
OTHSRxFfloJJhKMN2E3YhOGkPczd6jXs/MRdtt6prtDcaFWxu2jWN3zIG2sl
U8gXvTM1t6x46QdnVBGg1YQEzZbepoFhUKP6s1ojULIyEc38BgVj2dcPnQg8
FOosvvMmZ7ePJXYnbNkyDih06K0VSJ/GOrTI3/h+uiYOJ49ghfLUJCgiDCXi
SO7lWNXaA+8vBI4Ztl1zFC4utBcZEj4GRHs/r69yWnM81bgp7oiHQL0xoR3J
jeAIzPQddnVhX8u7pqHH/no0uyemenX6LHwV4WLMrjYSZKYFpxxdeBgph/B/
IhKcE/i+K0jv529hlABWCE3qg1u03kkivZFGPk/e4ttMMyE577xrwgEuXBOg
TAGhQmlPJMJ7tk0D3Ad1RcU4N0XwGDTzyrXZCoh49ivjM67CtghNX52EcriD
AiVtXORquZ4b0fsZplhQtA5um46Cl2bMxb0Q65SBIE1dUI/wqQOYLywAgSUQ
fkjpGYvfHVRzUva7BfMTzgzC4qyH4IlyiCyPHK/7ArmCjirlmzefW5GlcCau
62N+CbOyr9raP9/j/sD9QWd++exeglvVanisTnwdsgsE8h3VmxT8giYALN6r
UvXPBtRnlr3TUfJdOiW/DTmCFh2ULSQOzpfvUE5rYY4o5+uVYkskoN3pmr0Q
dets44qxcHFAomG/SYmu0M1Nk7E8kcrvGo7LeQ1YBBZdpSoMu810vyIUuGjO
vxtdbPe3clRHW9mI6trGMbeDYgISNSYD9HKUOqsjc81PKRjDcNaoxhSGj5N/
ApDa/IAxkj3Ru4DW3UwkpneE/0wIo2nPQJO+b4ipjvgCgoPDa9v74bgko5fk
WWFu0EKq48sZz8nwF+9As2pW4ZiRp31rODpCKvu/4qfgazT6LzjOHhJWLjD2
vKsFUVx28YnF4Xx4e/Wc9Lit1tFKY9LFHq5HxN4vL4dJUXTU8k9jYDQYTCkt
wpDKPXmAXAhdqM5i1L9/AVqlf1q6OSSpoabeYnbCQa011EItnOJqlLjWf4Jg
Zq+x9reZlcZCBuqK4jptkYx0Uyu9wZ8OOxWfNMMBTiKPtRR57ShoTtesRsU4
Ffu+cyGP6ODrCDAQp3x+NOdq1Wd7znK2+E5my/sfZukSSpmJaXq64/5YU0Fm
mlpXGQj3B5Ff4JWeh/7XgNNhuz4iB+mnvjcfL0eNY64uAuy8TujfoYlBqmb3
kDlEonEiziKDuGrVMzSGWzLmsmCoizSVITtCi4Or8MdpC64UMvg0Fgmkxjk6
cxucmA+4FGIsXtWdKxTxiIA5o6I46/TmDBS+wh6w4o5In/ZRlFa6N258ZQch
Bp9Jtz7uLQvhkFrTY4TsNkys8D9G07SKbcMqH0snbNpXSvJM2Zpwhq/cUNcx
Pt5IPoFhZ4Y94z8lu5R7wvGaFgO+0c//8Di8JYm/GY0nxwagg0pNy8+kL/lj
2ecGolohu+Yl6wFvADkF9Rc0CdXe6F63KVBqsiAev5JSK0jFNyn5HA76Sydg
Rye++Fk4VorTWFmxKsNybcJsNUX+1RVTn0/1Fd/txKNTQpkUKVF/rktIk3Ls
vAMWNALtTGM5kZ+0k7aRAw+ngYqbrWLSH5dinR+N66HCyAAtBBvqtW4hBjd0
hnWMIlvZ2vhqldGmtaXliLxyYKoL0pWwN+wYqFbcky7EHsdTm2MPkgYzTP1M
jrq+5srfm1+yoTMU2+ZzhtppbzfOwkQq3jZT1HkOOZtxfSZtFBWxbyt02t0A
zY3suvxZXEAM5bjNuuU3lf2rjTZS7s+dNE6Tj/SgirlF33KmSqFQgDU5gJWn
pFxZWXLfU0/Ws7cqVPc3kjSB4la97ed+W50ckcIinBVOa5ML+2aLEKfcmJ3E
MXswn1+2I/PG7zMmsqbJ9x+TZUCNcT6jM8guXX2mvdJrA/eElUt9spZEb1e5
L0utM+NzBuD+sgaH4Ng96OwnGHH9ikgiFcUBXsy4amKEQAdFKoXH90Co/JNr
Y5WPpZwxQohWObzqDDVD9SNe5mhVDJCn01+LqaIsxxd72VunRAV/Q7tzgxGU
3DM+usf0vKDv0Z2+4zCALiqSlAGgNeukg6vYQjoOmUYh+jV5ilxhjE+A0aZY
faUDXbsw1Vn/vgRE8XfiURqIDOoFmdxlvavMiva7jrV5oqNw03kAlZI7XeFI
rjjByXwAecSfMNs0VgXHbuW1SAUW/3Png7t6KoZDyIm0Zt8jhWmlTIRW5VD/
aOiE0ZsY58x7Hm8Xxzu018UIlXR0oyzFb1cHa44H+Deqbd1KS1iIRf5lUjR1
fpFq3PrOdsfJaxk+rqo9rHY9NZOPzmhiEAQ3UXfTQe6YoLTWHdaighuBTBxZ
+/o3hNB01L9eZE1xrkKxQyfqQT1xqrIwYI/1QsIDSrG4mynHIdk+2LCOtRiU
mRgIB5s8oFp0hnj2+LE9/sM5k9VMSthn79Zab5sx74gu1CckrLPcSrQOA43F
Fqf1hfUpYZ4Np6hVg4a7Tfv593XQP+dUmrCmNNrMTtiYnFwuCwCeGpMPPKa8
ZRXCzpMqzXY1nzhwUbyiDRELQbzgAEL1NZ1jIrOf9eZ8EMqb/OgmIcCVuZBk
FFOQ/xnQmfUOu0Txlldhz81LWjOCQTiW4pmVVfwt3gBQJiCK2L8Wi4qYufRj
a7AUTDfBYYq1brvFkYwQ2J0lljwTtklBdaZUrxajH7rI96YOnq9XHOzDWlYE
1b30nUmDUzM+EwfGukTT6ppaF6E6WnQ2CFvhO+amXh+lP9Jbba3Iifux5VMW
xPfTjQLDqCPqTPis4m5Q3hzysfOsajV3iu5p4SmquCf2lkXu+/k9shYvzeH3
SItS+J95UvBMTgDmpss/1O3HSiezJAjCMktRGFaSeIoDTWGY3XMgxKhVvMmf
YBpEnhgBbEwNRnhVmJ+tLpsQOkKFuoikatj4KwwK9HY0/gIhNw3qNSjswWIg
wcohztbcF4Fik00pQnR9SfhMVPTA/z2o7Zb9PtpoROI3gfI8hiEljuio4e7j
vY6eRYJ9iUEyDyPz3CvkA9w+AavVGomGQZWIB+dDjSn/DCzoVkLy7fF/0QCk
VlLjHQt0jqZ7Ia2OlGiOGiuzOEYdNAL7JWkk/mY1VF01wSqjd/GGO0JuYsml
r92bEoBaE4dnAsnYtsd8Itn1aG1tEVCen4abuS6PVj4ms1de/4SKyDKokIKb
QNhFdCfRymEvtqggK1L06m0zlXg+LBuEOt6ao0LR4LOO0RGe3GGD7og37EHX
Psk2fyblzsd9Oub8mAHcBiiU1Mf3PUPOPDltLrQGVpXsVYB4Hbk1x4wZa9eu
uFOmwnQSrTfgT+Uteadz3TYdb9+WjGYjQnXuQ3tfZgvHHzW6vG5USIqW+/uD
6ZzCrEU71iPR1gAQOPOKS+Xqd5MTCvcljq+Xb0K64/iq37S0YWbSKgOiqBln
aKpaAv+fiLvIGSNX7YtkY+AJWa4HtYHX4eWZ8lJP+nVIEdybc4xw6Osu1ndL
0JE/SZ+1z8f6KGvmO/Ooer9XC3hx8pFbV2gKqDFQfhGS8wqjZDEAqLj3sjUg
sVrLmho6fOJMY5J2GqDkvfCadM5RAlJWVKzXrlK9RLEg7cUJoXwb7g72/FHQ
4L0jF3ufJ7oSgC8+c5dFbl/+HtXs6a8QFlSCqaTGEgce0mHHsL23CSaejNpb
YEpb+aEqsYlgSwXAcBQfArVuHnLe7P2BiT097ajj9rvFTyXG1tUQwlsUgPVv
5+qJPcEDkdmvXsJXhXYSAoGDoWO+tPK6BC+oBQYQY85+cIUEArjt+oFiiHeU
8KKR7wf+xYGG3KpjIblzj9SterhYJdMm2UhPz0ceFcLw1K7TZbhNGdKOsnot
kzpDgzj4bl0tZYWbu7NYCXu4eKNZIykjVTQ3UlsKRoeZJUyjphoSJIe5BFfK
FMbudsoHE3uETXxKSa4GKvg9OO02N5Ht+ZJVZBKFMZoneoVodVqlt6ynvCww
OgLiz6x9S/I7ZvmXE+r3rf6kcfP25UgNb32cvn7XFCpWwcNkK8CKBw21Dtu4
xzoxJtQbdNZN7b/06GlvBazTwPqre67MJlo0Z+yii2tKV4XznS/CSfsKW7mp
wSCc48e7J7a5hBLdTapPlZgItolFCe1gr5CECCwvLLhUKKDVRb6bJZrf50Uv
eTha+NVKeEiE46p5iJQzWg0LIG3MyVWlpfrbRRsBpJ9WhI3ZEYwCjzIJxzKe
DG7pwKABueb2IPHoZiFdXQ2DiExG2XQHO/upxE1NQMwYcrbQ1A4c1QoIslv4
d7X8G3W/+gfYcPrXjsT/mjaWWhhog4DAZUqQYtdEWcWmGN04inlPKlBZWD6O
f/TaQhVs5xH/ZUd4owgryOsrW9OjS8VXhEH8+3+yoHzG2tvPU16pigKOSwzz
b7mVZNWlu3b6sEuomAOmpskCfjvTLWZby3sw5Epk1K1yP/T7TYFuJr5UPOG6
gtUzV/a3LOfiPOg1fOWxZiBmkU0EaYPOXbQKgMhDlGBAmyZZ/XQFpPugFFk8
wppGZZzweFHaaK1BlGdzuGNE+QLGPmqY6FLJEdTiFfkfTPmXeEIG20vcjDuu
O19MD3B6X5oUOV/sc9fZa5pExUYh9MnYwQho1jQY44A8ROyuuFRQrtDH5DOu
zYrkwoJuaJxd3Y0Y95oTcrpiavIocuQbgyGWSMB3tU3nTXw3vMVBMAc78ZwC
4EpULXwUzONi09pMjUidFePGuh/+VRpVhpLk2hFo3RSz1ZJvVd4o3duYuigM
j5xkuR/hu2akYX8gHZNCh7cTOs6Js6AbdJ5uopr3qxTWs0RevnxdX2S7kfEv
wXR+wd/F0oNJXeyDzdfdu3HNrQwvTXAD/eZGjkGX6428ILYhu3g1qZ8TUX/y
99bcHgZJHz3AN20Foqd/bE6PsBAkyJLgIZ6/BNogJDJUx/lT0TqrKAzYJKHx
p4MabIm8tI46o2v6JayAdnYxjmwoH5VAlWE5fn9t9QYJ4/tZ30LZ/3nteUQj
BTvYJBR5JWtp6577jBkHdVGW2u4qxFDlVV0bQjSJrTl7HTG5D4HV18xjhevf
JvB9GzY1RWFzMxKmy2hNsnoCdKzNZH+RT5vQ5Q0xQOBDAIkQ7VQnT+4A830o
B6X9D5E78v/Roe/Un7sim2cW+MQrwhMsgP7DCETg7lTs/KefBNFZM2VjDn8a
EgCP0a2/C6TRp7N3G0vtmHovwIQxdATv7VdAvuF9QyyFNt9pgOKpgU0GjZ5f
1x85Ko0jrJFMlAYX1JZWAAKke60qkFrql3Gu6wI5w5+l/NGxpX7ujG2t57vR
l9bkG7JlwjFoSUKI5ljm23yfFUMHIkzfOCSTdO2HGG85CSrACqakT69GyvOl
/V/hTcJtz1pFBwt5zGlYGVaLJxkoPvWucjJaBiS2UKukUme3Va4HfQvQGuOm
SX9zVRpsGiVjizLp9hYKTTm5Msnz463xaM7yzsWk9Tchf8kBhZLoU84zXdeE
qC3rkExbQTexFvvvwPOVRSgFipZmamONLE0pHSEMxodLp2DEo6Up7twXJ6kJ
jr1TtGv/o3KrHi9MKStbIZj94xWsSTDwdeegMUGbQtxTebq/DKxBj8kzfTXU
fGFCPzwmMnvpGVmOc2VXs0MbRPZjUg6+uxAMMQTcKdrB5mn8m1PjoTJLy+cm
cyGv7ybwQWXILVnqIB+GFZfxNEs0hRgY5X2h+PN+a4jZSzTed3nQQAWGOCd5
641t/DdHFAuTqjtXJZlI+fVzYIlzbOXH+a6JRbZEoLrhgPXN6q4LoCqFCw6f
bWVoPRCuZEikujnhfTM+PsEIZrya8Y/AZ71zBr0IPz4Nyxd5wwyFEwGcyock
hmQu/uVjTvNdxFQMNaECGcwclvfE+t8NFjTn356GIB4cMK+t4BB5HO8Zbue6
dPxjHNbE8p7gVgkcCngNWxnVjP2057bbi/dU+e/egOoUPf7bFJ/oQzsnXqND
x4wr2j7tSRoAzLiCLbmu/gUPbrhpU/N7FXQW3qXSO1QljmLV6dM1utWW0Rqv
N/M5liv6XFN8O5ZACNq2Ak4rrO5iKAiZQBJKw+U9F97RozaJAy5GBYaRQTSa
WMkse4eOiar635P8kuZyvOkAfQ2ZhYp9KGg4ltRfrsGrco/nzz4VjDywVVqs
FZSXbeOEHPX2zcpzannmtL6zwmc99Qlthp/K0A0NDb4QE51hhrjXVdVgT5X3
NWGTmLbBtrOAUqOh+26MjpGZHe+mtf192CtA8e626jKEMEaklSlolxBm72GD
MutItG9vfCggii4AgMTmJMfylMYEACLWe6E8Q4x3QtJTmhIWeJP95LdIhmKM
FA/7p1KuXVNPOe2lKPDdCu0xXXFgqlgB5bYMVKc/lM+bkZ2OX17xQD0DfX+D
x8Ze+HnL+V/NcClm2Hq2Ol+co+GrItGnBE7Ez8t997HZMjrJWfB8jdnyxO61
4o+rxadnhPfSm5NBmCgrOpZ+ssZOtprGnAFUAKWXV6vVvTLcBZPD+/J6Dn75
t3BFO9i8c/qGKc69uM/j4T8LTStehmsieaAJtwYbunad/nBGCw2Wi6MDXXvL
6ZMDHKBnm4Q1InBnV0zqbiKOqIaqRm3mfI+o1WOV3YgkWgsX1QxX/NiQll9f
fSjDXiKiFJPvn6QN6/HABbNRnXYYLm4sVaQV85pt5jQugOEvMBOFjrBXsKic
RDpQOo1KYRiqQpEPNCBBdWIL/5DDNAGp4GnlqPkxPR0vc8pqJKzv6pWjiTB3
Xr/vZvOfd/39jS8apwPwqmYEBiCCTzXjU7yoyYLpzHg0lLCVuy60z3G5leRP
5a3IikLZ1QSGj9UI8vqYp9r1gbwj4Q/TbBLmMiWqu9Um6+UVd5xB92ig7oR7
F+nxdBga4A3qVziwALXkX7tVfxIbP/8Gw2tU29kPJ66iA6PqbFCHrz3gQpPg
c/O3fbzASNhV7UaPmbtmQ6rwiIYz8qnse1aZWzLdhhAtztf3S+uoKTdeCH3/
mLJGWY0963z+nIcC8li9sj7K2X33vKedsiGTwCQNsnvGOu2CyCwyIep7he3/
MBPvJSCwmP8xIip0TWKLZV0fT34Cghnd/e0L25bK/VQdX7SKpAI+PmLW0F55
MG7D0vXJrfmdeIMAJuCm6y19p5fxX5ZhWMWvwTi6Zcj0Wj6QDcBfI1ZY5u1g
m6GI/G34Q79Y1w0OT4F1WtIiLoGaMvMCEdnm4YvZQ+pwuo3wQtmPq02Gb5zT
5fI6bIeVeHSxWQVxRk6lsw9v5706c+cV6iMnCp8z73bEoLAImxLvO9ibxH3G
3eg/zJrNcKJ9OvrFiotsQerpHu1JK57iUkYOt2Q6KZjNdqZEVGnqwIL74ea4
sIQ3QAsSF63iDe7xvOnyFYFhT6KPFURexL/rof8m4KBPyw/ckG5+jrRTSBSj
5unP0Sr1WsWSFCvJ/02myQnbNoF3LndKZwz//gcdp69p1tgbKE5sHqT0XyyL
YkTZJWgZcBH7+QClHBRD4zsj4kIH5WIIXzppnt1/XUuvGU0jjSqFtcYRUrWi
JkASqoVTFpn9FXK9HhBFGhMOU+xCD/a1UWikEB+DpWrS3jGambxUw9SBqCCP
mCwh5NFmsi5+rNdVpcv1Sf12AJ4atkA0kVwyp4QngW3hYl3ZGKDMZImazzyI
vJgIxjBJ3YV8Gfx9ngR8nvZJa1q6mSfGUss++KwE9euUezEt3e5MdAB6K6KU
Oyddoke7ZzZ9yYL3E6MPufEI+YFxNloeZruNGaKH9sihKJy3YPXhPYzCq/t1
rtBCGUNXyHucfOIKAKMjuIswAwx0aS7rmvYGJfEE/kzJm0Mf3Y+8BqryrUsY
RwKxRNURHAboiWfNtEwPVt6IEN3+6wUxPtM/J4TOm/NpGSaOmsJ7A6YcWl0X
Dufc39byncq+yqWMf6KIOGsfESxgQk7Iv0X+wr0oCN+TfzWh0Nd26WfpQhhm
546r/kId/vIHr92BRWisrB66ApYb+Iu0WdLwl43kgcBxN27Pl/7mlnbH1p+Z
z4cMj4PSnH3Ow54um0YDVaeFqcbry3SNGbVFlzS3lGBdJt1sxXbe9ehqAcbm
d2Ofv9/jdf3flMsWREtX0mZ53hFGurg7WCA6pjat7EO1YzkXdAOnJp30a32M
xQTQkE26EQesgT2HboyamkEh6oUI1ZFFFVE0cmllsT5L6tW5k8M44RAMH94e
ucHvcmYxaV0tC862bd/wBXaSPCCRa4VOeyDBpzH+rhDW5JAGEhKNANPSGSEJ
1dOm1oYxTwORfweFyHkFWzIEybCh7PjcPz2I2IEqB4PsmND93oOmJEdNm0HJ
v2LXBWTW4o1JHWKSbRtVy6R40V9OTrFcGUxI2ImRbrteKQ1K9NUH8qNz2/XK
OtM2wKztfJGuzdd0H95zvZn1HGV8Prq3qU3ZT4ndAzrrVxZY59FIjpq92Ar4
jqxQ2lY6V847x6hkJ/E7qnbLh4CEMkgn9WkHJ4Ro6BfPYmVMAZsTCWS2GRZj
DyBMGeouLUg29Mzkv3X51kBpK5GNqPKyWeiLopUwSNJGTZflaxj4EBYHzI6W
te9xQEM+EtlwW+8QlBtSRN9gSHKS0CndknvWTr9mRUNUVyPKSJlw6Z7TBd9r
ifP1xW7/FWBLWKqs4fFVix5P48+5tz5O+iVLHWFi504KzawDG6DcGvp4iq6s
5pi6agK1REq+6phcfqR5dso1jGWJymGkoYiY6NUMAogYe50lnmgGcO8c9Hry
+5OSvKuoJUXlZgJDiNiF90tnZP4e+8rMhxpnA0qJDSOkTH8H1kYvCNkdyPXW
tOoNfpUYq+Oxj/0EgXKdteYop8Vt0J4Ww/i28yFXcfCIAqqZUhnROh+bqnf/
76WqSRQ6gvTGLUI5mFVVLyZ5xvQWNEbU1fgeGYdLKZyW5FiSOU1IANfWc+Ge
OkiAxTWEdrA0u2TPSLIq100SXMUJQWJ6xK+GzHt0yRiamaXcGTgnlp4q+ux/
quGVLqh4HltJ7BUoRUgEokLy6RlWEz5kF4rRs+KD0pIfgfx3bmLoyNJiDnWn
l0hgbfNOgREWIzrQtJBl/YY/EgT43l9maiQqLAOE6q2HmnivibXFUJEX10pI
znBFkT2Xy9uMDtF/droFb6YlIlJf5HMAKJG5NYVioGVce/9nzyh9j3BRo51S
FEWSo11s5MD9GEG7F6zlhSXYZVhtEM0dU+dcKyP0uJobOUCkNR3Wmry5nfUM
6eU+u0LUelMm0WX+HPcTCfTr7NtDLb0oTg0Fi8XQUbCPe/XZQzxOd/wWL6IV
NEhHJ8VfMSQPf5KfCwFsx1dp8okiB4Df5mZtZ0nFOIR4EXNIZqr/fb3cK+kd
t6UKZdPY3ZtVZWn29SXRyeT/t9bMESfk6JY8gTIebJto9D0JCNckg7y7p2QK
ivKs99XbFAQxbhZUkbWDQlqTRytIQfcn+/ddk2JVKmMIl7H0hTW/frtQ8v8E
FTSE5rMl7zvO2ZvY9Bvv8XPtGt5JkRoq+hNqUbPtcrxhnMm2DOk2LSF1qj85
JHxOhirwyCORzNhfJ1u+G/w4TvO8DSvzd0knju09ZiUJivNJI5YMxV48WAXA
vuX7TApFisaAL8TRK/qBCFQ79P/oThDEmPi9YZgIS1hJzXBKmbArC2wNmnhz
w+brgJhpCVSkKg8/GHCP357VqX06b2Ir63L/pp2GfnqJtilBzi4LFdtGbKxv
I7RqcT50nIgKt5dQqxIGQGjTADaw8XVEV1otaThgJg1qKijy75Va7JvvYyYT
DpiskyVmf2O1h69kH4y6F42F3w/05mjaJIgaRVOWaC0QodsA46gg3tVF6qLH
u4LI15rbtpV13HgYaAtxW+K8/x4AYC6zo1Z3WPtCtYKZ0UYnhTb2W2LiUfdW
2IPnTWIRJ4XyK+gDg2zsMXtRDylYZMFoSOOZRheBycXOE4FM3tatI/XFinHW
LYY4hUTt5/X9ZE+Bg/ip6VcCxkt59nJIdhGCFmPaAY8lHmGUNXrvLXw5UEUv
w7pqlvSbiw/apysOWTdHs3tR6vgPteyxSy5yzT5DPbDNrk+uTdZmEXF9omCZ
QA+ZX1OyYTmIRwbHnStLVClBAO6Ou23rGOOxmj3LMuLwlpvCHXF7561uD+8a
udETyHl+m3ImHavaqn7N1Lps23HR7K33Dh+pNmxGb+Yx26dE6vbNcTBgIqGQ
qJw+DJD8iedqsj8kJcQ0AXLh8Sa03lO1nTaJA0xNvh22/PHut91k9ORHeZaV
SZFqpYLsNs+vFewVw1SbzCXeIXExsSKFBSOiT+DvlfiKLqBCeVw03QIrneKu
uU9DRa7qvh5bhWojnJlkA/R4G70sl8lUqqsGYduGMBRQEVWtZDAh32AwTIQ4
HIdujzBTEfNs7codwpLxHBPMiiLrLATclo9didOQq8OFM/5k7GC0ZLIaO3sR
S5M+gTV6r++Rgb9MEAxakdm7fcqe5w1fGDKqLb2FNcacoV4Utv6AbdcuDuCp
LWfmmQ5cMWKp2NpBnvEH4azCYGbdJcgaw2TDbG+yswY6hEdWI6GJSO/a8t9V
D6Mu9dc4J5uK5tCKlGMoZZFhM+ACj1tZlzYABipgU/uo0rXW6nqlTvCN632S
qA4E/yVHibJI84Z/yykRLq2jiNXn132NcYGzuPli2X75vTCDl1DNP/zyTvE7
SapUZ02NC26nHcd2c6txIzY5LJ+I1uuTtpHEn4bPgqIBlWC87kTeN9yjCTym
Ze/5KdVlooSwXOsulh23WBNismm5FEYYq1UDTeZB5GHLoaEmU3+OEMYegX1/
rh/ubEYK8q9pfDtQZb5FDNOLrzw9lHVWAK4N3sVwzKLATpvamA9ZcfcIh366
KUwkHbtjYzTumVgcPp8IsbR8MU5A5LRQIU4F58ALRPt/qo6vWdkNyXXVdH4g
X55uaHKjh/9MeBhy7Mcl10GKutqThpY2GLl3jZzUXgsiX5D5LNfqwMFQOTHi
0QO4WIQOOjXsN5cDszGuTiY2wWp8+rJZ/HvJjeI7Kw8uThP1jGTeV+EVaoqA
ENl4UggMb9ok8gGqq8nA8h7Xt18lCoungZK2cBR3IIenIq8tmN8CJB8Q1i0+
jz2rAero2TzXpOtHuF95PqM5/3nS5lw1U8YgIJTK4ouGKoOjRRH7w7xYqrQe
AXaiuQfHZOHoONDuSRisY/onVZnl64sPDWjYZwsVtobbgAav9am9XOclG6cY
bOgXLZ+ZG6KQJGm4uQ+wHlAtqgk3o6vDLzyo6BIaMFxZAbLZbhatsWc7UEZg
X+k+lIgcej9Bwz7ZSMQuaGUReBgjL/3ShNs5BdjZVX9Jn9SeNy2mTRzNJQy+
oTD2ASQGvTJeL9I8TkB4XSGKwog2bKXuLhpzW5TslN7VikKfZX1/HNTJEkm6
S8Zu2SIOQYiHzR93U8qWxFcpxGeY4tQnu1fmQO9jK15k8acNWfHLYhfAw0/L
Yet0HU00hmqjcKMAgKrl6cATUFA1Xznwa5oZL4MP4XkneREwUdWxlGBU10Ha
W5g7lCHi0i58b0hfzwASvm8GdQz9rqkkn4ec2HT2LVq5488ncLJ2AxglwRVu
maVzMhM+k5GewAtlJT9Im2gn8XGMkyTm04wOa3C6YJYNGKNP5HYiC6mA+nXC
GA/8lbXX5vvNTpZfMl5s9Wbq86q9ZrYbHh0EwfCgjuwzJUDnt4p71pORp4rq
QJUdbYUGtmWE1R3Vt8FTUwge6jK41Ezb+98fzji1H/36YWTKOHRLpvhyUZ66
jTkeGr1fkkmrFwewmyPF2haWEltpV6pPxTf8QoPfqIUV31qVnLnu6a70D7Ag
jv1XamB4LvsR75n0WZ0Mk/+U+3tOddi689fgAxsBJM15NREYMpS0W/9kzOue
6VuB2DSCHkiqTgLj473NE3zW5xggKWkS5u1CkkD48xD0NGczxLsu5nDNxTWh
3ay7WQH7siB7JrPSQ/XSG2f7Nbo41y+wQ9edtbgR1ED9Q1v/jHfKUsnRwHXa
8NzVkXZz5IK3wC5zXPXywcNc7BvnV10D2Xfwy0Vp6alBr677941lvKhNZF2y
GJnk6K0VKCFWBzAYj/Lzu36ep2ISvom7K69m+OsVAKzyB3hrryyh6AQlZU0s
zagBFJGTodS9jLzoj3AGUJ5aVTn1HlG/gmLNWewbwCneYGiuQyD8Un3Ao+d9
tyuQl9zUlRmVbBkL2R+kWWrsisKBtvrE4wx1c4l2KS7CSysJbp5WuXfu3muO
oWQFWvyPdUi67nTFcOQ5KX97E/ASaQueVGpYpSa0wcywVVu+zYuz6bO7doRj
/kY2oyhXDlzZrQghV5sXxagZpkeDRE0mdOtVoNtSs1Q11y5bR2A8bewdVzQt
Uq8ihdo63ktDb+/xMg6Wj0KcpJhPRftq959mTDoyQfiUlSVqUYRH3mBqYkYa
fD0vyZdjP0DeoRm4zNe2y+486kPlxYgLLn948lh3DUSi1kW/LwBGskRleo5W
2vYDiZZKIPs/iy8/0uLj6OIl44j8/TY3QDz0ymGlK7Gm4I02P7a71JyUvokU
t9wZlBoCdcm2LKcLZME2O+5wiji40mdF8yZuwZhH67t6KySF5UonPktFYhLc
PRUBpoSqOU8IZBMX4TtDdbp3yjtawQhMMyZpEDmoAZ4OQIut+qFblLDynqCW
PWFS1ydzk//kYBOt7qWmv8YSQ+oVNr/Af9gth90rDVOuX7BzN/8uIHaiBZot
GCuTQEh8knSlAhREfmcfinepwnGiV+R4ZO7mTNj3WJi/mufdpw12SQWj/W4j
kPHnVTnRlo9Q7gxHDgk1JN+T+1/Ojuqggj8kWAOjXBZOtQZiL4aplNUfJYkW
/O2GNva/zVe2DyFsedi+nDUg9r7N6YAzOFWf7PKiy41LRwMi9l3wulTnO1AY
YpcTThe5yVWQN+kRszmdywh0xR313U3cHav1tiFL3gVAaVxBn4Scree7H9o8
e07RwswNLqjmJRnUnpjfbAa+wRppdYd1ZvPvd+lWSVF/mSNtmi1GC7ElgRdU
PlyH1FNgVYNpgoxRLnSf4r5Q3MsJruRTlR1PQcEuVX54YoMaatiFz9jJfcGY
wKeWceV/2eOxTw2dJug61ItSCv219o+fnmLnTFY92oRc+/08Hvq9JrrQ/siV
v0osmoOineCcwPbLu1yWlwAlN2f14R5eP2T2EATiSCJ6GEMN6SEFCdwNSt+F
++IB4ZU+VeisRglnPtlN2FvRYNLMF41cLDWSk0fKbxg43F/w2/Yr3LS161M2
1pcsvg7biS5GJoolJ95Oc8RjZiNi+yYwPCxsERz352JQ1Ai0BMcZjwX1RLdi
041XMQ7OwQLXkpXI0sODajvNRg9HxNf5BmnD+7m3g8ldSBZi0u6Vt9tueu5E
XF/B3/v9FfvityPd41fCh7T9KG+rmRaC9qcAhjhX4K9nwoR2V75mS5++KXHT
Bue8XiBF4pkuzZuRn5FmnpvM80d1eReVErETlrLCietizMcEvUIW1tAS5CD6
RTbfH+0QJajGF4BYhNgUuUaN0KFbt8BnQj3rrMyl4xshiqBJXeDSAthDWnm4
UJcfCvc484lAc1lFy+iIEWiVJOkQxYUsrCExHEZng7DozPeqwt1xJwJzeLsi
vHqZu6bPRhcvsUdBl6w+xMaqlWDY19ILhWV2PlIofUklrlRlSmz/eI4ev7At
fj/uD42xzbc0JEGYXgOXWBDtFqydEm1RU1dXIrTnqlOC6nbUHvQuUjBwP/oY
6sPsbvte1Rs5K1phflnffDxoO3i1u+0oR2hGk+fvtqa9bhMPHps00qBxYUTV
qZwfzE5R19B/eVLbtyIF6MPaxZLV5SKQWSnD6RnLUobUkqC/FsWorIcF+/qT
FKojecYwASatSC46kYqcMyg6I1lAoh/gAx6ItgPTzLp9YAc0PkrTgHWy1AqE
I458XHExJNXnRdRT1/Mt2BGy643xBAauzAIZQjYMWeL3RNjiGFEdxPwT+Ule
KXntouaxAM71kjgJzJif+Tjul6EjPklr401u+cZNUI31hz+PuUBluhugyL73
C3ia5AJaDSUNSNZ0Q5IRBjwJtnh615X/W0c37midEGmE4AzuZ8YnEM3Simab
eGoYYmHg0mHPS0ZltmUMo7PO945BracVI0amo2LyxeSd4OtuKIe07O/QhP+Z
8Vly51yUi3ogd5PiiNiJoaBIAip3WEXM0wX8AIVxe/YR1s7umpd9WgBfRQu0
eHl1/LksspiP8MqsMfyMgQnD0EG8gaS0xG67gpPNtw4YuC4b7gYTKPEW3ho6
S3XEa81jFmGO2qR6b1jy3uB5ZIl3U/tN9wVn0jMSIYim8W6BQbW1Ym5vyJWF
hmg2ChHiK3zxncw/lckLwF8IQERw6Q3LLSZPbyW/E+SHgubZI5HOzt13kffL
gaGwtaSaTwDL9zUiRqJHL/oXBwnB1ATxVsL3tDAtoajMz14D7LIoeqagmOa3
fDSY1NYaQd7QW+kEJbfGwNf/b2O7EshObbCDgNFU5Sq5RUGhEKF2KgxrS/Ys
QdOF8lpauKxEtuo4hpXbhhXdzmy+hj53MTN6t0lFSoG2ehEDFrwAtXLKxsXa
7q9/HR4u/DJpasFHCBHxUb6x6XISiub3/0V5r4STppR5vmNlSiIRLcWompAL
2buACF0pcKTnCgLn23KvfsTEr/x3rbU8Tc2AYiDnlFAVd+SNHWPyzXqmFrA8
9tHitkGJ4/vSGxkDVtPFlLhhYxF5ZiLHZxNvgNKu53RZWClrwVl8b5QE0LTe
F9CPvyJmv1AjacRbo6j8wmoEv8fFbQ/jIdvWLRfnE3fLg5J/k5CqvRYD/Q5e
n6Vm48t0uxVJPUEqsvLUfgGPRvV55fw3bUPqO7rmp/3dTuiA+YX6ygnTpi6Z
prGcCEd1B1gYoHr7/D6CFDC6nmA/0qo77jgo+czHY4lpkAeOkBcr1iPmXMQE
xytP7ZodAqObU/2MNoHNbKNAEAMtDyT2oqmcB2gdF8A0c8mlmRalze+s9ZsM
WJh8/dxL7GbmLYBkg0CQn1vFfKZzWJElCuDCGo1rcmZDfGpn54voi6WTp1CP
G1p/wA6junAinyBovwfl+uX0drETBaGANIeYElGX3EMBrFCp9sCKxn99iAL0
AkHmqMpnS7y5pB5SkCaV5SV5ercIK3w/W6rqjWB+CPBENXWac0j4C4gtLU1g
GWRNACEtqaa1L9qZqeD5fd+gTfuKF1CtXOebDANblz1MC3krW5O+t+s11S3v
aq5J+OSQyUHg2nskjFGYIdpBJThmNr2UjAqhh1Q3o379b8r/ERFHx3cIO9ic
+MgceEzq38+8zeGe94yR1a4Nw6r75q415Yen6iRQZfx7mtIXlmiHejAxgt11
mDPtMpWJeme1zmDZW9mcKedAphAArIgXBmYhHBw4E9srjArX9CNFSFUQsIoi
+mdopvIvfobQl5xNcfXL8+vINC3Cr/UHNV3QJZgfh2DB3BbjWoPj2Vik59qT
IVxGgrorkoM2ezDnsBikp67RnA88SzMRJMcv06B/JjHwN4P8KGymdxlQMMJY
ujOxJblZi+z2ExsTsRRrF5gvJi5jN0QMFKy05ceV+gk0DXKdCUCwScEwf2m1
MxB8i1dC+nzaZFBIjtOZ1Fo+S/2TZoWpO+r2QJ2nLNIHHw3JLJRMO8bLRKyY
l4Wcjn3fAMLvFcpsyv8bZJxdfdKtZXREeqq4++qCCOwHoUFl3cwGbsaQ7m4s
zbk3ceo9tJannNKJ0cMUc9/Ss5sdk5puiTvdrQJ51+DdoG8PEueEHGxL+S6o
rVlEa8oYYzT7xfZ8NrwxtajDJbIWz59sm5M9oJ3AshNR7YMuBvWeKKLExibg
ifr+Q/Fz46lUsOP6QaD7UmFutaV9z5FABeajNZs86igH1ZsDmjiBEWknpWwo
xm/kIHVxVeXHaKn9+LzyrwwPfaHcD2PvOTG2RqNBQ9Fnx2TXc4gLgLU2H8wp
LHPDgi2LDRRrAROhzFZ0UmASBRrTCKNOU0/4MP/vfhtypD8f32AV6lH+VsGi
3eX4eEw+0sNZbJG/dsXDjEds5asCDKl2MdJLFXsr+wFTvdh6XefeuhPf+qjt
sUdMrGQK9pZ3XP/Bof9IZHwenmKHQZNziMvNd7ne5czafff2HnllMwkahE/U
LmKz80vRA6YYMdFC+lCTPXW0Pn3vMt94yOJR16qQBm2dPueWcQPp9CG5VAH1
3DmMEYzjsGrepo8TADoFv31N6nN8hRwL1fAFsSLSYa75O6uUBuKHPXiqVzHQ
kZYTwBAsvducEIBhOAGYN66hvo1jdqB9UlaJqPCfSaqzmNICOQOXuxwd8uDf
7RqFhoMiiuvvsLOP3AmnF5T0VfAkAjNIXZlXGqgtg9fCON+n/21bSaGSdHIl
ooC6+HhrNLVx/SlFY9pXYJRXlyCG5uKwtMod3OfZkxN5n7UAnXiuZWlQAsvY
nrZoTX2uW0rF/8oPFR3VXwhH4HMmlFhT6UbLwW484fSgb6N9tK1eBhPp1v1t
SrJ6FnLeNgAgU/mOjh19wJgs5aFdroEhSFvvSZ79TnQ/F7Pg/yd532cGMVZC
YJ9C2jEcwCU2bUv40jeyVfHwoVqkOC74UOsi4VC8wrIgARvbXwchUqkXRwaW
zzh0SWw9791GDFNrvIE8C0gjBL16GuS563S71ETN9B0g3sO8mXCxoE7zldnP
aQGfcYf30LzZH5VqhrPqdKs1PT+bgFkmtk9jW/sDnzjpuZIsP1oLN34pKMmr
cJdp8IWwbBBlLzGUchZIbTv5nF/qVVRN4hcK73JmXbjdCnLgk2+hi86tWXs2
64IbVPiu2NyAuuF77zJPN+y9cyyUIDlnE7+nQkTP7NgzhR8NZhm690R/QNiV
1eDQt7Y6pTuZy5AjokzXHQXW2IVh8wpwDxZnjjcSpjIt8ar02I2xgjtom5a6
2UylDh8cl5HMgLA0JD/vHJZkdanVI2oPzusQFJDrbSpQDdzOkrQ7tWg440+Q
WWEigglL/ky1kLLdEgCliqOSmNWoLjZbOBblcnMSKlJtFvnjyb9imoPo+uyL
crJFhbgRI+E0dk8JCVCbH7qg1CA8klKzbm2gJo+9koZLgC2F7QxXuK3LMIsa
PO/cI/OuLJskZ/HeJ5+Elmn8BiIjJ1hIvi/HWHdE10mF76wlyUXQL3wPnq7k
OFxW9tTJskQl70APO2cQ5f3UMPH11yaFsJET5FaoLPqT3fTm+dFScEZrbD2g
gdMsJCzkzNxnwns8+5RXgaxjQ1UW2hBsgWwszVOEDHaxj5YjyGlFdZmRjhg+
2hlBhlPkik4+fmJjVu0nQJWHPta7JaPDl6ts6WJoioCYe5KCxYg5D1VYn61y
yOB6awe/Ub+9TW+FwmZfWRbkQiyoOZq31w1jpIgARbpNi3Vo9ubNPdehUNu9
/CplGWe7xrY50AF5dQaEV+6NleA+zcNTBkDEFe6vi/NKa72T2Ki6A/eKNoYw
lGm6P1RDMRmUwLL1l6RGm0ZzNP3XUDYgdi8sKmZpfXYzaFgugQ88k5h2QsF1
LG3m4pJ2SaSA6bnGOMNlIeOFitDjqKHQubNnP73PjFJ1aA2VlwK37LGLqw8r
j4O/HwQibzrI4jJW5rfAuwjUfEkMbXpjfqf3eQ/+J054YYO+9P9Pm4NGbfEh
T5DOnw9/h//nfMPwNG2R/ZB/buprcbi70rm0S1E2PuoCxC/4Y6ai896huk1j
apjancupNxdKqY9x6QLzCH0cmwoMZz3Q/ivK+zSPUUgHwv+JQqM0f7jzw+w8
3jvEtYzJK1idO7aFwWZQs3g4YMJSL1DA0AIHQ7A7m11koeHZ3xI6EVJYTx4A
14MiatpoqulD2m/LHpYKgQWm3ZIwNV0TDNZq7eWRcqmGJrACJ0wEF2jE7zOL
WnBffZorNXYNyb9Yc1Att3S2sarTL2RwSFhdQO0EXES2+L5tt58bGKQPHJud
obKIYUHqoInod+XUPpfHMBuyyCEw0VbAWk1SMkMVeGXXaO9lEli+l2HdyDvF
ANzxgLiHcgy2M4Xu8wyoG4bjIxzaz+FwNF9RGpWM2Xkl/fjoL78qo5k2ESDd
WtMAG3EQpwYc43nES6O8MgvDSCcU8RnAZe8DmHT5YoZPNPGzu2KoQEWPTwql
owEwVxykTHS8CxuZyabnlvz+qDgbCpzXJ4V3G9l7eTg4BBtMZUnoWqEIABRN
qiaB+iHahksuVbmarOKqglio2S1HrPf9ZLzSRT+1KNOJAhpFtoZvbP/WMK4r
P/cnpdF3Q1MokDyVw5Aial/UKkPmGQPFQsx0Mspe7A+X+PdEFQ605qlz4QLy
QJs54hxWwdTDH6jmpsrhI8knWOwuoZVzOeKMtGHPsfi5MRMtKbqO01wztIcT
kFYKI/+1Oo2D8avFwobJ+lGdZfQL+BqZXUuO0RmuO7Zcg9ezpEdOVCAlfGfi
ZrRKh4PKOiZ8wQqVpteOr/6AmNmsJv0twIn0jNHZVBocZfXTqNdI1nlbqWl+
AbivS3UcjSM7y6Psd4Pzz3AXDdD37SkGBfc8dbXeqOc9YZV6jAgEMT8Q3zlt
0xpMgIhyQC0qtlmOhuTqQpPc9zln7RV+vbudtGgfoqa6Z1kN5Eb91JnzLZAJ
X2E5T7WXk/sZlDode4XOR3kr2+5B3G6Ri+yXceeoeGbRi4mY1pV7jG/UmE2l
7z+ATnYVCrldhgppcC4zq2f2j+iBjVhVZSM+JM6uu7eHuyfcmiN7hFGHqZ4A
2m+icnEgqYrUN4LBWtYuNys50PrnxZQlEJ7reaDActDANAVSY493gk9RcD+z
VkRU66Yw3UK3eZafhHUdFkgG5o3+RdL4uXI2/xTRxYd+qq46BtpnNEZ0vecu
qBuJiyTU25KIYU0fFBdo9BO81bFI5mCeacc3dBGKIrHcAJz22u/GXxOTjSKD
JkpJiI+AYF9c/fwGmvAv08x7TdBF2+UZMR8fn3LA+NHiDPpDlUVfA2ihaVNB
uEwzxpnO1zLtqgaOswAmM8KGv9920ddf5gU/1kyX5q3dy7im1UGDRDoNqEag
J/pOssvFX7iCkFA36It5rLJpdb2LScPvztRtb4Hv8GhTBgurmxwfbz93Duc6
rtKVBQaClWlZUqmgycthzenmIojPU4+vWn1MJiOEaPJz6VNhDX9YdPF1Cl7A
X+e1HPI+97aU+DqyM0ZLv7/Iiwmvhgt9WSPcCuJV8JC35/I2Quz5FGPah38c
fvTD91drFy/ZIs2gS5X2hqdrwQX9dZt4lokoWByGNhp/qtySEcwyvNyBWQhR
1TExkWtyY6W4KEmTNWmQa2E06itrnIVXy8EfaRre7TdxvncNjf0r5ddCHUDr
/IQ3H7hhGSBNTExrV4yf+11BjcKTzglONh23kCnAv3Jg+CeV9W91qdWh/8T4
DygIlgQ9wk4SG2Y5W8pZxi68VPrzOQDV6dAvQPQQhn4oPrs2Dd3yZkXRlzU3
YbAFj7pBbaGYzOH/UBlRr3G/fU6OK12NS81ZYyL+iiz6NhJjfDEV77IixP8j
vC6inxyA9zhhocPs6H9MSrhwxP+6l1KT+OHUIzUvVNk2S2fO5y9bdobB9raZ
b9G/HcUU5j0CbB1U5ZtOkUH3xXPK9I/sTXcpoRhZWd3BCDw2jE/sKiehvVnh
Nh9sTYVX7IFxpOjatxwZ6iK+AWOfAhAPbXopytf8O43P1WSDyiyuK5q19Pox
XjZ1oMS0DAf1xSrID4gU1JYZYvG8XO+jAKte8HUDr53Koxd7IqQfdMFksWxw
Vp2lVvNiq0Cx4dkwo3RCMrdxAi4Ecy7gDZMJPFUC2wFtpLSx8NQRsTDxRD+v
BUQC8jo/dd+1zcCtzUIhcskOXet1zPYNIiN/+7g31xktzZEBzPu5M0ac8Na6
01sbtVXOC39n+hrj2x/BX/NDJAnsDi1RFDnKeWJ9yrR9tul+TVdUJl1y0LSX
dbfHU4303mil87B4qJJl8jvvQ5hMNfFLNGk4tXbNdlizot5/GfUXuVD9Y2M+
4myOcV9yyOSl7U1UJAMNzdLajjqqOxJn944HqpAtvb3qDFclFuNeMXqt6vc0
xerfJLlKNQaWgIUcpCD56vptmuM4ZfE0SXuZgawCWz9RSzRijXs80VgF+7bi
vQzG6bbsaMepcodP+zaYmB2stLkeMm1exg/mJPcfS8QRiYJu9vbtt2soVwm5
cf0lUWW5o24QTLs7c23MXjCo0j+DtZF5WqEq4sUWQq3LK1MkIo90poL9DQm6
5H5l6+AunyG/zpYIDrmK62SI+3gAs5u6fiUWqBuyfdoLaFtWcPLqanZXStCZ
T6pTkr2kSP3lgF79+zpAXeICy9KOWM8UF6RlU3rhTMGtNxMNgbRMvYrhclVv
vFK/LC2oqTdFNt7I3DzhLndCrUgQG0EwrA9aM+Cf9mP1Qn0iG3pVEkLiE4RQ
WYRakHPOLvyZYH2MzQFXhpYEBen/GsPGX0bAqIz2JP4FffqRVI/VGxzBYAyW
j7ksQPWFGjVtEamnKN9qwx+qzeBAI/qab2Uu4dWfYERMTEsQOcLjse4CYdqU
FaLcxly1ICMc+pyb+B6/67rZKahlvoC+iW6zVuutW7DkFNC9UNcef96Tt6y0
kLcU6ldLIjvKZ1HhUGS0MwU/RJAB9yCDkjfwI1oYPMf3Ban8UcbjBjUDzLCx
b07BtHXR5+5nySATMP2cY5P+E1o9iBmgtPhuzU1vD9JArOT4z/UM8gtu+7oJ
DfXLo2tOMsX21/LChWpmx5BO4WQiWCJ+BxiwQuppTZkNfUzwgxNhL7wU1CUU
EHkdkC+aawmVBoPhtu2+03XccEFEfTbHo+EMdRIsO/re0EDHINwn5/0rSBkt
aScjFWhTuo74+Us3nrTcSKDz81rXcRQeQm3+kcsMxhm8RzFuRPg59KSTilEw
AgfAZWkPbSk5/YtoSy0/mSq9oEAwWKtIC5/txtTL3ebQ256bR4taFwRbPEjQ
6QehZGvZ6GcmJ8unpia2GivbSBp0JALGjV/E5+MvsgaRdcVCyB+1dX677825
CnCa1RBkCyjQAUnrIkTP2YbzJBPyHUMutqpMmy9nAERQyZklUH8rcPEgJvwW
RLSgHJJ3It9yI+bvwJai4hy8ohUkkW+z+iMSvXp8epysreUUNJscub3IgbiE
+0yRjlgMIuK0lDtNaqcbwWAK7f3qfh1XMKGM4T755Rw0H/2BpCtxJX29XG0X
Lsbcr0XhtoT5da9DRXjj84gmKgAripUOO+gekM7Wvu9SKb7k5DlL5zMriWn9
tXqiwyB8DrCNur+bLAiabN+tU2s7EXEvvPMKPcKeWXcrPm/ixu/w8Di/Zng4
eDoYfn4fmv4YMPcDCVxKIilH5aXWV8Olm4lTfAbkIz0J3oxHjYWMb2oVfNP6
isfzCZOyMIhUZCqKENq7TF+GvowC9SJbgBuyd0KmOyGCMXIpIYT8Gfo9MiQo
jsk4HPm7WrjQb1p7n+/NvSz5yiK+T/Y0Olmy92hdvHOHicAH886hJCOfoogn
cj2l6L/jn9Gk+PstLtpdVgC0SO53Tq/ldz3juqnjsqV5gPEy9zUDEwKGjHT5
5YTzFItv2j0odR1pYaeYk3E2Az3grV3j+mnLbwD3czgUXPUke5483AIVHvas
1EVHy7xSmsMYxcBYduyy3D1epqqZ3tl73SyIjwa5uCFxVvgCP5frv2B2ANN1
Mf4GZxOBxP98OuA1/NZN3WXcSmpDfuMVwbAHohFefcoxBbNfLHScetevGRIE
vi18V3V9cG8UmQoFyHMx9PTf9cOWyUzbKk+LzD35Ct8b+lX1vQEYvtjMuKuJ
io/oNqkyWCslVFQewV/A5D+mqoki9g88dsBRDaV8fQsanjGrRuJqaXaqJKQk
/1qkHlTPgYbqnv5+XlPZBvLQQsnkf5M2WcS5RduQ/hq8bF+KtYO5d3PRUNPK
yWXUTJbZVXW0LKVWJKwRtVEcoUnSSkbAdqRUl5i/yjBpgrGg9UyStWkjsrPv
qrtXQ86QuWdypqQOzWAOhIhB35C1J2eYxgjWJOcQCgS0qWsW8GNp1PZgaHu+
67wytOQm8nCebGZefdwsC9MCpNx/ggmueL9j3NE2vgwmaBsn6wzz0SoD5ddm
7RR78kWaMHsa8vdbZ2L5KalF5XBkgiMd1NTfzrA8nnZWF8MU+4VKpzovoUOI
xlxXUA/xGEGFVorBBKD9ci/B+NRsOaaLENnHtWKHYp+ba99fp+oNJd8irBnd
qbdwSn4Ddvb4Yi9uVxMQJLZX5tMqctvv6GddZvjTUT3L/3IK6K5UWEI23/L1
Rgpkq3gdO+i4iWABUlTi4FYViHn+Rl+8MesruiWkPln4s+zV9Ygr24TLgWu3
fWCWWxCTtap+8PD2OywWYcUmYDdiDkPgPqVohuWnvsIzt2xdb2sB6Z2AZb1S
GY8Bdf/bNMH2JrSQYHblB/WBnp+IC9Dpsr9Vj90SdipAL4ox5eLQN/bdGy9X
Im7MxA6naiGPn0ynGnJgpTHw+XHYBAeZTIB7VLUx4W4SfIzf0CKq5y5JRHPO
uwHpsLTS3Tuv6BQiZCi8YrV6Xjqv4bhmPzW73GO49y3hCJDnXivk9cpSpO1u
pID0m6tQMVSp/RA7iwuShzl67rvUw1jY6SwCyfPFA7V0eZZyiM6/T/Y0gaEi
GcQYZtMW4HMPa2KXMx6zMSeu9YgSH8ItotRx25EEOQWx8/SjOxep2N5cGMD5
Erp3tkWpLMwJpFpr3PtMkuNv3mcAPOMsF2O+gSn2+86U+N5qIYA6HiTc2Tq+
TJjCAlQVk99a6GE8zcrW1IZUpCi8G2cvJIdyX0gadgMjra8jfki30nSmmhku
V7bNolO1TXc/NB0PSuy4pHCrNkxU95TNF27dS7js9TrhcGBxktsyFBXxVIEb
j5B6sdsQ1HDwr/DZAGES04oyY+uoZ/87kbT24IFGJZx9Udea23ecc6JTbVD+
ABFXv5RZ/lMkLSwUCroH9tUBRPzYkjdT1z8+l9ejO/78Owr2FjApatW7XE9a
8yckvKrrRinwFqaT/4JZqG8/xpNhUukeMEXjaZpQydY8C5YUVZpQzK9x9yTR
omowU4JVLqCcdQ5JrckQuJfnoJRbZEKyF+CcpD/Fca0VaXaGQxMXXEieZ+Mg
U9qIfLydq5mG4WElQd8s60g9b49yFmFV3WuaLxza9fy1jsdhTjPF/tC5HltG
KmANCTIzJXcUy9I8HTN4iS0+reho2XUnzRyBDCzIM8QIVog3oayAg/YzXdVc
GLBo4F+jm8Ij/6qYbwyTlQIEUU1vL6xv0GwOc8Q9RhSyU25b8jHD1ydrnNOk
Z3XoOQWGEFz9wpAqAYt70/FHULl/xh5XARzJOdkZdwp30uzubrj+OSfderqB
DiVweQJEWWsU4SkcljbvHL57fkrwR1jhcbO6ut89LX2pL4xOwPlWvj0wJcNS
OQIBjltf42UXKiBw1l/3JfxC0EHyVeP7MvGXHGfRO9eu1O6bPN9G2yRO91tc
FYut5j9xivp/KJO62Od4nxCdJOhcq2v5d31rZWiHM91IZuuPiXyW6hw5y1m1
hL3MxK4f0Ld/CMv8pQWXNqJkOkLTMxRKmWzaQ0wb86eAA5g8e0W1mzAqXs1x
4TWuB3w/dvm8ruLmNhvTthmqx2+rfcPLn3su5EVDW/Lfq7HycqJt/iqpvn0T
QcgB7WgTxZ2CFxHrbM4tpklcg0G16WEPCZvSkou6GZGx7M0WyHHx78Ka/wge
FCktMPWiSuhfP/MRMJV1nFgKoWTiBy0YG/w5frPGAA3vA0kYTZLoIjEk8gJy
jdO03yy2EBwJ06C7NsmtSaI5AaLbq3ii3mwjlvwLmlyayjANm1QnwIFpfcsC
edATNAzj3XrGh7T/WDkrs5w2l0nI+Xh+sv+OqjMsftZoHJkHKzuQbuSlSDUW
OSakqK9D1AErYpiq7zPugahfC4UBEDxKNnnwBoaaP5sxIznwRmBQt7EMPgUQ
bu84+SKZBI+IDneNF6Y4bE78R5UwDnOrand6u7BE/Uc3cVRmt2iaaUuDCBSE
umqQ/CbndA8ORbi77oug9z1EbG2Rr7QfOghzBvbZOIgb50WvZ5p+qN36U1fb
ThAarCbyWKBrSbctJ7kGUSDmfX4lJZIq+PW7ULyiAVgUq/IEidxBZBFueo7G
u7Eg/Qgu7EkzT3TF+qKhPBR1BQsV1c5DZVQmQ/ri2azQsh78blEkHCgJ1WM2
WZN8Lt0k8wDwO2zOAniQVwGFZtf6J2U0NUGuTxTVknogG9I1HG5fUpJoS5Iy
pTaW+VgQ47sPUpSZrfrQa3DMLB7lHv+Z28KtjFtlMSUVzveKrIk16Y5nqEp/
QZqMnrdrpXlcFn8pN5zgkSNbJ5vWUJsKFN1rPj3YmnwZHYKHOT2+dTqbNpTe
MSCfWXsJcHD9lmhXOfWsQALAwa/AIX2TCSxmWTywMS2CejP4VnKXYwxgk7uM
aeO129Cr4540ns4kS7A2Nur51zdBxw7jav76C4EQwSoz2eL2yCGqtKwcyaN6
85QBdhzHKesRG2ddoVxSae8dnFOfySnrYdYqtwJG/qULyazC9mrQuqjYqra1
McouPz/7obLl7JLr8/sgQk29FeVQUpJ6WsI/FSXYsVU4Jlcsh3SauWKp0gW5
ZFk+mYqB0vLxCw4kewy5q/a88slAmsJ0LfnC87NAyslxcs4xdGvIZRmusb5x
I19cbAm6veAQq1KwGdm8g8xfPaQtOLbe1EY7kK9qPn+c7AYbh7xCVlhW1pdC
eWclqOiY5dz0+QQ4btoJiLdeyzufmnuOwaPepa8e+P1GFV9OTOR6BRHOLjn1
6epE234/05KAXYoQtGU1lsIF4MoCd2jJMM3xfBixPssWjVZ5yFIvMBqhOU60
qubdvtDAWJ+kUmIkInzPcLefziSqEO8E+MBXC+UhkkXoKw3x41ZFVBaULo/F
op3GNyK46Xyfn2lgk4KNDaIyZha4wtDmlMKKsUpMGxJ845rnhQnyinsGuo+o
X7+9mWomqJe70wkxPP4QlGfOTjuciOcvV8vSrKa3xbYasL0cKtCaQZKsk7yk
Mhvu0bmWKsrQHrf5XvwMVISv1jKF0l30Grl6JWn1VDfVnqCWi1ICBRM8V6aW
UVty8F4YUzyMLXGkG9XRD8w5BbCSeFcCogAXuV69hh6UU1Vps+Dk0v1WHbNP
gmDRbecGJlBFcegLDUcZJ+fp0fJpXjERNydKKYd2zSSS0XBM+sPpVMtaUv9J
xg4q8iS/6zJSG7AfziCVGzixGrIj0v1YGDv6a8zFfzoqILs5Kn4savNhr8XA
bZvMs6wUVJrIRsoeK6buwwXs3sd5J8hImIl/scBuct97HRBunYUZkqxAGqaX
9897dOEt+a63sKhB3fp+L7c2iouQEqkjRWfm4ejJaLvmek7ambvVC7hhzJwr
O6Gih/p2fQJS+WFge63reo8ZiuTiJCVTgjvtovvFmgoQyY5WCSd5hehUUWAT
685fRD+FB+CDu6/i+5p3ZxEXnjaWTJNc6JazeZp/8d4x04ApxT948rSbpsC2
KEPkhfXXnq2Idpjpd2TpSKVSXjB7DoWsdinu+R8w1ktKR/9EJAHDv3CEq7w6
757ScgrviNtgs0CDlvAG49KCNn63aAMh7IQ76bgnu1HRlpMogs81h5d1u38k
Z+VivHewOtP8LKo4tq201bh5nkFBPKB2Xoqnm2jxZEh9IHPC5DfN+XzjTrju
KlLb1MNNSlzJZBFM3KQBGqz+t5Nv9Rfu3vMAsqvGZTvnmrjwUd7jfKM45b0T
hocop4IcuVa8Fn4HBRGHDp8YqvZHi6EyiDMhmXsYo5pmSTbh+hgsOr3vbPEl
+pCoH8Heq5Y21zjhsJqke+VSVM5VCWzmnP+upBWBM7AYNU2+Kj+UUgqdVwv3
zvhQmCKAp1Mq8fg4nGYSHpPiquomkso59aNvJMpvxfz1dL0V6PT7N2r4nB4Z
XniAulQbm8ar8nC6uPOkeFs8ZrgC3uZt8ilaaaMBXYkpUdn9WnERCx5Yuvox
nD3XWZFORVi179JUh+1J7yWIdd0ZgSbtEmUgGWbQpqBsYHi+pTnkHsVz/2i8
YjYzl4cJ637MkqlO8ozRYJUer3g/hTEMpGf5vkrOMAlh/p86TXKBjI6lnO27
9MknocSb1b93G7yK/rYl7SkjXJocey5nOLMXGhECYWVgrwgS62ydwj8oarat
w9xKqfe1XEIAEnj6SGhlm76I2UeN/xKT02wN8UMBLexO2672W2bRNpaqS8zp
G5a7HiciDcHqKPRowlbXW/a8XvlM5bFMntx1vnDxWQ51RyDiXxHOl/f92b1t
SlCiuUsLoI/KQcaBSu5zxvhAIPqJcTU8jkEyEKqne5nXj4yt8q0CFHyWMPaI
EZmp177N1w2lv7LBsOVyG6DlMZm+76M/rrPBJJn+QdAES4h3cvV76cdLb/5w
n2LWll7phMRqQBwuHFFBtllraFClGTMg48JLatyGFrl1WdgDY9sZLyjIYatE
a6kUjpG9IE0IGBsnEGiHouCjYljzE+tVwTqWrRU8A2zaKbgd35BhlKZKkbP3
DPrRnEJMJFZcvfb32fKglEpKqVK9i0pS60qwcUSD8Xz3w7L+/xccykGl7a79
El7obay1qzKDCMgETmiC4/ygPn9pIDy4XGIrxKYY16CYas/5l4rxIGCP7uh3
qYDzV/h3xgwb/2y/KJIowln3oQEq+u5HpI2DZxuMocvg5ckUnGniY5363KfA
K3UyNmevvN9Yk7JBafFF4Yutr0rrAgT5/nqqA/Jtex6jBEnjMjbcz4jz7GEk
KAGhsdbIB428egXv+/k8JayU6Kg4ryTZGN5c/sbLbltV7kdOkQvv0DX7ZXCi
NbDuoA8MukIkErvVqP3bPTFcTA6+7aIkf3V52ePeO+T5D/mKl0dHAnNDwcP8
CAOtf35nkvYf/ucZRjwfKpW13kxRz9idEIyli6442Ir4vQQUnY0UcVBqyvX6
7Pr16p171KJ6d5FFuN+8yUPiAdtPq7SBCcM870oN8TjHJAIKDSEZjdvBtI/t
n+OHXlCrSvuD17UxFWxNw5MiV+4+2vGECNMgfOCYkl3YJyVzC9WhzPAd0l9A
vnajAeR75Pf1R1h2kSaI1ZDhmp0le+2cfsSe84lAwo6+dUcgw9XEBpT5jRHR
gnZGtq2fyjXZ0ir8mz0GH/KDVF05ZRfiSCcFw/7zB7XRZ0On6gAtuuitJM2z
sWRuJ8P2KWohm8YbROzBnkFjkMcDUPc1/pBBbMDY2ZoKfDHxFYPgu86sEara
766t516xgh4xKq7/GVsNSUzO6ixDeEQcYqG3b7g3xTD2ZSxm9GbFM38odEYY
sTkpt8itJS/g3tlV4PyKvDPOso4hRFytq+84wGcDOAUeBTPtIt6iXx9Kt1Jw
YkU7Qm86GZbjXLzODpcnWJmowqH6gxDuE6XAhA9ZWfzpyT99/nov2NQhYsvP
lV3RpHcsyFNhsyswCfSp9tMA700zUudHvMTzwaFO2xfKE0eOqe2Lg/w79+3k
hhMJE/ZS0b6QNmXMFcOEAoRGRC8nZY/4VKwaYorHPTbITQc6GE2caaeWg/Wx
ykLTWVi8u208ZVx0pNQRQRpzEKlNgc6hvVuxqRBk7kurLiroRBW/oI4qifxt
gh1rcjwxCsv7u5wfeJadVrKWkatoL00+W+RnjpgArW9em+avJSL/x7BMb0ta
UxDkH84BrjappzLhs88OLDZ1MgIVv3DNj8x5fLR+OqIA0fJ73JHw7Z96NiDq
OwxhfpfidIJjhq0oUlBVyV9pEjiX1K5zWOztzJnf6AeMe3YGf3FWzxs+W1ul
e/NzFu2kjrSnMsWwAc8F7tBLg/aStd1OzLwScCBSsprN4lQJcfz3JhVmuJVm
64JPpLL0+cFBkc6XjIluAaNoLmLSRwh9f/9fso4iwu/qThn1B7pxOYhsSnzb
jA6cbE+c5RQUK555Q50pFncnh4VT5mlB6mDx2W/h4k9M9LowzU9z9vI1dPIM
V0Deb8jiQeX8HNaK7vzxA4jyQ6Grs3wiYcPURJJitSJ8gG1jSzCHFTGjNEFB
PEFbK/ahn1eydBflAYEih4iTdMBZloBZd68g12KeXThMQaQKrwcZG+8If2kr
g01ff9kDCZN4OOBsb2xzlJvXB2ulLIRc0LsnHdBpbsd2ic6a1SFu5dlDSvt8
xe1/90wJZVh4X85ZiAKYDciOI/h/MGNIfAqBT7Aj1UePctWDuinjYV+W8AcP
Ri4BJxWO5BMra57T9yDiuKpxgpzDIo+9T+47QUMsOYVHNqhTvk4PQ58Exwia
kySFstayQbJCGMnkt36wzf4gq+b7N+z5l8d9pznY6+nkvHOIY7iCHpd4wjG5
uDoqZp//VhNEF6GF002TuoeC5KLY9vjaFa03+QwlUtiFaY2R57Avsv63fvMr
Fy5HV+DcZre2EqAIFxC3K94E9MWjbcll7aow72b7iuX/3JleCR0ypz6Q9LxM
/76ujIcPtIPEOcTUsbr16RZBGG2j4+L+y+fL0nEw5MbJkqyAsj/OsxgBDKAF
klU20eKF4/qBCS1ePSCuuV76sqAW2qODcn8M4tfrPMJQEPhM17AkE9oTJAwj
C3kFNHqVtoQgL0hOcK+0q+iRnvS2k+I5WRqftSlayyFGH/Fto9nEMGMzM0PC
8Of2eTuYltPaDo/x+IYWv+nVa/HNcr9RbvWc36cbd8ix4U1kHPlDzw0BU9t2
uCZWW1Z2OUvVaSOZVQRuDyCuFEiJlXqZXO88/2QbEsw3B+1M7lUO3D3jD0L1
AiI6dcZrTWJBjcf5QpbPksryWO+EvlwbtuzNatqFLeVTcTEj56oUcGuASZpl
6qyOzvNCf0EsYqRamzbm18vvHHan2nDHoHH7sAe0ZenFKlLd1DVrw7Z9biBu
DOzu/H8gMbN43/ZiL5W7riRSIo8iWtjOVjQjOa5ZCpSkj8TLVhSppDIYFdmF
cVMtkr4OpE5AjQjtiglegRQwz9SO3TPvxiCzvvQj2veHmmR65c32cQlh3AR2
Cq4FahwcOmr+2k6EV4Xxq+Fz7a2uRUoJjxIStMQeIgOaHvnYMW8aqbiuo/ve
LcpDWurhCAYXyRgiJ2isZii31kbOcVIQlQUFQ7kQGmUbk2VUSnrIxwqeFCPO
I6HiLT94ujdWPHusmvEiX1h3wpiTochnsAGRg4nheBckOEdWyQUCm/lhWgE4
MVTmzsO94DdqkvMfoqMSQG1Xz2ckcB/kzTlBD9T2HX6Atz2Saw2jNq24D1do
Y0B8cE9AIxMlULA/BDfkpg0WjBgPgUP+Ep56ZIVyY7MyvN2yDiAC4rtfyGds
gT8Al00SnLCnuIbX2TcirdmUTg3GydHgeOWNLAB5/Rm0c33ezBrddWUCeZmp
8z5L5Kw8s6f/KSWv+ISFSe16oOtAYS+050ELLk8kKxK1YAvAQEK0ckTbc/0h
X8B8j+PQhDExvijK4cinJPlOquBfIDbO+bUccSOccuX4COM5KDiR0Oxi3xFm
X1j7dRkaZ7RgtcsgFXLBrkerluyiRd7y0z1XO6AEgpTHooL9BA9PcM1m0Cno
sE5GmPiasn/BIbgRGIzifwekJUwAJa77p2wQPX/fJx2tlcv9Zt5Y2lVVBkwm
vS4i4bpXkTt4GzgjkF4/iwbRtYETO1R6hz12yODdeneKFN5ouX64XlhB+Ice
LBwX62FzpYuQ8/7KELgTURsIDVlU/XNLlOU0xGxx1w1X3jEwhZAmA2PBirWn
WUeqxfaMP5GGlWGcUHkxdSVitqlUibdHd02kBNcCOdJJaKki94JbQ6aLD1m9
nkTsWQFpwytpVrFXNy+edq0bn6aPBH25ZAmzPIQlZAYijLge1iAscl8Zthlb
5neZ0LFbGjhZrJaTvynF+VRsGc53YgVqP+PKHtamRSQqBXPqAasOs9gbVQFc
FdvxwGY12H5aD2g8v7QwU35DyMniiM1iDRjgkoCz52XHWnQPTm8Y4eulAkRF
Un2eGemb3YAFxsSMDWs7YmKs/rNHmjUPZ+prV1txgS+PHn84hy7sPO3CWcnt
IL2B7s4Hvk9BDPfSj9fOdA/mQARRfj+2e3DE+xY51FuXnnCYkl/oFx1gqNs/
w5AJm2x2ruFjnuVhmN1nLn1kjV2dLWi5DLJ+nzqO6rmzjmbd9bjm2sfRLmf1
LBc+lGhK5CPGG9lNGFG6QKUNlzE4ZMHcahBaFVFWMquKJ2ogWg/+03ls3hz9
LkoHxmornr7WdhLH3bU5aNdaL9d99gVlur55UNcS2KR/OP/b4RtlHgH29RkR
uGH3JM1rIv91KNdE1s/5sdS2yR7/ZiSrFhJKZnbD2FlpT0X0WrPAPg9sgaOr
Zlqzqv4pq4TkhcMmqatnMHTtSElWTSJaEONOoIKAFlcapPmuMruQnImr3LJV
B3LXLZloGc6cdQ0XGdwcLHme2rqn8saOHeziDY9nkzpou+uLlTvOJEpeg0Xv
fMDRUWIXkxgCsFmeyVYnIwxg90fM8++BMwdAXnRqsIAuQB+vRroL2vxnUV3i
q7k6Mu0hzhxy+OtnLRWhWnY7S+VIDYMrzn6LLUfdqsw3RQQ/h1sj5i26Ool4
mYgGceJWPE4ryxCVM4pBDjBzQMjtsq4Fr0KRWRf45gtDBLX7WPOc+6XGPxya
bLr+aASzYUkl3X6B5ETqqS7qxDGa77hfzRnqmdQ51dXYhp4JMZnXb7GKDDvc
HLV7yOuyZSuUB5SrOSJH1sfD8xZ/JpVN4GATRPNvjv5eE4tHYCQxXexg5a5i
vs41+nbd8boGLyRwaERigCI5xHBdqdi2YqCwsif/FhqJSxNb5J16FOB2JWnp
A0NuS/gnQhuJeiDErs2xQfB8qcCXgcjQE6IRlRxFIRHCLiygJFJNNtv6sKnt
8yuAa6N/R0+AeofukkejHIdGxxTK0jGAHy3I+gdVCFfc412C59KhmkFK0L20
ExoY8kvCBX6ZtfGrke9WF68Swt2mq/flR0jrp4OrtueIRYwkgdYdc/6RzARI
F31kQgM+qb99Eu/pvBS9Pb6vVE0iNIdrdLI52vA+Hq8B7hM/mo3dpY0hHPR4
g91K8rM6Sv2Ri7mrzvf08syTo97+Y2wCJBygog39nug9MYH6LHEuxnyFq14K
jvzQeOcjVdxisu8JDYPn2vNchUopJHkecxdLpG1dN46poNhsWY1nukqrfwSI
IPqhaCB7LPPV7AkMIGkjv9MiWZ2oaZcRphxmnOgV7Sxn0hmKOSUScrlKldcn
eU+17mNt51JJX9tf3CokndD9r7ff6+ZwcbSoPHfcrDAyJPfcGdFX/5LNhiup
Zwg3jBnltISmfYjj455yx5BK1L9YkHYJCpTyPTVMwCNGmWIBoRcM1MQ8Rwcu
R5ZgBYenWCRGMxWPnkDrDhZ3vsgOdS3cSh4oZwIIIRd0Z+dhncIkNDuD2BDS
5cwjFc4iyL1ExjATIjgum5LgUfD2H/evaAY4ZFdK+E9+OhSs5wp9BD6u96Q0
zV60OFN4DisFlli8fmxG/vqfRrp+d3yKlZWmVRS0b2FY3dBkCqybm6cJrjhh
sV2ehKWuHPXNFPj0lzd6GLpBSFuliB2GjzR+JxW8826rHnB+grcqSdOjVblD
2wcx+CH0vPjm/QDgRIU2/uujPj929LhIyCgj6p2I+y/uz5moUN4LB7Ntb5Lz
nBr9pjqSs8A2aFfXo9LnnhcxPjU1HpMrjrLX0157ni9RTA4pd2UthuPWhucb
zOVqMoG8U3IDGmtC5btkD7RGrZw2gSu6twArK0kqkmRgyp78uHvFDcHnJw3w
Sac+vzpag9mb/fmFD0ms/Avflz4ZMKEwAA0NVn+s6sIwIRwvbV2I3frk+O2r
C8SyXtWb3301MLF6p/E98e+O5633a1k+qFejQbRG5150xbir/FJsQS97pzGX
hIUkPSmPIW1pde9+XtFa/ghs4QDcSxyRsjbp2vYoSC35XbLJqzFj+pN+XeoI
eKwc/9t6CrBlFbyIj75if0tIhNjmQr8e4OoYpHcwshYFuuhAJ0dw8F+/0Joz
Fk84DCbLriblKrtLqKgVKIxlDtetlciKUHVTCl10SkgYyFWsJ8Rb5d5o8nZz
Dscby/RC3YSFf73fyVUdxkuTeuDqaML5vDmy/DAo5TO2PfHzQwXoNJE9EOZ0
c6ReuPbGTb0oiMC+408VsSHdy1AFJMUA2paHT5qv4rS5M1SxUd6GNo3WaSgv
ENadA2e3gi3ahdqraGSvFosVkxtuCCYdVZ+4L+YJSRYtlk6yOBaAiw719YWH
INF4YYbNX9TS41WW2n3OQIEOoH/kCBmYv+haG/Hsb+WClNdrw9Q+GoVgfawC
KVeGgIlooGHVtfUrczb+7eYOuAavIwlOT7ddthNHFv958IMg0gXhmm/VZh4L
D56boTvrdBA9MikPyhRI9/gyrz6IanGk0W6TyC3SJmLDfM8sUPYLRB1TEWe+
ZDzBTw/j5ncYJHDQNqRZjvXhZuM+haS7E1HM9HChR2SfP0djEEV2HWwg64Uj
aaBS7wwtgidYfHKw7uuqlw9tC5DGf+LCJd8KIxjLtIDnqWiGOBxo1fM3z3Rl
szeCNSj2HaleKWe74bGLv2JJTQprlnd5wDC9qQkw/tYzGzobFzdYl4EgvLSQ
v6dr4CCXJPb9KCUpajL9SrvEKO+ytkaB2JCjlia5vaHP0M66wCIC33dxv4pf
zqsFQwIEj4rsLcdQCgZhXGJfqvrKVtPeIXvhArHdE3NSljZZa6JRTylNBDV4
NVTdDW1uOA+0sr570i6afAtKXEAeRAZYOTmjGizEOIFNux9icA30qy1wIVSK
x3VUvymlYWNgpFFnRqXSuelNe6NaRhoA92cmB9qwWQ+DpAkzyb2mDKH5B2K+
UmcWjCApQhYHEN39E/OUtw5jF/BtgdIS9/kRCQewPJ7CVLhtMzpt9Db+QGWP
0gPths6GgKk8KD8wCWkeJieoJhopkGiGVrd14iW5C7mgNMYiVm4XGdFb2MTf
6XwT+hsvroRdHB4wmtIgLMiuTRufw7emKh0K4Wozv2Hu17dW07sMX71TyTVc
CfT3EDo5mvf4+aErw8KgN3ujVsSvTxCTRvpkGz3GbTXg3Y6jn019esQOJqkY
xu6xt03eGUk23WnDIGJAwjpkl5CJsYSUJ7v01u31xr0XIJKmUsnRf7n4hj/4
pvPU89wszDpsPRs2D2cH4rGIyy0yMqa/eat+fLGU/CVt0e4c0O3gZfcmCMpT
emLKbCVETgxB/2IeYTowmyqoJkAh/jdzx9gaRnz5+Y753nOiWlUp9368rB8o
zGGEWk+N3UfL7deeOrfAfaLVhWLDYAa25xiIpM3sRy/pA+xmQMGmgijJ01FG
2iI1SEf/tTOie84JpQdWJKyyE2jRn9Xccf8yLsenLrQnHV/qgEC9LhXm++Qh
dNtVUueM/wBBW7y7Lzbthdb5Se8BTgHI0dYj+qThFB+N+P695Bh6SrhUZ6F1
TtscHiFfbFTuLRGAEcrEnHtae++P3vIwkyciPDFOoOjgjp4L1u216/eMWqyj
p43PrizT0nlzQtjXZDvU+Lixcae8VTdGvG9FPKYTeY2TNuu3pm92Wk58ZhYA
m97oCViSD3XHpG7ZmmOYx7UawC4ag1kzxhIZN7r1+WPIW7GpFND66kRIwSgh
kIFiMxQHKT2uwrVwH3G7d7dXLF/iAXPO8tb3qdpnVzOoaDTDFliqsovtfmws
Yb3Ya2w2bGDceooE9J+Cqki8Bxn5JYEGhQZq07CBPhFvbA0ZPi6DV07YaGsX
kvn0AAZwcFK9E5sc7KNrvB/V1i17h0ka1GTWTGWx//x5fTvlSot0l8cNpc6s
AOebX/U7oP6q30PpAv5DQ/HVbHBlH64nFe7CRGxJoblCET/X8pIgOgEKnZ/h
UVl5eX8Ms+YZaJhhZudHUCdFIyjMNO0Ot/UJ4/T6jsgfPyJhb2xjShy+j3gy
fETZj+WuELAdqAEmqgIOw5szRzVGS9tW0+NQlMKCSj5Depv44UVR25AJBo9G
eRtWzyrvVRaSIsceQKfXU4UWhjDCCpZt7GpbXCC/59991bMxWoReGQHPrxSA
IA4NtCwSYi/d2ek4H1x+Pa+v7BAlKQKs4rPCbflptPXZ2NxuqUiOQ57PTol1
8pHRdhjTXZrIbtjhygGdiML6DnaX85689FWOyHpgNzN5tXxJo6Jin7LEjRJc
9CXMtKsPH1YTOQtvGKhBnysPx7ps+yHYHBvz1mb08+IQvQZ6txoOnJ9mJrad
9GE+hBhZBJchuFWfyWYfbLPbq0fovfMIIivIF8IHLNRXh30HVzXco+JC8bVs
RR42Qa/31e1u9MCyVrX/HFOJhuOUH08UxB7u52vBDcnLnq1ZgmADx6VgTVvV
lZFKKIX30NiQfk5hiCeZrCW3+Kohg7OnhVtJ5h+Rs5+jyQQDNEekcN3gkLZk
YPvcqj94kl9dlBsca+As3waZ8XOebcQM7X2DKPjPqFGNUM2J6aY/obH22ssE
whJwotFKBNSZ6c33BGCVeLt+lL5IP93xw5Ph1P7QpE+sKpOJQeILHqfkrOsK
6231XBGPqvsCyfOcQ1fYHhWCjDi/W8Sb+aqL+j2dU0Fojq6CP76w2XJ0SaFO
XtMjlEz/Nt6d3h38FJUo31kKDRjvtYAN7IulajfUnMZbKt8iguufr2M1XufY
UNFq9RCg91enH/2vnn94otSbQNzPRgfH77lmlblPwE86d2BxeQSURfW4oREc
rdjDu1TSElRyTUS7CArVK1t4XaBHdF7ILz+1pI7kdpp37iVxZLzENKlIrEem
CfSJI2vHVXQyYUW9tt+REqbVpVCQgV3R40i2oOJeLyIpm8AEKC1LZubZy6kJ
mCHiQAiyZBJcCoDR7ADw823GN0swLqMwbuNjTM/V75T9v79VGcRjIYLqpL0V
8zkGfobyl1wGRECQ/qfh7ACO0rJNTCUPTXB1W9SewXzVFw80iMxllnuhxvKB
oAo6K5yfsIhsJjH6/yE8EQsmtIx/X9gfXhNX6Pdd3ZCNc5Zw/ZPvUDqtQtS6
qD4jEI2hhiZQ/KQCLSvsl2EL0pbRfA5IT3fEmbBmDsUFLD1aqmzeFWG6EMS0
mTaUvUY+WyAQJoTEEw2Dxlh4RCc0rKEUTENUw1OlQs5agDOFxgG0vyCZ8ihY
NfL8h3z5jseTFCnXar/9BrfJaC3HpZLdBDZZc1IQrs4/JSPicy2Li6A7UBG2
V4+HVEirM+KDqJDtM5r/vEvBxHU7/fuEIMktCvKtJH42qC9OfALs7cG+OFLj
zXfELLm83FVj/K+fGE7cO85od4qMuVqX6/orHnaRVnWSDPFOeqaoYyH9CWdN
6EfbViAKtq1fzSEcYipx0spx5aq2IFB3+q3+SGTuhS8xoz8wzBFNqQIe0Gnp
FECOtzx4GKYEIBzWfsF0NqXjelM/nJiXUIC+aJFYlZIeIgaGk6JvcH/dmsRG
h7JfL49Z/CqvrzA9FhUg9fE7ctqakz2SmncVdn7+D/PJUqHUD8wyUpCHCzsJ
pmJASEtibXgVJ3/XhIDfyJqsY02r0aAvnH9VpAvVR5JRvHJ92linPateewY4
KrhHBfifxFZZ8UZ0T0/zzIe7qxhpNeSV7HFyHdjo0QGf99baw6zCw3InC6c2
iWVG2qSD3y/w7KUjQn2jdRMv5kPd9pgtAd1bEFBj9YrFb/bsOWw7G1OMllA0
hZsXJ9r8b0DwlOpaYvmz3UPGJjW3O9zlPhnT+sCkNxKciIvLCsW45pfcJYbv
oJ0Msu9WEU9VMJaXWxx3r5/Pzr/kXiGIY0zk0mm0PU4Y4A7oFd1lQFtNSsb7
cJx5JQ7CxAIMslgAXVyBtW6iEZBDSNaZoaHst08A5w/4W6haBoJWghYK84ZX
vQd/gVkJvT23WDooYJVE2aS7TUxcj0DmURl7M+5NwZ9FP0tfYLSlw8P67a38
dQj4G/aS1EuUtdSvORKXNS5HB5NcDyoN2N+LR+jtM+puaY0FF0CO4+/BFSmb
fulv9cN2OjoAexrmOtyXO711LQd91XTMBRYWmJwmeQfb7UkNrWhSRTQ4xA9C
AmV8n5ZihtS/c9qiZEl38cT2tV1tOmX/UsX0TjLEN6IicPBGwnpLerS+eydv
1ux3qEuPwr53w1eCpDP9DiDr/Apm40UUbLKyHkdpUETAdjiOqo4026XxXKag
MDiGc8RRufyijY4QO4AJy0GRagbQ/fURnsjx9z77IFk5fT5C3BOKsRWSLvNH
ury0WYhEq3aufznFg1Ba/GaLmSKleRj54umla4WdOiK5xcBY7UezZLiOHAnR
fHMiR7a60ToN8vp5EHgBDU0fDmR6qJ1mCVnVxXIn+hF0W6dqoR1j4U2Ulqzh
UvqTH7GSd3gjTBK0dC3LdPJkKJtps3zDyPaiQTWdP8Pze81jXtBYtPzf7Nsl
Jhb5xTjIf7kC6aUlBePC/5C4wFpWPB8vK2g2Nypwu7Z7+8qreAzJVisUz51n
UCdVi0AcXV3PyA8n25YO732Di2rlZEGamXiLtIEBwVv3mmb4nYXJwMokrhEP
lMzapuwxx/NWANZFbgYoHQnKJc10T4YM9Mx2dBwTO3pK3tZ51gTX4QuXuG4o
kVm14UIf0x2OKzfulUo0YJjKgMls2Ke0qIp1I6qj12IItI3r93me4K9rd3BQ
AwHyeQtmb8uwhv2435A6nu8HEUt3OuSBqY6/Njk2aARJ1VFDfCUATYpxdcJ+
gQLbtEWkVVc0qthWEW5kYtRDspcPB+MH+Fh75KRxv9KLy48aKXPYoo/K5aCS
YukDQik/UDDy8QGLECet5hEgZqec9IyiyYyzBm3TJRgP1/J3ZAl/dgpxNRVJ
MI+2RaORYpk28pdhZEez4dIteDdHdElGAf2lgGjZnKZ15tSMCl7VUq9GYDpu
tZ4zfDLuQTCSV4bxDZc8A7dXPZLtfgRHF/9Aey7MrvhOcHRjbDC+KOg1x7lB
u+dI/GH6uUIG8NWd1xzFXi52kgStaJY9DkAGbhRewIG2jsKwL1ZWUc5uprJ2
L3Cuw30DNgTWxdZ9IoZ0q6jjYPT4bHvJqQjVrkIC7yV6SzJGL0Z2m9DqQ76N
Ya0HY9+80CdaFkUMjrVo96vD8hdtGylmg3q2v3oAIUx7hvhmCCyaB7C6vYC9
dloThZ5Y5TyDgB4QFWzIGksENb+I7y8lwgaCrXe6uSiixiSI9NcPpRc/yXwK
1+M2gkfUVsVk3/kdLLh3HXr2jFN9zOf7HqbO3gbgpUtrvsePgh+b6n7liDzp
tMx4fEngjzWIpQIfhCRYVFMXY8mZaIJYkKQ0oQ1Y9/DrvauBljq+2COA88o2
R6GskQrR6lASDc3VDL7J6paf4LL/qVYheNHTz4VW1F3p8mjZjrLcmOiQ5RAj
mHx0F8k5teIK4uTQLYus0f54TXY5HzSn4MxjtOx1XUD9h6mXF1gvb9GYC7CQ
IQY8STPBhnfbEC4VWrLGHiDWnls/qKNOibx0i6LtXUZk7r3/oYkINOeEKX9o
/xHQA6a9CQ8taf1xy3UYQwHeWBIuUyPoCQ8h3/oKwOU1txKV0Ty3nnKiv4OL
i2R06lITWlHTIEsYdMybWhKyQDbMwekmKzHckcpKiTIvt14eH4KTOeOPmQ6N
3/60H51SYuIdMHVUm9lzuPZEA01ck2jObO3/TRqM88A0MH28gH/4oQTBXnMF
86+p1pxm6qr2AlbrowqNhYboSH0UiIurkSMATvL9Ciyv9v28vUHNgwXqT52A
WLZhKVtvnhlZs75a9ge6SVQ0IOrH8ynLLG5s3YyFnZVBxTjQ7kNOsTmFNhBp
97l596K60kI7BOxx0nu0Vre2hFGBgq9Q7snoWdf+ehG74KEipnNNGBTHsZwo
H1HCkvIzJcoHF4By9NyXZnG99AUUdgE0+RXk2Xvl8BTVUKiHdZGT5D34OjnT
0g0eTprgRpBvlOmww6/waw0Lq1twQUoesc8XWGxAgOEzCXM+FlXsIc0PZHuL
/3N74Dyj2exxiU/9Wc7T42RZ7GIo9MAQKqqvT6hZSJZpw7GJCdMTgXcmp+Ie
kw/bZmpiP/82Gh5e1FJo4KxChkdxhTHTAjGkyo7FE17mIv7TABYOx2Rf9w68
dISLH+enfSz217NPvwOeFrdlOqrdoqyJBSUS1S/x6GxdK2kSdsMzwJhqW1DN
apq82xk5iKruc93+ljpRa5bpJRRBkdEVl0dBmxuGCIDG5178SAvhQk0egi5v
Mrpu10vbB5thPzvUE31jNYFyIJFz/ZaMJkNt4ycHF9yBiLuiPy71+Yep47PJ
gIRZd/BdRkWMM3mtSIKiCaldCu9BVU6Z0eGxfiGAekHIkUpJksZIsrJi4Iyw
TADiDqBDWFxuHsCgtZwsfPRSrgfNZXrq/MR4pEVIJ2UvWPACBqqpVnFc7Wga
kCWhbU87/pQlAFCbhf+JrxpxhcvKtHbX4CqYjNy65SwYL47MfY4+W0oBPSMD
6KioE022YeF3llP9yIvc/Irved9q9rBNDy2k8VVBOF40o7jGRyjF4kgDTYo0
nvbIeV/gRHoa9A7OvBwVUtiFValy8gcN/gGfwUD9BTSCrC7QCS5wCEek0m/9
hl09QLQc7IItNweQ7bOMVTovC+9HyMy/nZCYw5ixwEh/j+tsKb0n3zRJAliX
LRE81L9CuSX9Jpi7HKuQgpWGRhihDLn2t7NbdTA8o6UNw4UCasUpj63y2SOa
sD5xnjQIPK73K+mMW2u8CH5RpYY3NlgKepmWWX5hxD3VPiuiXhmjNqU5Mh9D
RbGTZCAyO4q8sYV+Xe2BB+lJRh42qpU+L37NH1O0zUzeStbWsFc2r3XEqlfe
jgzyM2N/5yxyFF9gSZBEjoZXvRaMZF94ZUf0utTaLI4X9l6BQdsdp1UgS12/
1fX3kJPDJWBrZy8IjAnggGzFz5vtbFRZoO273zeOphZ1H6v79/l9IE11bzyP
sqOkvasRBJd/WzFF5+S8OOfqnVeKFfCQDMSe3Kp+JpZWFawiUNY6FzAt7/xM
1qF6cVsSfxEbq5yzrbwbq3PybUViLhw7LhDqzsvZQJJ30vgsy4F9rv6YuKFw
66AZ9m48G7HXRrNHLboRtoo4RYo7xQ8StnVqTc7PPOfBZhWMB/0UKYthlr8+
zghCEMetXtbRWfrgfEJMbgtUjCgvDU5YT1vYuoXWNIdECzDnju/SV4P3UZBs
gxyTtPpmxMmBKMSGPagubKJ2pIFCsVe8WBmXzsHa8C1RV5MRazMC9g4/qv9w
ZwtQPIeIl7BV71J8CSRoYxlJNXvGkaAioOtE6G7KDiy6PNEH5VVh8uZV/uev
8KaMYCNQZjjhr56U6GiE+Kzy2rEdidgf8gXo4hlQq/+XlP5wW57ZzFEgp9nb
W1LbN1lEU7Xkq8/jzVPAgiDFVj4XO4eKlE0qfYE9uEh0s6808M78G6gHzCa6
JesprlVfN/2y585YbE5WiY8ysYiSYPN7Ft8BywB/cKLiEAVvr83fFBH57LCL
ald4QiGzBepGBhA5ZO5TFxasOqPFFWJQgovDxfFJwaez2KjfHPAycgmHVlTs
p6CYAIGR3XBvi29AvQqtbyHNAm7bkywiDN5/OBypXGLevNU1pbhaZYn8TUId
nhplGumZNU9Ho+ZeHbIM3uqwQ/1+IP5D3dVssZkgmBmK7r2vCx0SlDXCOgye
EYoR8hcZ/6Jme9K3ANU88L5e97U6HDdqZUo5Deb3Q/g7Aj9kFPSSWw7ZQYsI
K0VM0ZZJTm+UNCh3p6P7JnvCiqDc5+WkG4Y7PBAAfL1vkXlOqi0FpdHxiIhA
55zTws8Z/uBpmCzwWgh+Vk3ZegBEZG4UJ9BzRRls4aNuFN0Rkd+PpbhPI0vr
lWZ57l/EU4EDCDHDgYP9QcP3rNdvtQMgZysuYr/UewppHIsqIXrtPzs21UCe
Fg3y4O8sevIMDo+E7qhzexo6zMPmZVSs7Wz3QsBEa02+xpl0Pc0xF1u1ELdI
ZzdQZCWcvm3Xg1HuMbMuYQpQbOK3P6nyh1u0uRt8MkBtaviYN2CwmZQr8spZ
O/gZQqhvmX+zxYWTS0boCO7aeH3Ldd4GOZW/siC5XPkWvkWW38RVDCV7hKl1
+lCY1/GbqXkyE6WarNjlPjBdCpx22Yuw7aa9RFZ4gX1qxyEsPyT/+PlyyhU+
u/T2mbdUou82Fd9q4aT/JrKxS7t9GfgOY/FXdPFihB2Jl/SxyBIfd1ae5Mrb
nhPCpg9jCS1Csdc/En72MrljOSayJAw4unavlmilrXnujneEe2NRhwGDmBCA
TPArOqUoXGxPVYKCOGB6AmZLhYfm0BQt1URTigt2jv+Kw8lKrvO1ePaebCew
Ebq8cHBFNk9zm59i7Eoxy/6mhbx5ttpspvzI/MmFUuWYr6FnqhLS4E8GBL+g
WMwk6wNJ3LBU8ysi1vAXc+xwhUTOk2C0B+3cZQbGle3WAc7X1u9PCA0ue4Gr
yQ+IGj0zQU5yWuCFNsVpLwhYjEb17s61Izm+ItxbC703HxODyzA/XhcgV4AM
k08ZHw0QZVgJ+uRZbuGkaQ8BTF+BhVF177g2vk9w1EQIsFZY88kb615c+fOf
MAwhrUbuQiNysQZcgZjvkD7ToVVDyGQb/sJfsbrzcbPbLVO7S0WF59o/cdq0
AhXObJiK/d9W+upSacOnxShve2xrw0p93moCSKtwbaZ3iiFeQwU8kcReodkQ
aL4PKryRpMybUE0AX8OfaHwng1j/JgIVV3WnmwyXgwMfOznCJTWeywSzs8bh
Zkm2d/9M5lK0HpGfn8zfOwc3OGtWIVdswCzLTXmNuLnsvKAj06KkfHl6JeE9
YjN9ErHAgcAUOziRZ10oMp3jC5Vw0KsRHR8aZK33dOj60xGLAxKgd0WA2p1E
nCcGDl8h5A1h+G/ozjzHNDvD1R3jMmxdkxNIUYS0LzKRnCscFizlh7AMYG5F
jrk2lKC1NEMpZqHamnrHB5TUNs7OELRTM9yOPlqUikEwHkeBqCaHS2rqXKF6
DDEzXCdYr532jFKezWKYHXJ+Nut9/FN6JW0quhsoP8rKEFpn2ChrMlO8fkNM
0YLaJwkNfsWyc97PjGb93vns/8/NndKorv7ppd6yRVLg9qbXIVrUAQxlOZL0
RXdTwSwcdGo3SWYS7WTE0hbA6mb7Sv1LvWalYvF9jDMijz1jEwTn2nV+oCGH
yTGqPgSFN8D0c6VrLOE6YiLcAA1M/0j9S9bILMK928yFPrIyzavmkkomaaeK
jP5dE5izwyDfo55efndU6w8Kd28wtGgfz6njr66u2Hm+sgDz7xe3QlYEpyCB
ayLO8gwJR8DRwZM2C+Xu4SCb4s54Kp4vzRilqHMrYPFFC0krht7gOcBMF5br
FSlswNoADqgIoLCLfEN9CoxKKxzd0U+GY6Y9awtKcKKmA6Jmn0hyU/v+4X6h
jWHPY+ECx1mWfuSMa81fSGLCkHeAyCBsHjNXAmhzXYfVHgMHRp7sPPiZBgmO
gGl2VrzwefcX9sxKuidVwkrBC9Uql25uIMNqtdsJk4GWwpU7AE3/oIhV6Vcn
7dNfJhMusV7IUdiMYGMAotT7hPfYNn+d3cTAusjrEgWdjJ43DRmptbqbCdfP
P2Wl+ExiXi7jfBwC3l0mPw4G6Q0M6AeOaVMskTUMcplc4EtIRrQzV4yv15Wh
3yota9E7rFLcFWHQoYT6THNyOKmxBTeUwtLI8pSnLQzrrNWaGI2kk319NIGu
t3HETEIUcaajtyV/AwNACGMwCEZq+9kOyZ9iREc+sn8wBHXpWZVG+yvgyCBy
JFhQa5QLhSgLV5D9eqWoWaJbBbt15YZxlc42Y3LzVOwcYg4TeYzu+OXQa/ks
F3xYubzF8RO7M7guij9byFxMJdfrgiyIe3QlMr+SbxeYaCuAAMVvOU/Lc5Ai
4bqTbxkfulxTvPlwkkmAFDWWz8+LIsp9fMTF7ikcWsrE2stywy3UiNGMIa0F
4EtJRXUIKCgny4A8BvzEz1fyxDGzpc1SNCC+yV4hBMXORxfyk50fb96GTuM2
VVGJ4w4J7gPF3gJzoUQGMnD/TVRwUbVh1JAOVPqCjJPTg3tKQVOXpYVn80D+
Bup8gMnMhABqTe0O9Ou7hWhnVpeRvs1b4a/tDSUCB48CsCWpI0mpUAl1w4x1
6kLm3t+bHM3XwC5dJbuf6ixBEjdPuZPuUU4BUFwZsQMYrwboFIzXDbXbXFCo
/hTBJroYzfS9ndeiY6qIz5q545hrNDbf3F5SBNIJMPfm2X/JgkCugRfYJyFH
0EA01c+bHsOWyqzCdad7R++IVW/eKdTBMijUvcpSezV/38KFpZiaYBCSfeK6
A7cOtC7He3x3AJq+R2EYerutBiuewAfOIwGYmBqyMfHOcg1AajjK2SUkjp+t
Hn8humvP9yaOsF2RDAJkGtKGPYz4VHO2LlOxaywa2c5LcvE8T93OaHSzGNBF
4+5+HJ+fpZ7/YauLlq64ZcD6lPcFo6EhVhPYD1y2BTT/5dSwC/LZ5Q+Xz9aD
//ZdetVv1c5ZEzz7fdMPvmb6KkBmS69jmYrh/e0CrQk9sMfU7Z0Az4703cd/
DSxBGA0/TYRVngN8c/Wb2GLllai/P7QtM0Q3XV2rSNETNcW0HlQD2x0kA9by
IrVT1fmTRepNE+774UgMsgNgxTRmOeiqeH63V/b3H2FdaDudGM0oYykFmvnW
74nTLCiHNLXN7aY0fS7Fe0mHDYzWnWeZ08BZXhPHUl+/Td7erACMJ++Jw/Wn
2CGpq/a/7DSqGrnp+Y2df9K5Qy2SNWgudYnEwm+zAO43WCTCCXi8CE8rv2sL
SzVOpXwiGSHU+/HfpTzkrNMiUl+trctcLYmR9x2sdYZw8T29qdIfpIewH0R9
tGFe+iIZMaWYt+e55krPZYC4V19OTVT+cudhjOCqIrVP2eg6dciRcO8w64F/
kpjuyKaeaYhqEYoaOAEdwNApku7W6v5fv1OukFMkAORnZBVJG5Ol1yozvrBl
pDtHnWJ9yTLaoC+C59D0JVgpz/VXQwWlvO92T/NLZq+Gw00RQZkFxmeg2H/L
8ykWvjF2ay4FBsb53KetDT5J0wrHW+NlXafdNboaCutk48lk6hYR4av+jADf
HgsE9xukFaUrHgJ9fU9SbzPRxncKdrx8MRHlM314HaozFohpvT3AAb45qpp6
5BfRfC5SPxq+GBpaLG8Zi1iSr0oEICSb039nLI3rV+HAtQdOUmRJ+THnNDzP
FQFa4oI5UmVvWPaLGihrk6RSIhH9otc6PXwzNUAVm8e0HVdB8oiDUbPHw+AH
UU7taTYPxw3VHlM/VKw/b7v5h9rT90KAczfOcI2mKTZzoeavZJjJ6kT8/JkZ
4P2wrcDg+zyDOCi/05wK5NpFJeoEfDaZZZqO0X6ymIEXPEFyl2uVB8qzk/bl
NDtolxlIC3waJnkwQ2IwBRcAiSj/nCimwhujtcty9BbZccTp7PcNJvy02h46
xyvshg63Bx3hBc/jFzYBXBCXyRMu2rEWw5ofJS3GJy9+uGw1xe39rPeOhXcT
7uuoKLjwO5TA9wcAT/Yggj1PTfZIeneKsmvsocFJJRFdajG4cDnT83jwAewg
p+v5weSa0ehJesW4ZzTqA0WGh/yQL2nHfEBKD87+7dgQUaYWfQNjP8hhWjnE
OEFtt6HgKRZYSiYWdkWjDTgER3AhnQwyW0P9rfasyJPa94+Mocratxw9g8sx
Ffgu5VvHjHBn1nvCv3ExoTxwKxCr5f9zDBOkU3yTS8/DkHIv8IoD6PHtMLYX
W8G87w65uiYK3/hb7zeJkpkt95o/DiYDHtxGuxAb80NYG6rxiuYOk/QJ2FDD
xW6pViUtQIneWRSqA9cQBQjmBrTJRPCux7xciYGqn3KzLiQPir0egaddFyzB
ePcsGN+iitAYgvyrq6bnMcViKgqD1u0FifGYkz/CkXQv5fVppeSeWKJXSqiH
aES7FGKjySfOXrGI48QLszPzmc+y+8yqEmvpm5Szy0QzRJoO6DGsznip1d+u
cxvoepm/k57lYZzG1RhDrE+N8Owrk8jhW5RbmwtgDqevR8t6D0S9M3MT/5MI
9d2C/zx/UabaPkvb6WHCeFkVPnObObRWAIDnUhfVoW9QacgXMNt8jrki9GvW
2iwSFvUsianT/nWzp1nEvDFHKIXiYWXHjd/Koxod474FQ7yp5ldFL9AINVSl
nKBByDX3FJxHgOUdDfgYPOK91UZYD9t8vwMwFq21GIXcFx7TQtUdygRFi2d7
wfXVbiQYT/1t4je/Xg6ho91Ksrhx+My7Q+MZWDqh5uyXSQyFno4/IjovechX
oGcwC5TCelI2BWiCU5YO0tZMsutQR+dQArxBdqZLT4D4JzdwiL+RLBQwIhwu
yax1gr2IfWBBZhloDB5lj/7cSXijzx97EmGKEwHPJnepE+i3BMkFLPR0I86S
KOYP0eTU3Jq6GUnIOGhNRrO9qcu43PMS6PTW55wCHfHcsNtaQynnnTiLAmi7
T6xFZvpWM4YVFaLxAsErcGqH+ecRBNDMqhdp8u2zr/Yf7ntXamtjZZOLDJUL
do9lNpCPo13sQnrGmfTDrV2GqkM8EFaqY5lUX/HbPmw0H3KetjmJ9KtM9vRG
HA606B28RJGqGXxhio9gKlfd4P6/IpLb/cXOwWVq/sZ1iE/6Aw16zIZmVAIf
k8roLZyLdRbZF7gKRigPLs5U1OhZtUN59FTEvW5DiK8eShXl6VDzyamrkFw4
kVK8nAQ4LqfGpJfVdlQjCsKbMp0PIkekRyhjTTv8MJhBSrBjpgLxaS+8dsIw
2Ul1myQBD49Htp010pBpOFjP0pj+JIGonPjbnqTiLDTxrrYYPK9IMcLwpAi+
DHX8V763ik51T0nbscBPGygZu/YmA23q8IEoOrxFIAS+7Yl3xm/W/jjar67Z
8UWQ/RHtYHrB4sSuGO+gwEAkNYer2LJMkMPmHhpaqjPrAAzChKPEuE+yJxwK
KHTQMfL8IbmIPwW+BeJFcX6UcMDy4XFPW9iaFgN63tCuteItSmEGNoU2OIaw
azje7tofId4brC+fzb+7uOnf7DvA9lVpxTrlD+XJmauLXdsCamOh4J39QoKP
zEU1a88Yep6LFnRday61rjSDqcjMqgv8PQuCttTHwbrF/jdoQNQapMSUnF0z
w5E2eTD1qRjSHFzWvXexgH6fJXuaOIPxD31LegOivk52rC7BPGj9pfiHXpa2
nE0qzcj0kR8oN0hziuXF/Cg7i4BfaOYLZyJ0jnI7KU7yl6GOQLNR3DvwYeB3
ShQf6AXjAQ6gbkWB8tr9if7kBF2FnuPzWVjdn8n90W/xHOBxshmSt9lgWy9n
94JcvfNT0Ty912vwmtLAdG/dDYc8kId9vln6WRkKjS5qBHFyVikUans/nBKb
S0T7DSy3mYsBYKovOoZwsvQUWmzp0QJgsJoVXh9dZ/YaQ9nQQV+Whxywosmz
0PQS6T0MyaM3kz8D5kZF3c1aJ/BVsEJq4uIjRpFY4EB4KxRXJY6TJZfecdHg
l9jUqPP9jdTE1CF8XY+loi9KZoMDYyTsdPCye8ZrNAHxFzLhM7Pr6ZBTErRF
HDvX/93lhiS2uNYcyOQ/mxe04LpM2YZ+KoyQGIB80ZoullxkdyifHBNNbl1s
DB5DJRFJBvbsH/5hwkOkOS6Hk3XGt4arYs0Bn2mL2TTv1G3hWl9YqUYjrJyq
QcGnPYPgAA4yVE66qZEEYcrT23AaXCtPmWJ3xwemYnWw5UhLgWr+YmaJeuhd
u5OmlEBodH0OFpVMjL7ADIgF7+TQ5ClDsF12cF9JEnlu0+MssJLxikDKV7a9
H7O2nPSMWKneGN3x6D9JW9aCPdTpbB3e5ILTOaczuHGQ5IEehj9z8WwIMCG/
KIe9gDWVnZ3U109W+VdyJ7R+0geBGWleJcgCH40EcdhJAuve5HgfWmr5PIWj
heVPWqXip+aoYlOXAiqaut9IO5HYDWoedpdOkt+LSS/g9VWnikiNLtLo9WJO
fHbhTWQ+oco+VVcnwcQ7SYc6AiNo10xzqJPXHu9PqmNf0qjyXz/YxKSLrjo9
7lHJXj4t2pXRhJsDVFTIIBCtiHtfsAOwVn6fEsun9XV28GiGKeVYp7cQrCB+
5fE/U8OfNTZ+QaUWf2pixkrB4wt7DIsKKJphsMDRPfwKDjcGuQjYJa2NYVa+
zgwil52yY94KTz6QEH33i5Z7+dWgSgGLTbaFr3LirmnhrnvdBSSp7HYfJoGz
IsnlX25pR6eGjv+cML4dVr+s+38mUvdhIcacHvCULjwt674g+dWxhyWpws2K
eKuH+9IvyXYVE50TflIQxgU2XOGcXO3Y7h0QnOfUQfAwGVPeTUP3P+dyH/Sv
QMfbJp3dT2ZOCmEdaqKWVFCpb0bn3y9WXDDsxnkTmD/tGZhW4Q8ZQLPlQzhC
kWTbw8r24eZ9g9N8drZvmeuxoNhsQDwemlqWUPn1DE8bEBXRq5zPmYdEztkJ
QnnYFDNakjyhLH+hKT5NNksnYiiKYMl87sl1O5s28/hs2nMqt1Pxph5MUjeX
AHXujMPtLBVjJqa8rgJ+ClpHIvgbDC2NtCU2e5ipkZmJFrqkfNjAJXVA8/+J
MYEBchg8LLH1XizrO+UkdH+B8uUQ5yAfT3jdaVhG2MiOqy2CcK7Ep8DARr2n
XF99n2WI3n0YTOQFZmJGFtv7l4qxLQwaVY26L+MHKkYDEKznjy/S9h0e789D
/k1vFQn331+W6o8wnUjZ17Wc5Yy6tYyWR/jR2VecH70dGKFFGsHwzOaEUqKv
cdlJWefbMlVYJ6MK9nnu1L0UgC4PgmXbFSo1sregbtn3AGO9XoWNVgqX27iH
4i5p6NW/n7DAjwFmYGwSzFQauInR2h1hWs80HTZllegls3W4Hw1jGJugFYlZ
jZhUsImf2Cb2MZKwPchS7/jfeZRSzQAo5UlIvhAfhiRXumpLCdEb0XLMiqfy
rcXKwdriOilmh/9uMKYYLYN1N9KgQ33uxVrtZS0bVARxr029SX9ZaLjlFWrk
6Ua9A8mpgTWiSqA8GoX9vU50PHrTNooKnUxdycUVqRrUeZWXF+jzhmq43Vmn
XxC1MMDGNN6AmXnY6UaSLqdx4xJh5EKOcNJJBXbYuwEOxqvNzArMDxaZTcwq
dAu14x+cGS+pj4yp/vbfUKz5G9AT6ppq+ROVs+ArzYUnDKbhke1yBsu9xDAq
/XqkaHdnHiMqm8g3fnHVTO0y06ESFaS9Lp1MESnbiaypkJynM/QRitqmDjg1
R8nxb9yQIXZWDsMi9u7zYyUSa4bGJMKlvjXlbJxN4qw6vqCbZbhepitgI3M9
wUMAJuS/L4NdYk/yJj/M2bcTK4hPr68FriYptbaq3Fc8XqNcmRp2NO40wRQ9
zEFdcSYQcNyk5eN533tGpxYbZXmGgW+/TXRcrpLVmCZsG6I18yjlbB4gegsc
VsqVsNziK6AHNsZOG/Q3MQeSWQ1J4gmZ1LGSe73S5hE3Ntq4c+bhmPaWFNTo
TtQ0Dqw2pue3xVYiuqUYm5zN3RY1pmch6SykqE0UDsMQGO3LGjyO0QVKAwUG
kmwyonukFkj1fStnWIIFqBenRvYwok5nCJxywg/vGjeC8b1wbHaml141ySG9
fXadgs/+YquYHBqEQ2G44PSycjiU1VI4KDCvfx1j4hstYbtnmOrfDxPVe5Fm
ucissMz32QS6uUq/p55REXovhH2BU2Q6IIgAo2albLR/aJ9Ic4GUDXKtQ7If
mg0ld3UIOryEee4relgyM/Re/U0gGQ6RC0NjTjTgCoH0LyTvks8xOxX5domN
qXEpeQCDwWq6YZp5DzyIAC/Y4BY/MJTuJGUrQo1isdftsy/T5YW7SCsh5IIi
dvgE+b4p012tRl2ICCP5R5rAK4diHfH89g6QUQ2TYoarFzCfA32Arb7uH6XM
90CZ4uTkjhr+MweNQ5QzXtQLjlO0O83IKu+yhO/kJRqb11Qq26zlPLwrkkI4
W/A9SfjOHZpNh0S7D9fHSkGDdRcPeUyCO7y2/rRpCY3jmB46rVR/OHNi3ZRA
99bRvN1V0WHvHEUEchI7JdMaor7nyBQfwTyEQj0JgC8Ku1UzSggpUoDJ+rXx
iFlYL29EwGOGrz8UJf4iJtWV6E780CuTjjdwBgaHSxY+7/fBEq64EHAKvCH2
dWoDh8Y8wSVokxPWdT4g8cDdUjdV4PhNjY8Yuk5MUOYqQBKyW91h7AoENOxd
NBgEABQXWd162f0Hbq88OUwqtujryq0q4L9AgWN8EY0C4i0/lup1QeDTPjgS
U+n6gWNI4cf58aHseXcuA8XlakSlhl8DfWLJDnE01GRr95qhuCr0+UeHENN1
AbanV8NlCQ/d2VdSnIn+jrbtFfNEPKCycTkcdwgFZNgEOkO7fXj8zUSJjR7Y
DxBTtcCUGAd90X3Pq9Wm4ruiqS4n/Kv7vifjh/O6/A6Piz80ejcs9FXeqaRi
sPCG+ltuCD5P7caA2Yx5ZCgCgEj8Ysvm8xr6VqlBFC5t96wO1z3PMcZwmpKY
ZmM0B0wpAPim0n1lkpQUU5w6RbeHKXOqstHjQ6pl10fUISVk6AU8SoLF9heH
bcrbnKM0dXqUJcq03Kee9NhIGf24s17r9LQQeJonGQ3Feam9ntPMXDjU3cRa
iGhCCjn3SSVk2wF146hlSagQjtFk5+LmHp8ggrPSCUW2RlPUHLnghQEoAdmx
RGXN6AR21MNu2MR8sREVIY49SIdOYHXF8BhdXIIWvOToLbw/hiN/ThCaTqzW
KIwdVfRpSHGuj9DVC/DvTMKtuy+2foahss3t6nEAqxT+SDUAt9tQLzQInPDL
sXwHcQG7H/C9J8L8KMX9cPtFpewgJfE3JjcN9zsm7i+24pDj9O/kEoubqw1O
xD0+/BFqXh3OaNcvx/GeDFDbcaOk6ifIWbHgIBQTy1zhgXQmSbYqd4vNr7O/
XdAPDpkP25CDWpxUwaE1QVHQ7JwisgQF/PBpY+iPAJZmTVjl8NMfx1LFKJ+P
Y14L0eDP0rxa/jK7GzodwNuCULiesTOjMRuCVxGHe4MEkSr5UBYvKrCN+2wa
qctqArBV3QcrH/cZP1CHRY/kiC4v75oH86fDGmJVvaTfb8MbH+myyL2Bp74l
ixydhjbxvlSAtwD9o7Cht8ZheNFHtutfqOF2xjz4ZNPJ7UNxjxLtqo7MHU+l
B9tfnwd9BXFXXqmDbJ7W+uGVuQO2Sp4cfskfE2BCh8wt6PQd+V8X7MdpgjYX
MIkb2e96b9bL/GEEVS/7LoTlazyFWWU6uvXEhsZ1mn0GxSQLa8HMg6jr4w/9
OWYWLj0++YAVKqH1r6mzISdC+NdFgyiLAvX3qExtCrQxyqvfg/5AnkdK8hQB
NOXVfAPg5cv7yZzD8qnNw6CMJSnyVGhP1y0SpQDhUSCnGFAnhPbIYGl5nLLe
+Mj4J14NBGDtMiKRiuDgmMQpBskjcWwToxUgYmkcxk5U8AF6XVtD1jnOlV7y
wRDjAUAPwsQ6pqVEJ/sj6ccvNVHOOi0oSgelINz1eCBAb+BMUlirz7e4Ar0N
kEau4OkZpf1QfBQfMyWB4y/KFj4MoAUfW9GVqgLPlK72zYdLgIHgv0o0Ky6m
3QB0fEeoYEgbTPeksY3moB0wpjwl4YJ1WvEg/JmdDeSWnQFaHl04t0Cw9rqa
TOMi7l7YLe2Rpm0KLiQaLgL/bctuu7AUZUKm0GeGYgoITAg3LZ5PC35lcnK+
PPP1DwrpHuJVR/rTJpn+EszJBHLQCc9dotpk63312XgKpYC8+5yh07M41ljp
6GbG1s1db52Z8ZfmduXm8q54NwMa2Drj+XW8m47Pfk2uweTsag4EmYOWcZOr
IS/ZbWiRMKRw2Sq8WfDqK/Tb9+3c6sPqvE/DGalEMGeKcmv72px4HPQmBbVM
bTcoV53d5F0uxWjocSfQ+hOthDRyXtSKm7PJDFAf5eYtsDCtaAPSjedopORg
3yp7j37dMQ1lqboEQkzjVrClXputyP93ieBd/L9oLpQI/zcInBkxukt+TsU+
QRpRK9v6ybrd1gLkpJkc124rpCG3XY9Q1JsvuqXR/ZqFBkhNoXjybtbtZM9B
7lmdsp/Oxrn+3flrx7I5mQGC1qa324tFFM3QjzOoTPtFCSNYzO88hpeMzPXa
VijJhntY1zCUGErX+QsFDOCpUNqyKrt459lfyi+WPPrrZ94IAT8ym5fX9BEG
Hy2ZKg955ClWijXZ6pCRjB9PrnUu8T+HfAdwU54aahKGlwQTiVsZowlKymUj
sE3dSkXmuFhsy3EiexrFZ3kbjRvoqqab0TJVPB4g0qgc+5/6fFMF23njQJOE
GzSuFeEUJQIrX7JKiR7DNPQ4MIz1eRxw87cccusJuNi84tBMm3XMpsDonJ4y
WoT76aS4ncbaqgXeHma4htnDuc+fvXx8J3uCvJa4fhVoyZ6zMvBes6ohkJmI
8qQmwGfOKM7o3ELpDrURomb+5TQ/K8OS+ny4NQ1UXr+mRJ3aXhCWOH1+HsoA
KWniUnENnq0H0ZIswr20uYQnxCbPIFfXCT0eCALB1pROlu9YrXLNlJ1leWir
TZl6aIG3AX7IkECBp5FZTl8Ex3pou9uaNEMFPg5628Pq6ev7YbrZJrjaENpj
GmjI9/rdPGjLuDpp4O/+g7oesc0vz01dTsCQs+7p9b5lq2hDSpg2za7h3CGc
pS9+XcaXopUou9rDrGT+o7PM0SsJMYMU/XN90IAp6R5lTplPQmJ0gLmIQIRo
S+8sruNXKOUSXHZUdGF0wAykPAmvT57mn37YFWPHVhwJnDclT+8IoZDvQWAB
XqstDJnWMSTDI7wZ73MCA4yth9gfvWjUunQcHMDm4qTtNVM1XxuF4ZIC7an+
k3M+LQgWnNF6HST0TZaV3ms/aZ4fB2lYWPYp8ekDu82Y4LQAPRwVRlkN18DM
u5Yp5sclpOx3UhIpXlfP2ChtHEdhbDcjxo3pMIhqD44WtjuYSJgDIYktuGtk
hNZeXtiaVxfR2ioUX6EbTj6sWt4Zfin9OLz9fAaRp1IrrcM+r/t2m7yxyYZg
q8ereW0vKoe0h6wCcI9uQd1Ybbgz+RtH3tD4BHfASRg7bOCasqRI4gWSCS+W
fh1vOsU3rLCS3lo6e9AY4Pr0hee347zNGTMQvhzXLHfgG9LWDO2lXKa8HKe1
EjqfQeRszNejcUyPip+HKCuGDgT+utVn38y5f4KDSzVFSFka+1j3oYCe5aOe
sl4doyaNXSytrd7PB9sM2wjhVa9iBBGaFJFtesp3lQohuVa3mrAHOKJEJN01
PFo+HYAK6Plt47/MQAGzc16HUT6ClZuFpOP5NZnXW5mKpWv40+D1vlLvGZVb
ZNtwL1w9QJvJ7KJoh90zB3fZNBeWabJ/uj7L3NuSiuR7L1hJsk4c/uOxUjl/
KyWLS+Fj7Tfl3462+9Ezk2Fc4+TJxBDH6mUAmrYobKMA0bNfxGmVeUSaT8vs
slbZ4lYC0XUhwvJSC1Z947J6qW3SVZriMPF4DV4pUvsMw5DbcOqVt5pWtUkg
0drUBmtrQFccZ8h29cX4ATFKyaosp50CwpUKgaCbxe/cBB5XnSaF9Xl0O35G
e8qjBVPvPyDEif1M6xwoHypkTUk82ZNLbC6ryAhfH5T8cUI4h99rBdGgpJ1I
5NjE8fHDVAVTNNiyuCbI2ag9RWkVbFJaFOD5vtwcJdBIb0gJpzGxO2fLh/g5
Y7MmZ9LBT1HBj5i/5tXtOL9sWSRMBsy21VIX7lYn+Haz6hn60bpERtO+ZPD5
6KOhEycmbbtx2m9zUGF+La0KT6TB1G/UKGOL4pREpDQDhR0x6IAXFz6kyVFj
6kK9iAX8q2CqW1YLl9CwfwqlP2Kwf+uqCmJOAXUlTQIiyhBs4CW7Ih4HzL0Z
juUsxUaeOvrtGEpEocH6NyT1e1jlpAQ+dLUIaViQMkP2uuy4w0LlOvvArzn8
EmO0QMlRwVL/JDAF30BPR+P2uzhPRmMHHrZiTibNM5qvd6YdEFdb9JiB8sEZ
XcI23vhruh85H6dLeDgcvCH1LliHqP9Fp08C0dhKeNUojDsQeUKRmiWeGJIr
TfDG/Flcy2P081Y6TU6ijDuXwSDGxGt+KqMFHaZqgDWBJSzz/HQ8Jp7dkzBW
rM3aNoaDkPTE0IADTdFBIjRKXRd1h28oIebMlxY9nxw9SkTAd4LF3345KKGN
DOfdUZLzqHkeqL6MVyB90+t9EJemH430lfvtgKjNu2H2u8OyEYO0j76Eu9Ca
9qPJb4oDsadj/DhgQQoLQzRTIakJYh6vBuJtx/D4qfFjLcB7d8HW5Gos37zX
/prsRHr+T9lOShbNnhPak7R2nmm2BxhwvUY2PlfPZr9luFyEAbY2I3HSGY82
Oxw8n3cU9ZGOlgWrGZyMRJEqX1LNAenuZBhv1+jGY4THGXzciObRRQ0++KKl
Wu+/1EyRwFQLQAH+y0U8Hsr+qNDzqQu9McZ5rUVoHEopmMhTwr3WOTUcGCNJ
wXI6r6RfXRiS+wNp9/fn7PRyHI50iaeIc1TCafWZrlwQ1C58l7LdMV71CLUE
L2UAp0hljgAu7+oQiDsIKRYb+RY/Kzdo3cs7kvL5rwE8MVu6oL0t2dVv7RQu
/OQswFNzXEAs7vJycp4NN8M+y+aUGmh/e9A/m0wy4Bt1FlHY2jkUYaVXW/rS
OImSplhTGIu7bqXtcOHdpDKjwmndPV9C0rQI76u4BspW5UuN82JuE2OgAP6+
hgGFWd2rr+oLCp9fb4oz5jLswtW3Ic4/mRcoD+eWZtc42Rp0AcdFXSvEM3dZ
+VrgTDMA1JVc8S17LtVRN+TAZTaVaoUqeteEcXPuYXGpzkAhb5CW5gS29K9V
2pfyvGnUyVhlQeCqmqz/XDYrGO3np6mqsooHxFmOrMsEXzuB/RXn6m3FmJey
d5GvKO5p76HlZTvA85J6Z9KEmIYBInEGTPH2uG+iXH38L7kFCmRetDtbAP0O
dVc0frY3SHVatgfqAbIgtCpMb7Icp83Wv2qXY7sjCWM42jyKRPNUopYuh9H0
Bl0CL904zabe0NGu+QPsho1ziXC6j5no7/gflVNac4HhxTxnXYOKkXnkYDEd
x8Fwfv4UWv0LbpPikxkLp1CdTRrT4K8ZIYDbS+ARMgk9WNCZhy2vNTJ4vVIl
lrS8Euoe23ee5Z2ykk8ljSlNu3DNb2/8gfbcQhYy0HzHEUrU/7OlOv95o6u7
DVL6n3QAHhmjy5GrecB5a8TlEeN+ago4HXpmY8ZXkjeChXEf2OtRnIIvAoYI
xuXcQFepe7rtwrGpv58oYgHZxnDHSGOw62tYsfpZDhT8r6igfZiVzmVioaPr
+ncNM2we6BX5wbn8ITgsVlO/0sVqa5nduBEHTTQUsk/GXxHulGz5JfGDmlfh
y1luDkw9cfwiibv1ur+zf+6ElDYcyexKuNm3YvcCHcSHpnq/nS3igj7nejbR
ISRXFqM2uSJrzoCAISrVQCgtVfeE66aYc3zrw2STJ0y0U4DyoPYef6oFnENL
1xNUGxN+CxGvA78pUdo0UAO3iXOKX6KJ0ECuKJqxliN+6sbDYv4cR1jbRYZk
naPN7LQOPOZkyPO0NQQCmAPiVpbeZZ6xMI4dVyXpLmJatf2h5WMb8nMVgcxE
52LkrG2/BYCot722tXflJqLkLIvOFH9pj1nh3pJXF6zLarT56w3kC4gqZc+2
SXmHSobN3qA+NuORaFcAWXVROYmMxhupwXF8lo8KP88+SwGtseJw0bKiqZee
6GIBXFLEx/sb4hZhIHSo5TyvFncn/ZGQxn0lLr/xYM73YL7dVgvKohrBrcNX
hfS/9rRLtss7PUEbPDvQ+ZyqjfL4NhfUHkUyvUJYL2iZQ11AmCpsgSTQ2Rdh
SrImZgTIxcMouC/8B5iquOHUgT3e3s0OGRtMoTzpV312QH0STz+z4HD35e8H
yXXW0TK2h4eKzfT5SJwOu8Yh4jaZXEVvlI6VvtpB7u4b2+lAVj6cQxhHtHcw
p4m4Ch4iq5AWtUP4ywlOoZuqp5eaElNaIjUgol5kEJOJtNj2T4TWuKZlZN2s
gizhXI3Q7L+cVmHvagbIT06Qyvf70q0Fk7VKIT8vB6hNH12TeEXVdzahN4WS
2UrLFIc4rBn1aFxWk50XeOCy6Alia+r+kaue/lOlwXFMpoM+uYCKTd91vhUb
UwoCPDrU9i8X45mzSAx8owcZk+7Lu0+i82Jn2SRHHj/J1v8TEbeXQHeFWYqE
8qAItCekMm1RHTEsHY40TrPMOcUehiVt591ks9TpFl9GYx7ioB+2kS/oTmGj
7Lf04/2rOM5dUQ/xUv0L92YvRDC0pEkoLpPlpFQhl0dKOciQPi3ku5c2JPFh
HyyJyW5hn3Bk00xA+wGdlDQAfWgFz2fMgnECwjqXVyUmOaSi+RfUeMlsDiQf
B+hPIAEvxUafJ9OZbgwHEEKSP2ffasH3llrmqkoX+GIHg9QC71ylbFy0bbMM
CKwCmErbQnE+g1SXBHZ5yueT/aAud4ll6PoyKZcQqdPNDAYaDuLSc0Q2bnrH
aXI5LXSj4mscFmRYYRdF6lo7H7qV4nN7d3WT8xyWpFqTGHY8+6xdwp7QVu4n
YACl666TfnUkBQ1SY8C+qdbGg67XpKQFCDBhfXb6x+RC0pmDhfdEm0bFXEJV
+qH7hEEm5Ze8OyTIYCk+CuKaK5qilayaoM9CKctHb45WbK9l0M7WBvxP8rnM
sjFiLYrM9MH7jWAHk4q8MctWmQE8i5KV0nfpKfyvaAUK6BX6yL0KomxAdLdu
IfE2jiHzZHQYOauaQAL5mBwDwvQI0rVfdC8viAyj8YsI8BMffLzDXrN7tijp
2QaJCkUgYpeAIffYhFL51foA4FtnV2bfYWRHehdzHNVhRX3/56hZ35jiC4v1
KRpB4gCPL9JFKG2T5F5rY85p8FmLjlY+SEdmvwVAhLO+QsEWAqCVT5bASzhj
ntJuvUtfZgbHzzy+EaGoJ4CHg5jmiVCepRG4bEUxtL5Nd0rfg/uabxKj9Yiv
6Dh7xQMRZK/LJuO4c5UR0n2PIzav7gPYpglMqsCmI80QzDhGUn/27XGIOwzw
xsdUDBuLkSH26ASPllLfOak0s8zJLzbNa73t6dm4dTNgcxf6iYSwI+7TQI7I
r0w0X/KW3Wk4V1EwUe8FHVGVtrO1MklVgX9AYcNXAJomwD93Svoe+7vdRsm2
1MNuIycbMdH0qXR+iLa37HMZEc+2C3ZO9m5KVVcpOfLmtYVWhvpEEMuvw6X4
TCL2iYcIfsevV8MrXn70z5Nxv5AIqnFH2RpRX8lB/c4H3Kzwp5ewy3sP0YvE
lvOKUbBQYogvUnp56KuvAYH7xptO/jokwxBhPT3qWi7eEjdi+eKn7VL9GWoK
24xRjlrdXpRdy47A6LFLqKiThtc+dc/uCqZqw5jGwekZlwHziV2BQUIo4xbv
7nA6ELxj+EwPsNz+fd3Kf9nN+NynFWMe+we8/PDWYNxSDo+DpLzp8ejbtPvZ
z/O6qDYOBLwt3tCNRmjurxUkUzmZuTHSh2nVOCHXV1ljQPSHdzXJLd5ZJok/
gOBocPgfUjcfZNkwp5a8wC/Ept5XKwAbePVnrs5K25698jwDqXz4hxA+B8Z5
rGQCCv3UYoTqSAOrwt0=

`pragma protect end_protected
