// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HqwS81dBvphQEvtfzOuiyJ6SnWBHRLQVYZ6BTNTjIbSchpywyQ81ieZCHE3u
4WRh0lAweVkfDKNTDDRuWatIakADXB77hNDvn9L0U0JEt4299rr5GvUA4tMP
RxjQpa5FAJZgBiHmi76f3/7lXwzOMgtwyI7D9YLNusrbTtbI5kA/CtThta+l
0fM2QKbxv9IMLH/EX/ozUL8DjL1uTeNv0XnJ7hMwBSw56+waTOXV0KznGZmD
YHfFkkedB5RpYTGzmD4Zr/j7/98FoRgfxPBBlUQL8wCxvgEJK03l1n3w3342
ORfCaogEGooali8kPI+E1w/TeVt4hxHB5+3eLIMofA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LgxCI+y0nXmA60ov0TCwnpMzqdjJMcFa0uE0DONEne4Mnd4Ty1L2igusriCm
k6Ff06m5MgCs6PyaA786iEMhy5G7GBHoRYXpFLAzPLz/Tg/+NxkcBNpuEHwj
s183r39ACV0tYANeQo5OdilYK0BRa5UItAQLF4zZ4+Ii/LEjot0sSte0QH4W
BQNBhQd6Xr2xov+Kjdw4F0jD4hRXSY1FUJG23ID5CMspcVmOFZkJ22HWZy45
rpUYYvLNjRZZCsrQb/enZSYxASixaNPX/BMZYGvDYJ3LAH+xusNGQZhauQbf
0cjCHltx74+kO8baV2NbsMimHKRcmgv1zNUssW58uw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LT2m5tx5tWPWdZlTZKB1TOuxak/fEnU2STL7ugtA1xYKd+JlV5hi0DoFrg3A
UGznfE7CbhWzfzH3tPY7Ln+q9aCuMaaHx1VWQ7OSqiLQ8cwcmbytfqENaOX7
u5rGYhUlJKD93x5ZW1NpiSuDRdSioZE20L7n27a0sqfm2SIbcrx8Z5EE2N8V
R6lDdnyG9y/1lOq76BAJgnMh669HLcQLOICTgZborJbEs4iNPI62wXKlTlrn
MgePgKMUIzoNkLthJm3BGFNG3b3fiFAKH0jlBEd2DvF0iNh0A/QFt/e3ZRXg
Wdm7lriV6Id/zsLuMEM5leh3CSP5nrWKdxvlZe80Ow==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sJIv9x0lADzFntYLwTvdCvcaUmKaQGTLMZ2Kxl6DmGcbvEjwU8RJZQjTWu4U
CdRxgRsNFiRvhEUhYtypCCK7oOhev0jp6fEA0/GvYjPEUUIK22i88QA+p5Fh
v5C4J5rPXp1qI529cKLRzHkmWWOtRrRj9X3yHw3a0A48m15BbFI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oVrVZFkJ+vVAZCMU4OHQHH72pfqPpv2G+BBNBzgsniBdNbivslAZ+3xSPUmO
8xT44LkS1nYYnCnegtVU+wYwQPOQvGf+HQ5jMC1bVM181ad6vi+tjJ6RL+Fd
KOaoEm8t8XQON/7g2e//kKbIIbTxdqOHin+DSr+edyR9f5BnQJmIuv5/Wxze
xIJ4AksJ0aFKYxbZIjzPIYalnjpJ33J6dEXQIMb7d2h8AXbeNnkacHc7Rg+1
G/8Vl1CwFqpw7iYbhu5AeusKM6z5gDQM4G/pJ8+MTpCKibQV1m1GCbIV/rsm
vHvT0FefBCE8i3T4rEQ6XyRVDgABCKS3+qt3fAHtFmjcgvtH0nShx6CZrtCK
XPg0trGvtuJ/gUIwK+V6baD6VoxG144UBiGOt0KM/l+AdDpKtLrDk3FkP7Ft
bjvHqfW6+Xy0Jz3LYYJUNTJ1iUNgzphx7QulK26tG2vHmwQkspxPd405P9vD
PzLCCZPX1NpmQw48eUl3eVV4PwiLLdDd


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sWteH3CZIiiclPonbbUaGY0k255F+D2Bdux1hKhjGUciIDcdcZsz7dDrOmXU
21E4dRsHuxu8n8PE5vVFr460vKZVMxeLe+Buz9sbMwyZnjbNhXVoXbGh3bhS
EJBTK9QQ3imkIeek4VO/Kr115T+8qGvZ4o3MBPV/jy0VtyV3eTA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P8foeF/cCQfVSXWtxuqwrFOG79TdzNBTBGR7ZDCn2bLMQF9xJcR0tq1MHC/I
kR78eOx9kNdbXj+IoxEdJ7iYKKKMo9sgqjfm2QXr6xURc6gkzdxaUxUg7E02
Np8Nvm7CWdoxgxbE9TfrNhrvWXOY7zM21EkQ+gHxygRgGLzISGU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 55904)
`pragma protect data_block
rX8SnCPsOH9Z7tMLAEujbPnpOGe2nekCrTzUCzuiolcRIyotfvn1H6xHhHYj
0HLYJb3Y0oogOQRtHfoGsHvIJJsR+xxh2tGlm/PjQY6MFOsla3AiOZCMOSNS
PIG7OZ8GzhxY0863JtqPoLQYjyn1iZpA3GDkdNws+t+MlyRmetbVeJnBvoZv
rNFXeE0u2tyhvL+xg6L89PNSVMIm4a3iosGl9EZstu/6U1qF5TmlmD/wFzjM
n4HRsLD6sSXKu7TJ+4Rf6nqMwzblQUWUbhjUj1sFgHUttUd4PykNse9eFiQC
FSgqAf+UCSE0r6ltzHnp1YlcllWH3G68ivpLikFSVOoGEehhC8+rk5hE2x78
td/HpLrjLY66J1z1rCw0syg3wEyiH2BBNrJnC/7pNfy2czONhQScsztNDEtI
iOeKWcqOfCP4ihYN0P4kwxOO/0ZxpbbBabyw2QRMRB9K7lz9TQS3kzeqKvbj
8olwjmcRN+067qbIDUocYk/3OPzn4AStp6vJWWE4KZEnxDQhkUnAo2OqJrAn
E+CR6ftNRYqUmgjvmZijPJW8gewLAblwg7ztM4Kg1/OgKC77C997zfS5qZR+
LEroMsiX3ygpOpe/Pibd2W36fts8Xu1arU40BfAxdukvAhHxIKotlQKYJf07
x0ESyWayNA8r6daJTy6DOYX1zdflqb0pGVqiCrY36N70hxRHdCHDnmFMEgq1
8GjN+gXmuB/Mit+ICLAPhZdMeSMTljzU/xu8y4Y3cK0r7DVbCssJlAZj65Lv
VE+D7uSmtRcyeJzNs9KWEi3q/CqibDM/7tqRFeXIUXs9/fwOYL3N+wVbUvdf
EkMUZP5vnC1Ct0ljO31GHAEIcO9XsrziH3YpyYTxZ1KSqf1008JWRfjOd4fa
orBoTBktdNkUUG3SdkOHpeyCXmteGQWSeqh2slxn22UBsEqgVnFHTtFTUMJU
bkT77IBqZm799u+9hBbuJxYocrOLhMzxOVaYdFoySTHu/hIEcq4+o8+iQnNC
iAbfdVspipWfqZjg/rSPsO0t0LuQWL+DtnBjXiGzA/fI+KrQOoieHQN7xmTA
YejezjHkyUJ80c73lyEGWjq7CVS7Uphf3oYuuSorU6CT0m9OGC2Slko3Kwjq
RUga4u2KWtd90YxkIk9WDt8W7TsLpl1JbfmvfIv2Zns0xPsq9/6vgdmoY7hg
kr2WVTlW/Dq4tV1kKkODKgIvMkgD+OXenmvYAhTf325fYsra1jYAnONIyK2x
u/Ry9s6awwlI8+Karlvn1uHqo8/NYfmq7CKALCFPgaFPS0tsXFX5INIxxeD+
/40ilj9cNMLYSi/sKaBji3XWHYpefN+/qdWvyasnHsnPQYen+yIBTvQ4X5ds
ViGzGKfdmenIj/t9bUYXuEnrgM7IwnJvmHUGNT/j0d4tLZyMxUpKFBflyzA5
BjvKYny6Li/IcWIXy0sWyBDq0OVr+eT5mMh7ODYX86yUPv3DhPFf1eULSgOG
TqXSA0leT+9Te1J3HS65J5/se32r45sps3BBzFRUa8iCMa1VMFEuvVyJ+rcR
3Y8M/4aedICZLhg9kTTZyrnAiZoIomrgi6FMNPrrYimeRK843s/hq+T+NLNc
in98Q/qdNI4A6Bzrrx5OojZu7RN2swDZKAHQAaxYQmubQsJwh6ZAjbSV4NlG
qFto7NyPlp8fMd4zUUzoMPUIO7HHRIWRqlzsU9EiYJ3NMbc9M1GI0lNr3zJs
xDLG584X95YN8pOuUTsKfI5aDiPwlK53TzJYdWrNM1xSwKzzkvRVMpgBCSB2
DdKllBr4RDffAflP9TPw2+qoBuAmeFP6bR0uyYNX70zgO6UbG7QOjaEe1gDJ
MI/nrTQsyjinOQGw4soNLCR1iSSZ/b/D18YEobGpz/OgsweUrygy370SaUT/
HV1/aiIVqjlTa7b5w//96lwmbP2FEcIJ/aNG0RjRQKdXYJDnkJ46m5oRHd46
KQPouIbtqE+ERwIpugMyGDlzejxNC2orjxEUsGci3u7FXTQzZYr+DPk3htqW
cJLxh4+txmVoKWh8R0Zjf0tOnfgtBVgJkPx9yPAnDn4mzk4GL0QnW7CBO271
Qe2Ff4JcjD+Y4IgQuTYUDzoaP/m1iq1Vw7nPcntAxSepg/NnNO33XceJiQot
HSWyYMd/hhT2K7rbOvOPem6rU2RzwJ7B93722dKLJGjBL4qRy6HsQeioLXtp
FPZymTFPIiQjhY72Y6tD/P746fteVOdT3IZoBEgotBIwAqZEJSBzUZvXaBut
scKstf/E+uA1qkE3fIdrQp84bVpZVHSftPrn7wSvFFlWSz9v/c48KPvyrzzQ
XFXG4a8z9h70vokfS5z0qabLg9hLXJof+B8GBFyQ+ZbyKputRTtWXK5Wib0a
K1iL+K5hHMwqGLHMSHIEhrBPC6OqZ3G2DU0xRCL8tfQtIfgVUBqNqs3jCjDh
Ux9Uz1nelk5Z8Mhd9FFWcdpyrq1v7lVrIp1dTNeYJjTzWaybDVxFTMoHzWvI
inSXYEN41wbODlY9GM/ekIclm0+OHyKSBLCER/AY8bCnt6o9Ox9Q205Y+gW6
+4lyHju/a5X3zQKPiCnPieCWRzVZVmiynZru1K6mjVP5cFW/a1fbtv/+XXHW
wbXNq7Rld45cOo4SZW+JHesinqb73ardEi9ngw2psrzGmOFuFAnxmaWYb1Ux
STG/LnpwlHh9+xu4JLsANm1ZfsdhkV8jKUh133i/cz4xp6nZBDtxyt6Nwj6y
tQu11h6j/oqLDv1t46NEnDdffdn1MvECAJa7raK6ki1DV07/PYPoMbyQlkVR
yZj/c/tDnZGv5RLrNcVSgI35c4LgvLUolY5maVTZCuTFWdpxgK0cqOBssOB+
nDlYvLr4dGaksKSjJvOWeULRWT9RnftWrcUqbRjGprT3UH4f9xfqGn9mjVk3
4eledci0i3e6cd3LgoqeYHBABWzq2O1XIMk5/MOzR7eHUHTJDH1niPlRAzTu
LFqN0XnJrggnLHh3AFOZklFDiRWY05TgNRKyKPR6t6/0+ej0l+MxYrX3NGJp
FZrY5C/5tZVxVAwBlb2iucTu0+4uNnbGkJmSFGxGah9QvDjx/kWSMBoN73B+
G11MLZ3DqEY6aih6V+YMBzYcTeDc335w9doFeLXx7g37tJL3TSGIgvD/vs5a
21T2MQVBeHyHKNtz2s3l9pp7bPZdgS8e+IycfttyQ2aXEqWmw7a1959RfTAb
nTlQoEYuYmgONpgxfsR3TCoA2Seo305gonaEq5t4lsb23+GG16UHCYHFdzgB
4mo+EsLpz4e1LkIEcZlavMX11MLMLBQLG6dJauN8wMDoLTNdngwePrsBlNil
bqRzv4sx1aPxQlD65H0f1nMmj4Er0JttGcrLY4evXmmKOz7Bh4CzNTB/jL+/
EPbZz+IUQc6laizehgsb8ejb+Tl2i7gOOKPPWz8RI+7dwCvzsxyVKDkGWSJ7
ijnxHSpUk3LTJHSslV53Gf6/Q6Sdc7HNm2AbvN5FC3//ET09I8Whc+uUqnsp
/R9C/FORD5alguS86APRzIY6xuTLCzRyj77qD6Wuu/m2nWMPUkNq0dhvSvA/
bfTDniTbvbkNJWrZWxVWzRYeoVFR9EPIvyL18xnIoVA0VYZyRXF46m+Xvw51
r+u2cm2difIDlYxqYs9JegtSvErRfCj/0rAKwhC0Nq3jA8oL7oL+UpJpKe2T
oxf/Y37c7S9apdrGbnfWGl7YCI19fZHi5pGqBFJfDvp0DVjU8xNw3vH2zbro
mIZYKZKPiqvBn3g+TpTm/6lFHpcLd3xnUZPSuXZqA9fbc1Ch3nAa8rzHoc4W
elrehzZ4ei2+iS6h3UNKSWoWDc5kEvon4JpPjFlb13ZSNomxZb19Ved+x98j
VkxyE7z08ZYlpF8hGfYFXvQWXZa+HlxIvWUv2QgttAyWzzBnF4I0Oi+vQxKk
ZinFbE7qu8gVMpC6qc081xa1or6sVv8Zg6v/P1pQmjxLbemBok5gPiFqqbhj
oohFqufAcYhWRyPqliTkknnju6JBqUvEAl5ao1rq1qszO1nf7G8Ut5igeZ6I
kfSMpkIqGisB2y52T6Le2pc6R9SKMXD8t3M3y6BysyeAcYJ91jpfv/1TJgjC
Q30cEbIVx9tsazEs+LY2J9GQC29pfUTbx+51kmJLfgU/oe36TitxYNaMsRNQ
FbIWT3r7lP4OJaQHzaqVZzPDJ+jfl37/DK/W7j1f5sb9lG8b3aRD7X3bQ5T/
xcQggrOe989MqNEDmJir4EdhABFpPikBGY4MtaHQPh95piJuRaKAi+rjbCDt
IhxWFpfXjGaKh0PKWrkGROaF7GsgYrrDB+BngFI3Zs+oduz1VmPlJGPZIzYG
YWDLYci8thg0WXr2fN81DztddkyePrdcNC9IA8dOEz/gofkhLg9nNZ5waxUz
GopiT5dj5TklduRIY0zDTl9toVcgWq3oomiB9ugB5L26dekdbMhG7sC36ls4
DzxkmT/1G/hEsz1h/ORVqj72LHbgJmMkVl82pKMlI9Yp/XdlIwRCj2LkavoT
lyqANQ1Uj1eeJgHAeA736dasuRS0W4XylXpYaPVtX7IebLj3ACVLCQGZmG6P
euHX3UAvqFxbLxobfbGo6IXkMJnbayg9XTwdY4AK85D0F8bJaHQ6TMO6bK3y
89zWn/oG7ZKr6hJRon/OeO7+vVkZoPpzHk+XkiTkTaifNCg7jaz6BjlRLJud
/AzA5Kn8NPPYbt5DSfvYxEbfKCaeaq3OH0XrEKziCKpIU/rBfFg3dSJO/B86
9Eb6sN/gSipSgcVOoI2al8k+TCo8jDakzZrXk9/o0Lq2sZqo9aJaPR9LdoP3
i/IM5ZUpObqGSA/lNUTAs4aZbIqQnjmw//aYB2S5+WZckTw67SosvJnlV2iR
2tqbUrDAjWb5WDMETm9xVEs5B8JiO5etioEh35QNsan0UfG9S5uaR86O5K5I
+1p76qO91Q3Cu3yW35IP9Eg68F0oOZNnc4YLu+YlMGs0zhx8iTv27PLI6tnR
Bq+p/1UjCnQKBxcZwK1wWHHF/VjRskqcsBb6AWMGTFK0L8FCkKcFYvKPPn4/
1Ji645GJj6pCJn9C9x+IlnG4EAj+UWc7scsDz/Axb/HrPuy4cjzgtvK51A+r
bmHs85nqk5N5LoSmufkYlUGiMpT9NSwzUVOcMG0rLCSr3LiWRCRTkADrwYzv
N7inyGkrVpF/o715mK5G3s4+0O+1Bk2sBIqSGukJOi79qH3s9D4pllwT9Brb
wafSuMKTYdwsre1ImNUmyv4k63/y+mOwuFKEpV+nCig8tnuQ7lFOFdkfRaFc
kLJCtZdx/USwt9hYtZuXxBZGdbO3kdTE8+S0dgShUVc9BpHPA+sacaTNNO6b
xC6K/kdvk2YZ1XeTrDznaheEuax/VkURXR+8F4n56I1gPWV9WYA3OhvcCjRs
+FODBal3mLtZe+9tKKhLPRvaQrSfjwNU69MJR4Cf+E3kijAjS09+73HCorW3
EieWV9LzAYaLLBRiigl+haWb1MoM4nKJViPIAlFqazagq7HU+AZ0iPHMbk2m
CzOOS2Ml7lD+LWJNA2M7reiQ4eqLVwMg15uswokOstxQ8pRFMzmA9Q55wXzr
dPgj0JSoYqluTLJ1C01LL8JRNUAaiJNImlsgIIEqikFpi+Ejw6DWLWwfbx5+
oXlIgre7LPDiWoamv3ByZb0nbD9Z0cLObYwerGI9gMTFd7o1Zfk4NQ/liXyK
RyLcALfh8UGUWskREcHQYcX4NLn7N5mGdDs8ri4U9GQKc+IVGdmsM/rvSajm
aKw+ZNvH6ZewhoFU/MbUu3qm7WYyR7iNt3enhXkOXKBsmefDfexoG/WGDSxO
kWq4ipo0UW0IBM9hLNBtfjXYAAoVM6dhWWhHkdVHDsmvzz7Lq2no/T7HFitu
fdFx8MAlHDpOlJztMFWa4f2jUUtl/Do77WlKtZhe84P1eNIRt+MzHmrwyW+n
rccFipuclYJoFwGea56wmpx5prtaySPLO/0M6zTpbtkiIUKWePokz5Ity2VP
X3Zc+btJiQjwlfBmBo1qkUo9PX9WGziuvMjMqcz2jf04kcKwcq0UDvU6DCeG
HmmRSIFJFtW+mZhHJ/xKBTb3s4SmTXQt+VssHZTJTd5Bjnmv8CghhyjLa3Mt
+B6wT8RR/GoRF4iyc2HxOzecpwc9gWFVHa3GKL5z2JupNzjuCEGBw1CkBGlO
oPTBh7XtrIIgikNfOPxwIMWPAk9qzhK1qQQv2o89q6Er/yEi5eBuftyrUgvz
I9h1xqboQF2YEm4VfHMILH0bAzaNnNYGnKbLlH6r94zig4DYnr0Qrn5c6eLa
n34KQ0AIVSEbMpsOyxZ759fUDBT80QRE5usoFMBeocOPhcEmutILB12eV/UJ
HLUxRF2hMfcPCW73OlYcfBWhRcE1a+FJUm80p5uqA0lR41jwxxTTXkehwKyA
8BHNGfM3xLE4oBQmaF75fmqOWMk7BIMDsDJM/2Loy7oej8VSHRAdZeVh2Apz
zXa/2Owz5b6aE83eW+s32Hmt8j0b4ye6cHVpnVi/h0pBXGlZQKFHFdXzR6OK
K0m1+vZyEY7TYFVxRcO7BSH5YtHFDut17fzhYkzbvJSyQLWmLrtkmJZhhBYd
AVGmWMAaHPzOICiF0d9MehOcvf/EHK6KBp0pYMOavQeZl4FU7TGmvVQMF0X1
LswOJQlEJJJ2JQM9ZchRHq9KQWlXD3cDp8Alpd1zb0aIrAQNVI50Om96PbL4
RDIa+Fp4T8fHdd/SXsNQlmXoqctU4BLVcvtJ4WdPe3PCIS3gioGkOJ4KRP7u
FWWmL5flgt4BvFHp/zKPJ2qzuPXAvzH8mYvZQ1hxE6hThMQvqo4d0KzZKCer
fseQnRwkS1jfMouDI4iQ3v5aTOg/dUdF1zxeyOSuzOoJ71vSxADBgogWcOY/
G00GiQg5i/O6kyIHiUstlfors9XdLgYe54PBqrZpB63AgYDPhJSoM5kLJP/T
0rf2Ru/MAQij0PPYa2VXpvOTUDA8G/TIC1wEEQo/sSQA9tkhmExe/dU4Hu7+
2Fkrfj8x1Zs7e/PUTiiZXYWcYfpLp8TnEYpaAikqgJN7Dc5bNGT7eDbEkSlV
cFHhWu7LU6icQkl/Z+wWMaK2MSyojQehsTCblLeufJTT492naPKdTYL3DdNR
yhti3KK+CjyTUFT0IHS+DGrvs0kKH8VkJjdNaRMErO6Ah7H/jC832mUsoIQh
0gtL+7PNMdFTIRC2JbZ5rymFZi+axEo2+U1Bv2mb7ysO8mVo/dP0RW65bqdi
lZtz9rXC6vgwJUHWiSUdW4JnDNXp7q1H4q29hGN3Pu4REQKb/6Y7iGWnQnW4
VzTC4jhMlntzMJ5yqemN8yJa7Z+prX0iWRATDy6hPe+KAmF2GWubF15DLClP
8lR1brPgnq6VxqMs5c3SfcEGjpvhknMH7kNmUAKwSm2X+OoXpK0E7vesiE02
VoVLQAq80D8fuygKah2ZsHCFKxA/+Qnxw/DNP39KWT8+I/rFdaFK5XpEedWQ
bVK5ZZqXU+v2iFKYsbKX+2xBcxB4L+dhWWiRYS6OB5DCp1xWmKivTF07Tc1w
1RtDNnfWfA/w8rggRcH12cSPBeLbk0Pzivx3IzYL6RPrOW7zEbWzwccxyE18
v6vxM9oYpcB8PKTvtX/HOrA+Er+SsWPA0VvH9XXXXPyNZt6kMXNuY594g5zz
U8eUHnXnLtN6xAQjYThkFGXwn7YOSQnncbz6rWbuY+NA5bg8SWWTraIkixNV
0tw6S/8Vzlhcs893k4QwvqdooLn0HLe3WyxMx+37pRhwc+u/CBEj070blSAx
TeS1vx+SBobP6xMzto6L5bvirg717BrP5RdO8TZpH4TZSiTOIhjoXnVXT/ea
vrL2koi1yxCzDwTCHYMbvH28tPNv0OpLih7+yBLmUMQ1pWidjeonOdbio+kA
sFepP+tZ195ABEiYjmxf+S1PuF3hRLmA/3ahO7myLsPDIvUSHXLXLPIMZBdM
KpfZp9oeQBR4JscGfd25meZYq9NhQh72uMJ6+0YOGRwrTQbeK79hBwZh5d49
jJW7iuYi1edxlrIyAxST55F4qaAI5vtoEPe3avoQTaTbKNcfzc0K8JKFUQIK
i1WUHMALMNUrC7yZgZrmKfW9xslo3JyD4Q7ywJCiSZRjUCXiwZTjog2+BFSl
tZ2bEaR9ffcLKSrFzdDE1Y+pEkDZ3Dx7MFBC/h373H8vkLBe3ShAmTX8bSY7
nC4S9E1nomOjNqlhuCFU6TZa6h0S0DRatpDPGevSPY8egLeE7QM5L98XV3lS
IpWnCIZMZijRoFxDy+wgqKODR4oPSMStZQkRXKzExwR+V3Wh6qLl9tb/bpta
nSXJXTcnTPYsMWMUHnoS6ot1weZP6CxV+ee2if4XlZmDmvmS8frQOMnXMVaE
bpZQ9VVw4mqVZ6lt98b91ucjPOK7+0S2ZH/70zaD9r28jWMilRQe7Ke2CsLJ
gMSXn4DCPz9QngtDtWMx+d6uiA2lQdEPdXNnAoH9kz5AaZj8T+is7Za2QVUb
ITtGznupKBst65jjbYyLYPHGj2cc2srOFNFrYOUwnA/eNo/X2KnHPBtuv8Au
1LfwX3Crw3YP9I11LIOuCrSZEARrCdoAC+aqyzwQo62SFIwuv2vzx2gJpgOQ
o0D508eYnrZG57YpmuOWTBdTy6XyKl3LDHDjKmVCtBvvqx9QeFGslpir/l8z
Lvx+sIX09XRVxFK5UJt5qqVXz8Y90TnEA0Zz/x7djg7yMBKDhzV4M1GnOOun
tEHfzcrS03rCvYnmbnmG7uFfcRQKhTPGILqYF+TWNhEVA2kNH+q8XNriH7Yf
grBl4vNTZjB5521pjMKx933AvIAMqDmEYAyKqJ+p0eAqt8GT7N4CzlaVcUph
HC94SlR1ddHTTZRmuC3Yn3iFuDt44I0H1aCg9gpJgPPJkAPPBJ58LJij4DwD
XnWgYjL97oqyQDuszqRw+BDn/DR++L5n19PPi9maAVUFy4fbwQfdE+vjke4U
FVSA9aaemCwq9jM0/gSWGbrzBepcGKB/4Z9lYeR786KyLWmKJGojXMSLEUg9
ZRykgBHY6m8jfIk0o8ndsfO+9AczqrXMxqSVpBdxronJlY0PzTyvYNch/qhL
OgmOKRvDe7zTFO327E3V0LTykeCZsmyIuIImNgFa/Ie+8FaYldgnJfzlf2TL
PHyc+Q7pDPNLslyF4ZFYkccw2j49i0+RvQr98LQuZrKFm1ov900c3NUckOeo
cjWVvf46JYWF9rrfPkpZZSvx9hJVHZHjlIKFK6E9/GID8cxzP/S+2zmWQ26P
2EdAfESqzQMpA6KWHVszxnqlCBkI7RTVPTd2donDz7ZCBlVwAt+mLu7rAAw5
k4seKmPc/SbiOqiqJYqbuoSdXGqNTqIvtOLCdciD8FFOFkVIBlu1N5/NFRd8
9ICm8S1kz32pZIhdYE1b2Ad0MPH10Ndc8jRC3UG0G3/MzEkGzqRhBsm7NeoK
qVhdfp8xAK+SElUva0p2xSAexIcP+WEr7deaMztalwKpFdm9HmIHkre1xs5F
DG3sfZmRNgdBLRJZwootv51dBaw8DeRx6C20wDTfEQEE2OIcnqBnO+7SI9Tb
Xa2A2BWYnBulMWXv4KcxAbG6L6ZHp/zqW9mWnK3/oPijsnTZOTM8xxCaHJDG
D7F0K7XbkPS8O98AXKQ35TFpribyTlHdyUnDSyTyJ41q37msQodIpdln4dr4
PYUkHep5HEd8EwHumT8h6Ko5kqNTwPj58b/m6zEVeSoXTkvP57SJIvOyCpr1
xLGzq1r2dfd5vbpZ3y17DksJcseoJkvCJTdCvM/P6/ty2wjwMVHN/+LhoLwt
sxhZsCLfnfqcl0ZqZweevwjdA/u8WqcdlbRKyDow+AITL1Q1SgCKyuTlmhdf
IPgcQYcOoDm9GbTdUegxXeyIYb0CIiY0pHmwg4E/rcORZFNvTrX2up2TWI6b
PgJqll+w9rr7/UjyC1s0dIzNKE9+CyfypKYjW8mkkj0F2X+1hlwj6n+PqBez
7bHpj3/p0YGkFX03wvsGwAi79FjbCv0qZwJHove6Qf9Lw5X8x9/JO3zjKUTy
S8ESmaBTkNMk6lSTc0nuXr78WY8hKas5fO+TAueyG+ArKXewxvZ8Nx+RNT2a
d0cr0YUw3U34LVEhQYtVo3SHtpTUy1GdmVi6wdsZR2IPvRcuhe9bOFL68I8p
qowqMUoW7+M6ozxjyxy4iEMQOAGmzsE8soipj2hoQvtG3rsrmckpd0Ezk3LV
WeRrvOZdpwCSk177lZOzLCvQbhTrwfzLq0BhyMYXqqBwUU7Dzv3t/qA3D+AO
DGu7Nr9GFa+9ugsKaOVAZ7AIzE4yq/RfC48SaqRNQRbT8WzFhxoiYAuV2stI
3t1Y/MtN8D80mdL2aMTZaonXasl87wlOJFY8T2/QWKZ1rwRkS8+AvOItG7x5
z0fTGaKuzuNF1KlWZVbqgDPjPRts/5dCpCwx4NH9bQMMRFk80AVttjGWmThF
a+xVIocCNp/0/SB1anS+koXF40Vlqo9AGgASJgU7iH3eCbzI1Dmy1Gu22tdi
j9RIQoI65EBv81JIBdjexAiOgqEbCbBaF28FZmNPa3tXl0weERdMfpj9y42n
ceyjv8x5KRWWvNslw1r+s5tsbx5V7KnB4BGYbqNXjgsVHdL3ToVXw0LJF4r+
Z9Sj3hQABBi88w+dmxh9e8AjGNVAOQy/B1aKhmTYwppoLA5xfhoAzLAuvgCl
NxyIxVoOc75v7GfI5VatnbjP0e5P9jUO3AJaLBi2rWnOvV4x0NnHT6KWxQmb
Rbchs+rmw7DdlTnXCbnlHL8J2eLdPcZR5qJaVt+iWhfgKZ093Nh7lfoxjRzd
db8dVv4qUaQjVsJ721RO+SyB6gXxCn94ueAKuJyAD2VBTvSjCmbWq09DUVkq
j05o66FJtx9Dt+5Sa0BeiYvZcEv42HGWUXkkupOrF0opniR+7iUR+vfNDCfO
/s/RmUkLoVokPPzE7ndIlU0TvP+rj/ABIil0v49/XJ3cwumw9nzrQl9aHrNr
r4CvGUvgOMPIbZIoqMy0ZdWsMOhCzPFr526H64kIlowzalH8OVKm8U3ooN0c
DlkbWUDeGZsrhAWtPCZBNQ2JTamWtWGZrh9f3gwnnyB4XSRMn9l82RSO5B/R
ymbfTUg0SNo9y6yYAjqhBoN67hNMM3/e2PHWqgQ9HgVGMe8X/l+cGIkq3IU+
uOZ/anlH9tWgvpEA+bZI3/ksCBTIuZc7NDjJcCwR2gZqeQHL9PetC1zzlZo7
hd12vassZRu1tBdwIXFt5bl5+RXi/ls5ZiT4IMi6Uo8ltfqtBmoFstBWzKSq
7h/69mfuKiqHcDc0/od1jaYB0lTJ9QiYhCq/D4jKDuFee4YtmBeCLV/Yi8wb
DV5in1zhK9MKEryD9G3kGtCULZkWAd8veyIqW4CFEjsUScdhrXvXxXsXy2vv
JNmxm2WZpY9H1ifDUV5WRw8BujqqYwK7xdzB/pRM4sknb7ysc+ax3nV90yzS
atG47bnMYYosGefis6XdUzjSsfhSW0mgeUGMvh2Lxr0h1yQjqHSII4GTRZ18
3Bld38bfiD44H0hsheY+cmxOEPjYZAbICrxdjASIMBsjr0WyatR+LsO0dsEp
N0F2CuV1COv7JEYrtDTLHjg3nb9VX2tHZ1GitMBp1hj5zLXdBRA5PGfB1o5F
vrGxznvjkw00hYcTpxvLbz7gYpLkuwWfBWAtQaaojOyAy3Diub6zA1IF7PU6
NFYT6us2argTl9JP5rEeEs1FK1V1dfccIbiTEHy4BDOV3od/Dr7XU+Lq/2Ym
Eg1zf8zWbNdlHF0hRmec8XYQrM3M5lTMxeb1bJxKznoRvN6Oh54PIR73+BnU
0RY67wjyyifJRfK8igvGkGhS73fdvlePSZm/5DCYOmkl9juCwGkVgPtrbfrh
eshkk3h3jZy0uWedGphXoUIfA3tEfV7sfbSZcFypIrsixSg9zTzKL9Fr2tOH
dySoKPc+79MKdh2fsYVSu0WTG4MGksHLdWgyTeGElwu7MgaUYhf6523g+yU2
cL9W4gD2aTGcPiFAz5eRTr5gxGHOFdUBrtK6Z/vZPQtotU2P1tRLOtRN9mKZ
2f94TpH2jhO7Pa/A0s5qYwtGbUblRoZNwht6uG72+xzpQ/Hg5dVZJNL1sk53
H5sC7PsDVzafQcP+jPP67xz6qssdiAJFQE9niY8zEVQNcMoKzEDU4Vd9HGLU
7P9DPqBCzh8vap5DzWE/TkCb7Jqhjc783gskzqKhGm/GQG0zT3Kry/NGYYgJ
P3KVn+WalEpkYpkYuq9bq3HjGJUD31bAoPW22W/CGScZIL65fDWqsgY7Mi07
mNLaf1Z0SHzvWhWHBkg305RL3rVzTfmE2YobgV+c1875fCuFU4U1CT/Zguhx
/Go9h4JuXb/4bncXABgMaCXYFkPMteJZSMsoUs9VhNPvRdscl9p+LB3Kd2jX
h37Wy+YiINC8VMEXbqES4HxXEUYI+bPGt0rwy40hlQHxHOQVU51dE/PMnu/P
Q7/vU2nmU0HxLSvGU0OXbd+SHBmltrPxIxlCt5JXQZHpm3zrxqlK/E7M9QX7
djc/e+vuPzB0KYpzAoDOsA08qXQbOoScaOnmHqs1bZexK4VNRgCy2okRczxm
GFEXKn+MPOFpZPiNihi+iGp+yNd0HpdgZXr1T4swmTygLVylWN5vOZangDI3
EwWDwkZijoSiIEkm0jZmIKjisd1t64keh/mitfS/DTjqbOY18HlSj/KpsQ4m
dz2nwoaMLTXqIqdkRqS9wQm32bqnjXBAD+1GVTtqbYlUfTfSOuPFI6Efe+pr
uTVK45vPpA7RJeJoYR8Pk8K3ViUuEeDhwBEUPGfEIXYNGMumUEkNkhjm+nb/
ZZKVhkspKYphAJIPr5Ihn95oDixBvSuvw+p0De38gpkEDoHUTHkuYSQUPVU3
wsRI6iLilWWEIW5OVq6SaG6ZYvpTwMrlu8thtgMn8ABcnrZfY8WlkXNPRqKh
HK7BKOWrz5Ep448spiurUT6VqwK7yfxnrhjTz9fh45aPuVSXpuMedZT7j/54
49QjlGF7tEIEMo5PAsTuwn/4mSKl0gK6hLAvVLnkxewEJE0XEGjePnj0qMUG
6k02mbKxVXDc9NBxNeB3IMaD63WUgPHn/9VVfYiUNxfHuj4+U5m6uE9ai2To
5l/1+zOTIKAS5JljO7x3ZqxQ9spQ04sjB+WtsQbyxRrlD0GI4NbFiQrgT3gO
tFe9v5wymB5LPap6wxvNhFhp3F3WX9d+a7dwwibs9tvoT8UVNYtnQoJdMkGC
nXJb8si0MOpCf2blmZeJMlAoBXqnP+eOX11DppsJYjUHWmVp+mQJdbkIzdjm
r4f1ATV0AO4MuTt4UJvUMbrkRl9hQPGsSBWWveu3ki3dUxy3RylWlH4n+q+9
S9tkmDK6DylYaiMekBurdxPPSXD40yF0Qy7Ca7X5qoZkf9oyjpRRwLm6PGEY
UqUPz+E1dJVLdeAhc+dfbKiCLLm0dXsNMyR9koC31d24Gv/VPr5RrTaYYzDM
YFsHDyFqOg/OjijRrH/RcT21hj8R0LSOJdKZ9fPGtiHibFamuU3bQnOoHEWG
VPFSWBCSYdORS0gQWgxE8xVhjF1pzyveonMn2796VQN0EBmnBusfBdPY7ato
Se2TbGj+nneWpOP1Fe23EPbqBj2gJ0WWTp252QHwyX46H08JIVGxZSMgFljv
xQnY3lgTJtT/GvuH8Q6pLR6yF1EMBN0Q9CKkyiuQgjACDq0EaflDdblhgSQf
iiVPRR+8IxIWsMIZxWdEZigMCN2ll1MWj69udI+eS0FreZ9ngjMN7lRmh+PP
vTGZLbgSyQHI8ov6eKFzmYwPv/EU/qyrXP502ptxoj11d2KrTots6iCaQ9ql
x5bNW2qHfxXGqRtiHMo3m5L3MW1Kymx82IqnfsGsn0I6/EKFPVOcnWu275uj
r4HBu39P6SmNUL73G5tSSNM9Z8dOazHL8UNJhM43EIwv7f6X+F1rAMyI1Nkm
Av6QjFCb8+AHDpzQ2RmXumawPAyQeGspmjoiGbhoAJYi/3WbW9WcW4FZr94U
6IlNGdv3vV4AbbL+3X/ofJxaXqWR5Sh1z9XBodeVDA7kZR00plSi/AmFz1kD
Nwnh4bQ/4h7mzadfrK8wOpwJB4ZjgFGMHdAIGnw68J0YSkVCSn4aJRAZlmk+
75N2c2on5i2Orn8bfFzVa2lUbJBiUAWAyQjqLtrK7rtNrp93a1oAWI6omCyA
E5goudcoJiy53O46L7j/N1XonQWl2wZC5eqNVrjbG/dqD33npxWzdFCyZL82
TFg8wRaMui0UoGb4sfurg0ZOXPWwFhUjwFHxTLcO6NAtbgdcDNjkaRZWLCN9
4K6czPZqa6Rdpxo0sOY21iP35uI2LkLVh0NkJ5qHLYLCrJB1olwfjHbvt79C
QUNP1Pa/oURwsEUU/eEdDcuZ/JcZbO4lOD3vdJAdLrcC8MuGngSXZetGC2gv
kMncA1kP0Q2UyPIex7ffLe9Z0LbmG4FKkIC5lCFCw9sPmDzwNEDQIwd89AQU
1fXzT0BOvUXCONzSOSjbSu2zB6rvfJT/u9MjHWbyxNHEJW7YbFsgwJE6MGq/
k3z/2RKNIxPI1caES/sm2BPa3CH2kr0ExCLMDiMNGz+ZYU7R3vwjHB7tnBN+
pQd5HrD2AzmWJjEzSAJkr2Mk5EUIiAUfQ1JeCvGo+jsw6tQSjgKKYQ21YOQQ
RDOe+m+IG7CkWVN9/S1WpGfwXDFq/L6/H1/fn4pWZ6hF56H4Ly09JfLXia2E
rw77fQGNDI6kbq0gfRwVM0CeSQBClWo0CpbKW1rhivLh82Drzf+jb2AhZ9Az
Z8SJNzX7+5PXu3S0+Tl0d2Iyfy1vd480XTscKA1LVwWW4M6rU3GCj6ZRrUOY
TcCw+2/UEQir8lKEL0pWY+qDUOA/R0LCVLkLaXF/4/hH0BugHu1oBdWtmvCj
Pr3oi/vCGjKr5u+o8S1RN4wJXthbj6Y9rdfU0S/w/vzcJAZMVTwav1b46/Hl
VreicPkjX85HXvHbZfaSuSE722LoayeQBx1k8kALQlJqLZI3ncEG4Iy7XdtC
WNJME1rIGjLoUYwVL3jQIzagcHjuV5UhtXQT5oMF3obeBplq+YubVKzXGqO1
+7yJ+Dwu4QHDoYcqeitFyczh99TuN99FOWXc5Ehnxw/3eGPChfvpTV+6u0sf
PSg+dJA+/LFqIasqnyqGH1JxDf2MPEzuCcEKMVCz+dp+dV3/vWaDRre0/+AS
F1NmjEds9mortIi4K6w7ndLZqRe/w5oJyKhBDR6mNQtsTkhi5IhUPaEEnQiu
qDAuPKmAKv6w38NPkoGOFCb6tHKj/PsD1LN8/gCLHuX4+2DfJAnGdj2wqpMF
zNx5jUP2OPeR5suG53oiL5xQocNASB7C7zAJQH5uxvmo27e+pu9+SoyVHTI3
JjEAXwHWVpl4QWwgZps2Nq8At0EB/Cs6LSBUmDCcXR+C/9FrQ62RIMy90aWz
dzQEDY1xck7izb3iAFoQntKxhgf/sYKtM55yhvBSXtbse3U+zHCCigx7P+Xs
EiP6+W1g5ctIm4JRv63/uft61KHeYNzqsu/Aikb9Q/bVJ2cFArfZpv/gYYlE
98UffTLgHNfSjRnvObSqeV1WYPlrEsV+3DlARZxJcT3VMOAlerF0dPRuz0IB
1rhvpTKf4rk1+mOxtym4k08EGxKF/ckLi7ba7/iENkpHk0S9V0d7b8aQL3gH
RlztyOVk232kWrXgPvZS68fBAfXI/Sx8olOGijrE5SYgu37Lnm3Zsmc/0BE+
Fnav1r2SFhoN7iTkvtVHcFn/GLR7nZHvvxvTzZBPbspgTlF6A3SOfQPiJuM4
NSDCgvciGOnmPyrzGK5M8Kh0SA3BAJTfEjgUI2ch2ZthuPg+9VYrvsOW/9Yp
SrXOxcYMuFnxe3d3Di6dd+bMZtr3mIbtPUz1IeO1J8G60BwoS9KCRFcgJCn8
48yzs50blA/mSZCNdeRsrgSdgfbdHutF3Se+37cEwzQwL8huVJgUL+GemlW5
GTq4hKcsk20UgILcyW5h5RfckhHejwdkWHrZ7qP/w/kL1tTMAPFMNpqjfuv3
0fkChl/Dzj+pgIN3n5D4IsfysmuStHYWzOKeueps3uMMAUfyUxBHSsuBTbra
PmMu6VbfzpiaVNfVnxGWU0FZP52P+HFWxRzwIZ3q0YUeeP0Qm555fxmSYc+w
g5Ji94E+/Uo+ZspLyyWm95gitM2DN92ZZNPtdGSPMsMqnyJUu4YEfK285oVy
LUMd4ms+RDJuBCRZEe7eNqkNowVY2haqpv4U/7mup1lvZAAiaf8DpjB5M9mb
w62CUtaWqNLtSPT1zhZNzMULogkezMb/J7OBaAWoTZDWjKSmK9Cs3mfIlmMo
7MKL3MYc+0kDGwTzX157SUYMQAk5nihiOI7lcIphOOeGEFp1kFMnD1+fgVad
BK0/VCGxRs3G3eqpHXV4qG9iZpWHtVjbj6m2dsZ0epxlVdxmrL1D/yB4nP3V
d5YymQyBuFqdkSrwwGZQlEtLKFIxfyoVDc4O53ekKEIPP/EO6F2KTHIJ10OI
zGpslmA8q7rvGJGG8oRo/d5X23SQ00aqp66emTYca9Pgq0Fo3Qh0Am67w1KI
5F2CL8qVyOb/PpE5byF5LljLcIChOZdNCOEgL6SK66UFNdC8HnPUkozkpyvK
Mx0x7/4fTpPSM45YsRvz6MWcc6c7iLSPSzL1ElvPdNbpgeH6N+df7zeRb1/H
ITNJFpr4NN3NPsI8pJ0qBVsE7jG3gVO5ICY9eLu4xD3uNapy9TO3QnKJvELP
otOduKSUmVhgCTtb1LAjx4g//WYrvxSA2OTnoITUQGTG6OxeJ0HbVK65kVJ4
7r3DH2And4CGWKqNXArEhWLmLD1EMU97X3fkRofuBJhe+E4c6vOGRcyT1EOm
eJfWOis6TLdJgs/JKsSB1xBQHPQ6QnGqReWbdOoreYKEdJpoze2ZFry1yM+G
AusvGvx7jbWLGoCkrlBw16mywNGg6zw9hiWjhIECaDNMSUzdm/UOW0WHIsZe
+hnkyF1WKE0rz7dsQC9Ik+N9vn/QDsvHhh8ELMS3HbqMuOLu7siYiCz84LHB
hVGF7MbwrBHx/pVTrTnGSM0CSladTii9sr4uN0DVYPy8Wz50BfS11sJZFU3j
LzMrt8cq38RAxsK0yYidD0ODMSBS+x6nUIO2Jv7TCfuIihdqX3d1LH8uPtKI
u0yD3p6YTaUyCNJctlyPM7ywFiQcelj+fFYB7QdzC+UyFl79NjE5gGQFOamc
DY2r1AXybWHPOhRVyqKt50BDLAlWcq1WTkPtDgvNHZsqkDk1bqxUDKHGiujH
21uFqH6qMvaoBkeXSbFccrYyaM5WLGx6GWgkRYfyee1WoD0PmqyZHEyr2wKC
08HmwmW4a2JvlcIWegLfC44dc6aYO3+Q5YZHia2WYDyS0Ja11Wa+nL/OEkrt
f1K7qKMVpUDkmv1eQcRiNNADIjcGTvqMQgdxja50eYND1ygxxe6y44XmMJHk
McYqyVeOYCWG7eRBYl3XjP91LRMUHpuIATgNaxxWXRzfksFTPS7ZcOnShQxc
hZIqxsSOkBMIoa0YzlNg2KjA8jMkQAY+nAsyzTHtkd3w/dso2voGLis65fMf
YBweAdcuogPW7UTqMCcveAqdcWF0LYcYjRVFz8qDGr6WLwCpmmEu+MFCJXCp
SuqcoGQw6W5SsJOoD/x4GKsCBBPdmSeB8Xc/EjKA6fzM28ukZGseQeT5mGHt
A2gRO84TUs98BVPdSUeu8/jJUjEJF0XA81aLHVsHZ7EuQJWPMdPf9VB/4yPl
RcXtqN6QNH7xxG+cLNl6wgpsfsamOIX67/Kosmu6KmyclpQgEki+3KQU7dhJ
itcsqh2HEYiBx5PsEpIZXXO9t171Dbw98GDBPnXce0yt/igxKKzlnh1jdYGt
LC73rR3y4F3d3Bievxr/mhNHWCoe1WFCZ5X2Ysa1fF6v9B0vwIqJIcmz6Sdf
adOrCClyGJp3huKcSFsjzyCsVxkiPUYqv0lwYmWaWzmfPbKUxjUvl7nl3fST
7hLN0qG2Xfj7vfZr2c5dI4LxOT6ku+hyRfThU7CLJL1w6DIfHgVHHEByloMN
0qsxIFA5xqAhcS1g2f8EB4cRwE5ayJM8ZiLljH10jBp5FPIRa4PQkUEmvjR9
TVmrwN4P4NxCpTE7dMdZrtDJbnPvwfFWaNUC8SvpTM09Dru3Gqqw2MTQPNov
hBtrg0f8rE3+dJ7Gqq9dB3knZ9IdT9IJVnHvyAYUPJp9VzUAqjozRrSy9EhR
ijNnT7ulDVjLm+ZOhxJvSTy7lTskQhG9sqwyTllvRe2wGBbbvej9KaUs2Iu9
d2PTImqlBXgFJzYM4MX5FG4kJyJJxSULX1Ge0O46XNWXmVCEaVmMpNym8k4Y
5Q7gBwdq2KK0opUlHMKxBSAyxFklKGzhbUrCudxVGo9p285XvCKL5VSHn1xD
8as6fNCRI/Sm0edzUmhvpmIlaOYPEpKEN5s3bfPJYknhq0duQmPRU4C5kqiX
cB3CJX4JcPaOuZPKNla2DCcH5bvbN3osRu3xnb19hf9X3vzQqXK0oKMPPJRl
ccJqcNQ8eK8yIsFZFc2BITH4VxOKGr45ufhkX62kr5HCLKELjNR8IV+RYoMN
1+oyFv3n4qvpP1vBJsacNt0cWiX05J/F31Y8AjPlz6CktMOVNBCwqKZatoDY
u2Gj+828al8Fqu321lXsY++NSWxNsIbd4iTxfq8YGRyQ61MfZr4qfCzHtY1s
p9KVaNXRaAlnA+rbNY9bpeSYtYLzfS1Jpr1V1nxmg27L4WUw0hQD7m+MVOYA
tAsZBPNwmVkNLt0zDACZM03Vmif4QtS+RMBWutipPVl1/zn7OMN4Vc8g0SG9
tE5JWROAFnBHU+o2Enp5AK1ugKjK7HhKdCyBanZx9M+UXuHoL1dHYxQ+GEhx
KQ8us01oxZh64tovUcZw++UDpuR7FjUimojfcTDPfRKxP7TdFe9WuYgWB+/9
WrGwE6pvGn3ThFIeQRWpuCYz1I2lEwudYq19tjF0Qc8IxW8p7TmoF+PQWr7r
7HdAykSYeDlinP485/S+o5ptTgzdqhECeBbcKH1ByQbylH8Ul+Nz0yC3PzZL
apwzuA2ULfH8h1Lr4h3fN8NhJiMcMO66trclNOrL9v/33/zebbT6GxW3O5T9
V9xA5WID/7W3V63TZzklws/nkz686SGBdyMLwN3oV8qly4kH9U8USpquQCQh
RRCo0LhX86pyBLtqKNuCN4Gl/D0GCiLG2wT4WlCI9P+zKWg1DtWSOsGGAQbh
C/RfkUwtEdjLRE9LUmYpGWDHmR76qzNCAcec3f0y3iwWAGAjvGQrlL7nUx2+
P/0AgWsVeJ41Tjisi82W2KThav9Q5IEju+DWIliGgr4/VZnfde/VUT2hHQUF
rnL7bbGwIZ4D2O7KjVoJQ/D4qBWWzh5LxVsIGCXiFhgD9ygC/kpHH7MY3aXT
YcGs/tItpxzBDuyy6IYF63V/QNXKMks8KBtO5slJJ0T8JNEuGuxEcLIGG3iM
8E3E1xkLkBKhVl63Ps687XZ2bA6iOQvwtGxQjzSvI66bbYUGm6lsdinwYW88
SChMYoeb4eekzsnYrVV76/hEJHOoh8uzsMfwjbe1hzqXe60yMrcoJUHfX3sl
WI9G8Je4cHYOph0NDhjR+iclJJdsjvYxb9RgTbkShNgXqsRWknBaOUlaoeBL
FKqmIZR28Bf+3qMR3uvd9WdxJAV8zPIES9/A1JarpingqWPB+ha9L0gk+kKo
D0eEpul2K9GW2N0FuxsazLWTEUIXHELW+Ll9fDC/RhyVWJDplgSYXybkYgqB
SJVtsSeJdPanLsIWExra6L6ADMUVlsHvG/gR1ikIhg2K4SWKxOvMjtgeU4L9
Us/tlj9+FmPTD9w1+3vmXajUeOYVlBLs102VcWUGMEdDz9JR8zcw866P3gem
fpUoAO0IqVEcADM9dYRX8f5Ii6gHZniA3lOHhs4q8O2p2fwdsmMYFBBG3m1p
eQKic2+merML3r/gYT6JhZRM1VAS4E0unj4DORfA2xqgVAEgiLv9zoPlxbkV
SjVGJ4pdkAo0LWP12WuSCZKgwFUUeyGTHgUrrLPcLBGXtAm8ICqZRAnE+feF
pFCWhdOUDpvhfzp7pqjcI/2q8YNAaoYZvTE24NhKf/omqCdow/taiQkqi1Ao
p4zcg5H2YFXE+fBXHrik7vwL2OVqEMbnucRCm5aVTj0KZWxi17KBPnhQNhtY
er9YawT6bxu0gFXdUSmUMmhJpEZYwJ5ovF0QcTVH6K6n9fajhW71+StLY1O7
WzMxeHkl+AkUA8fAtYGfOq1njPOd2HxbA8kMiyvZIJ4lWHfBqSCGChgZnHpp
KafUS+H4r0I2o7Zcm6kBVdBkvLedSucqh5gWBznDTs7tRWbymaWOLiQsjoLD
MV7VwtbHET8K9jpg5ZZSNQ7j51IFFD1sHkSz1F/qLzUy9TQzWgks+MpgzJvW
naF5nUU4hztAUohEZnpBY1pOKIBs/jLjGyiC9n7v+SDlan6AcUApgbu7GNBT
I7P7uDLBcSp+xsGWws3fK55yRHbG8Ed8ulO0YQI5UUr3ObYXXBY2ykVvJhbq
wd3bC931Qjjph7hKMjcPEvK4f32jfmAl/N5HSve2oi6hFWMDSaW2nsfOZ7sF
WNqmnIeTPuW0oXO2HBZVuEO/xSGLpWctbvDB478cR5NAemyuQBaYjdoO7e3S
Kk06vMtuLaEL6e/sJ0w78gs9T9Kmp016DGV61ZjmKu94UWSzOX91hvKO4YiY
yaaDqDmaRFOR1Uq1XDxAjAh2oP+BQvKgTDHuqwBXMrdoIZ4a9YrkbigoTGJz
Rwmpw7tiyGqUFamjOok7BtK5o/LEIKOLSkXBjU1W65uqTWlpAWb21KdzAW0I
YwP+7ChgK4ScOmKAE/AUDIOBauVqzBymw7tzq+gR3WtABHG7udMGyjepc+Lv
Nx1sHSEfZG8L2vIqi5doS+26A0zpygHONGJZ/VM2tu/ZbLxuTnM70Gli6lXm
dxzPpy37hpVHitJoqRKBp43pjy9aXI3OwgMY4iphSt4H806CclO+jVidv2Kj
vNQPTW31iRWNH1yay/+ASYtHtIqf3FRt1kKNJuonW/gWYX/pKe1+AlXluA2a
hZefZgvhqwDCf4cJlVofdvMe0wLmbGcJsMjYKpkozPnitVHkM6j2nctJ3P4D
9IAKiUKmRy62Vg/sUJkXp+qweJD9RFft0O7KrNhVL2R6mujZ2kLgWj1Lxb1q
t2Ne8RIyiPSW84d34epaU7q45zVZ34vRqNgNIZhWOeP8NIDcIuUatcDauKZo
GG8R2vRUyfyYiiCxNWFdoh/i9zVKyugHU/PU5JBpWHC/3JloWD6KWGCqvW1H
Hj0MV+AiZyMpudXjoz16N87ZUz0i9HIRZAkkDcBqQDbpCYHVUqb3jmhq6Kx1
SINs7QXbctsQYcecWZluDH0v03yJ05IZ9KBMovTGcNycOhnlaPuzgLmqp8UQ
jLU/MfTMAg95xwhR4P9Cm3OV0n+d7Uwr1OYZFLpggykct67VF3j9Szwqei7Z
k+qu4KKaoMx9odsL5JZRbaF6HALtgDwkQBHGAmHwxhJ6wuC+i7Vjp4yzzX8O
MCyfZ3S/fgLahBVPYVSDCXM5tTmF0rWHKsg+MD3WrYr3Y79qYhXDtJ2jW//d
tWhuWXiJQRI6vhJ0LeQjtJW2QIz11JlZkzo/P3lIHzQOt1wC7zTUUkayVUhG
D8GJUFyXaJrXp1Pz/gl+fV2WBIyZDutivVv1KSwtaHLHJARY8pKxjHoRi/gA
bqX0ElYbZeCy2OviKwyhTbRt5oll3ta6me2k2vdMBNLgZcbfIsOlgVnZgCyL
goke62G/0gmST5egLStYs9y7k5UMSGQWXmYq9YROCJw5jz7gjDwizSPadXuu
aKZSRG6yXRtX54FSVIs5t5ArEaWnvB3vSOGeeqPuk+WxrfVXb8t3lGCKoc/K
OgnJhSBLESFpQ0V4hEIDxqtQCKDQBU+DKeC3Ts51js+xRwySDBlGI5+JPygo
v/ilng7hbzrjV1Udh3QoYSv0R0nzG9pCINYfrBkpbLGBzBoJzXqZdNVyfGD0
MtOrGjv3FgRwxnI8KjuWkvDtJ8QBK2mm3TUi3kDEYFVeUJomlU2a8ermjIxZ
sjpz3pzcVuhLcR8LmxCMN90iQglmYDltv6b8C0BgBYJoH4GZfo87sBjN3TuL
cyNaOS/ws+KyqINaws4QbzhPHfkDtpDYkwC4LHyQfpINiO49gQgWXmOFGz0O
ELApitbZDRYeJgj4qQTI2rRrxsMMC7vMjwta7RF/NxIB2m/4btMWQTw6dhsX
+Zia5azw4uT3HTwY6vtktcgtKY6aAAqB+GTN1yeuk/sA+BRtjhDJPNhrfFrx
1Llq5BtjJv+hanuRuMYXcK4hsFxaOnWocZejcQ+AO54B6ROJZp3//gj5eaIU
bKxob0OpOtPWhtWmr6buMM3wtlznpvnPhi95NfrKsDrKC41VK5ciog4DLJ5g
MM5f1tYkfA4Q37l+ep5JEj6qzUO3GEA+nfRCAwcGjqdYYsTwwsZzqWTwJH2E
W6q08WuJJZ9xK7a8FNxH9S15o8lDoUx/iV8evFuuFJNaf1x/KiOoJO0JUHDF
w9dewxbrRhf+XZ1ciMoZmq1JMXxNfhF5vbWbIeSxgQ7LVX3sQxSZKQ8gUNYk
D9jRo24kDlRoNkVmLjQjqQw7DpgxCKj4qcuvtzCNFsRObiCrnNLL+3WYv9VM
DfS3rnOG0akG6RGfvUzKhHa4jbD7zq4MohrRs82MLvz8eBprBBfVXkiefBts
FrQergHpLbP4v+0iRLB0KrsLBLU06XLknMqhiHVdOJz9dGstHWOvEo+04wzL
cIX56qpJlDFY/KtW43t726TKUfW8AGs04zdO0C80RLu9oO2KKEx53gZF2aXh
vNDNW2qGeNHVzT9+HvV06RpPmhER3kQMP62Fh49VRiATeogKLvgsAXbY15Ku
SbQuvDB8TtOYrx9aWTtIyqknoG0EqzzexCS285IdUxOmRDUGcFstIkbipKxM
DaJwX6f2CkmEbKZ0dV/H5IiAbFSXLmvAUcTWNb7e5T3g8QHVjHqXG5bmEGNN
P+1n8+B4iLoO9kKWJFJjrMHpczQbBGOLAWLHNbvn0b3flDyDOyuIp1D8X8nZ
LtzplzXq/rWO+VHkmsyNmxQk8v7rthsMlpQJCR46gag89f/k7gvNgEztu74g
9MP9Q5c+M9Psl5I10CtkSIUR2jBbXOeMwqVzCMNQl6eLsB1ja1D0NJJDEhbS
Ut0OX94ftdaVZDm5lkzzjfnAksydaCazDrAWea4HdY9rwc7aBHbiGTdvo/ZC
HfTivrH3ZDRzu5J7Jp3KJAQJAPAvkz2dD0WsS6ub+NST8lQCG4KFVJVlzR0K
3GYrXOkNm+8p2xkCreztAHAdicLQkLaWFB5k6k1QqkEk5zRUcQ22JQyO90wX
dG+v9XOmQ+LLVbqW87t0fePqzoUgFlA29v+dm8zHTK65syv09y0sBZWu/RGH
th+Vni6iu7RD3F0KIb3qk3B9DC07cJ6c5ADhzOxleANFIULkQgtFfMaNFa5W
VE4BvUTWYjkoIjUPkv2LrKIylk1pP3Js/lIAyQ+BopySfVxDGAWPOuPxkBh1
7LeNV0D06F7Eov2ax2W+fb8edgzsu5QfD0BNCmUyvTtRTmT4uSd1MPJeKk+s
CoQxWOBTJZOP0E9NCrg63r97VitPsm9YMTWi1Gfyv8FljYB/IbQ6aHn+I/A0
FTMfuC2o0pXO4yfaX4KphSc6IvxG3d2e96k6MmVP3/rDYByT9EpaQOv0aSl3
1I+oqzzoC4sY2SyImM6SRRpRGHvRXFJLgQxGamXU1KoI8+JUj+tgLJ6n/I9d
k583WWGXhvo9I7suP54AjN08KfyDtfiz5mIZt61hbUrcntdtwQv5DgUISWHX
che4FjPgvp3SZPp5nYgj8/imG+kLQn60SJUtO57HWMu0dNmZ8XtLH4XtTct8
I6St5zqU/Y79QVVUazJvHvdkw5WE7wlT9PtEo7nJK+aYQBXXVI5dQ+A05bUk
+nxJKpSJW91hz3Y7KPSFOxX+/wPRmOpbu9CMmbntcu2P/Y2gugvf+VhClvjb
9EWDfRY9oalNS+9bXeeXR3pzqrndvRavZ4P6pJf9kD5sqHvfr44ShWOhHojZ
f3Yw20G/7+Ux4+wr6RR4Wtx59pcAt99P7SjLIaBHe8OPcqdTS2vakUHBmb2Z
aWdv/R/9PfBWHr1RG4/QE9QiI+1pkYq64+/gpvSDzQ4GqcC5hNyE0rUF7nvu
w1Xu4nLpbsYj1P30GSjOFsNn5xJPdkzjmpx9s4lgTw/AD8hfk5NLX5thWYgq
6YpBHrHrb9VgWXqXc1btwKPfCeEHRFmYiNjpxKC6PcTwyX2Wl9v7NYsDihny
jO6Qy80XEkKqqEi2JK70+pogENcLCjKBdEH6tYdCWbPvzlzQBqvL5uuWCV2t
REIES5qCz/HiVblmvp26UzSnnAthkUo+MPuYQh3jgAhUfs1XuevOnicwJf28
377c/pb850tQQgIxNz5X4Iyw4AmgY/MBJE6opdeRhGSX0iHlBrl1DfWUd1gI
oL0uvVAmHXm3p1iUDKJ+3NS33EOQucUyPk3Hwpy/dS1zsXdOWVdeJyPBVXRH
8fKFE/7aLhnYQwfFk8sef0lUbRWiglbhexOptSDt9wq73+gJvRS8BXJadgXS
HsCeIBogp8gMkeWkitDmil4nQ383VBhjQvNgqCK1q85iRunYhki/B5kOkrG8
hL4h34g5C4srD+kCen55yYu5jFob6tmgH21G/yfhdzo9zN02TWVWq2wxqEqa
Vv+0WJ+PvqhFJ0bmPzXtWveFg2EcOU7Ely5MHjwxSub67U27h9nUpLZXEFmN
lMumOz0ScyjlDd3gZ4QUEzMBkro6AAq3WAaWbb9nKh9lASQyLOYCKAVVngp8
csAE+TV2hlaiXtklsk0GiTGtIr2VdxJQU4l3sGUQrfPi0XXiHqLyWhvSRi+N
Tp4i8DYaMhMJ8Nzr98eQsRaNHglxIQv98Ax8nHY6AYAWVXa0nBfVTLSCKbO8
jvrKchqy5AJqM04CeePDK0363XH5d3L6196Jq2RXV6UrPM9u/f+EXMBDbCoB
8rL/EjboCiScCX9L3r66nyqwKxBrS+u86oysKvVCjfaOHAByNo5pF0amBkx/
jKS9abxFVCE8GXc5OjvjJV9F9jygpYoH7TW9GhNr50sB4M0BC9KoO5SmNtWh
YQ677V1VGaQ+/yK4dkg+IPn2ZDsJItU2OzLRQ70XQWwLhL4ePw8k/e20vr/R
9a+BfR/QK751a4a7tAGnp/b4umVJ0eCsxAHK33Ck15G/dbuTf6qi3r3uoFo0
xpqGNJNeqByfgG5Qhkx/ohFENvmWUaQ1uRT1Vjj7uIso1y9jyBhQ61omIV/Q
2mNi2eFi9Kkx01jqhZe/joUIT3HL6Kt3Za1gfup20mo3GzCzrLBscRrxkNIc
5mhRHI5hlVZ7PhsfP8bV9eLxeAedj/hH9wgyk0U/inL3e8p0VHQPMgEDLcRk
Lh1xVjfR4ld2YfyH4VA9e2VgyKtv3Kknu74C+F/9P7WOEF6eu/snWl3VmxcG
RVHKAKCEOIGBwW0OdPdnsDXeMQzvvhQMCsFBV1JMbXXuu/5bRxHVquK1Kv1U
WBN/6xOQzFsHvLAj62eKrSmWEhPjfSaqIKs0457jI1iCn2JXWaRBbgzM7xSD
ScXN4BYtpxMdeMU93+mdYtSd0RhC9zywBOt9Fqs7EKqIUr7Tr45+1IDzm9SU
RnsyTBCq5u7yHzQo2wqrvm68wKZfYgliTGyXNHAL+XrvurpsTPWvDVbvuEGg
/6oUf3Zaz+wIU2jb68L5dyhNycT8bli0mUNKQVd5fPBBA1NlbRdfcgemUvzn
ZzNtpBbkgASM4v24iRhHX3uH47dWyX0SOY7DUjBvmD8ynX8gj6C9YCTsUw0+
sSLc/4ymp03YO9AlDFL1PYVkhoFjuNrOGQE6ixmaOqSkY8jdwp4EOe3PHOOo
rZhKaeDXR6wtfDnix70ktefGL/t/l+TvWXSu/jPp+IuVhL0h4w7aIrtpS9eJ
7Qf15SPb/qudiWjHP/itDFhc3KcmZ3Sdt1nkXcPNo29cvPFP+f6MT/gUEnZ+
fpzJiSbYWzC4EnSHj5WLO7eVux1y9pELcV76dgsNAm0FwvR914sLbpEy4n5V
4VUJkp9tmbJPf6ZtOsnSX9U8B3xA7IHtlfXnixSZZseRHqUokEfwLurrxrFF
PWpE+rIhJ81TkkSqca3SGyChAr4+788Fy8s6Ydq6Hzm1osMuPJOfkVkQY66L
gRtiYuFCoKNvJHO//BKhKDNuLTMyrAm0euShjjpct5F+2Tn1iwbjlLz9TUdd
bul/5WBIVolk5h8hpXunxflbj/j57K54dmwtoKDa0XlcDi8c9qXVSvc4xK4h
+s1f/NY4tUympyIMhq3SQkGTIoP97Ohvtn05NQ6CLwajDwFvg98GTWqrM6Rw
ifN3njunfITd4p/PMhetjcHxfSxPVUyxBh8YkCyp8j7zAb4L+k5WrQhKCXCE
0Y275u85cyXgoKe5t9NFIJjvXtIcVR8sk7Rdcw/wSXznLeZ1u8Ch4Ob4mCPk
FCFdNeRMsdyvc+QEfDlbwlVZ9QfwkyaNihhjjbAAT4ramRRl+MBCCZYjYZef
J4hSH3ChbHu7oiTc3Gmd8I1v7BkYk7tLcqMm+m8v0JxFdOESxu/m3eCeLYon
LD63UwEThxUYggzh/tm2RAkK3iWExztlP1FORdBh1nEEhe5V+UXF62NMq6xM
OW1mGuSLs9LOqn4mXP6TsL/YiIZIIqK8bajrcY8d+jmDKekxvhO+qW7xeJd4
mL572/8obdrFASjsfzpZtRFZ8jzA1VelEarKu3LvN0l+YUhNYHcyFYmrqDls
+HretBWUjVe4SI204zOiOnZM+ldBENBZ9eh0huUKv7mphljArxkBiitr1GlM
aPsX5eRBwRM+/oNxXE3EpoB1uFwHcvf0MmcxqX1ST/ZB2dhHAw0apgN8wVah
sbcHn2rvJhpctUmbvmTERuy20CYms8PTGEGedtc/aGEc6YRUMJrhX6eHIPCd
mIWCulP4+HL6cfMSrfzCQfYRLaF6/Ii46ndmKosVP4Yk1iH3jhnAYOSXIYOx
ppQjVXbbNZ3WvAsNsVqDV/xNT2QcUb32xsbJXm+DeofXIzNrqaGnxxb26ZKq
Sds+vyofX3Wj+itBioJKMIReZpVAVwSjlNTfSujcmwr590snI393NThBcRcH
jw2ORckciM5uQhpaB8YfNxwWrevZdMfwjH6UyedLhgmJBhwtifRfFXMpD/hY
2kbr5LrYNVAHUb0FI8jSnxBm/19ZUbLq6Hd9RjBdFhlP0a3l1SjAmZcpmAOV
+oqj+tOfvS1jV1M07xMtksHqvK2zEYEeLwrl5X7TpQWTdsE4kFfYrbEBVRWp
ilPWQT0SGSD+rfFIbJ295Zdj9V8N4V+ULnZrs9bu3FoEIoo2xwCsmgpUgWEs
51cTwFVk33/J1iHL0lX51WEvEpE2HTrz+Ipl21zODlaIW029DzD4poRiCcVV
WxOFsndXXUzo7QvRdEkHgdbSqSHrbgwLlL3Gc8nAzuSgeD95QFkJi2WxwfZX
7SJ9tS0/0EhUMcc8N6EwCjsSiz2lC6Fh2onAoiSBXPnkyWMws32MZV0vK4UB
MudHs1YE3jVYlHRNiiEBVXM9oRFksbZpF+txSHr1m2O90IvNNWCLemUAl8iP
OiiE88Ndncr+siCjBnzCqvuTe9v10Qw+LOQ41okdN+AcCAwp74FavF5TBlzT
JhMEUfcrJAinCHowcVTq2vBv69cRytRu06ReKRJ7w3ZIPkPUR+/6kJ4W4vaT
y2N3fj+bW3pNw4t/JoqmJvMcs7EJ/NYQ275A4PG6WpcWMk1ClO9jbaQ8FA/l
Hzsc/VtNTcm2A8QI7S6a1nmUA8+3LYVdkMj6WVBiPnpmvTGXmvMa9QBIQps0
P7hih9YL0ST1tWheLtZdzBj2cSe06QpPSlQr1kysns/OpvaZRdpu3sFrkecs
MA6XbKjYuttNNp/I3qnhzuCAQdeBwwi5yQpGrnQhMItvH2iv3NAccKbB4Qqu
W0rm44N9urL4II3Q824e6A9uywOULlHRM7d26Y7AMXZdtbP88RU3bcqHewYK
tJExqJLj77KqC263FndyUc76/33KdxbYSJd0spjUECaKXm/wm1aEYjODpJG0
pPzdCtJCsIv+odDP6P6uSF2Va+/ltGpLNDTaMZnJodj4yHWriWNUW8/8+8nw
D4PQvHJKPlwMBB12jryPyxTLzpCAlBEH9zPeJCQLP5Af6fkAkocp4glXgfRp
AsdVllJqiG4W+VnY/l9Vp7/PdttANCb4kliHhXFYJDLpUu1jpqfeAduIBrWL
8PVU7BqOsKb2LwY8nM8pfzsA4dybcnZnBKxy8CoZjHEAD7w4lPj3rLzihz1u
JMPlFj0Vf4bPau9Ov9q5+9qVentTNLnPPYiEcsASlO+K+lgsmKbdSoX2YQPP
Dt2Pt4E8km33vIem3ngTKlgTiETI6DuotJkS4V7Wpvq0GcXPk6ioDyXhKH4q
3hTqx39eRMjoqdPQueIVxNJqcBbA6y5U1q1bxFyLsXz5+lPETrP85o9vVJ+R
FCmsj4UyXoGn1tP9fiW23zeHCCnMNcmBlgzUl5QrA5Pa8Ot5WOOU3x1TxShS
VwWwjXH4Y4qz9fd2BwiVZIZI/AojrX2jl3Y4AG8T6nxlSWOhv8AqnIynyxPO
PDC+0pwiHKmCY3e71isIu2BYlC3V72URvUoMiGM0hj2W1pgIGz5zuVvj8dZC
lspHYphdWEEFzImUAQZ7j40dbyMuri5i+0ZHjYazJO2spRsHm5q9ExSs2Kwq
oTRrN/68adik7SDT29EA+MDFNtN5zs5tjyC2UZZP5VqbUM5OiaynuHTyFPzK
TMA2VmyeWwrJ/Azw4YB80e55yXjAiXkm019YKcAoa/urNAIJ3GKENPh89q2D
WOZkGBkPaPXGmTPXAuPMSz22Sg3wj9pD59M6uFHyXjnCl+aLaYp9RF6Or6RF
R1acH5VzdFcyfvzeCDWxQUqi2/Bf+QgqW7YJRuTtOnkesT6G0MM/PG84k0rp
k9Q7cI2kr8BItDyvJtrOx1oBKz8aySu47AJ8UI8SUyUzF1Ou/mEnV+ghYIvP
Np/c868IiW75H7rU6sjU6J4TNyydl1hQhLFSFKNC5qH5r0eHi+PvNah1SmhE
5j1GB6DJ/3FvrLt1f23tx5UFNqkvsH3Gi+DYKnLI4gFYArMc7c12Y83k/mwr
/5qaRIFF6GRBj9xi/07RRv3XYQ07yd9Py6Fga0q2zGwEarP1QwZwGOTIot2L
QCme7KetPfDisKCVU+FP6MHInhuMCyAJ2qAwiUCk+ChPtrT4j+4Y+VRJzAYb
v01xs/yQ+Xkkzvo+rbTU/XU63bqtR6b+mQU1Ce5eCAXwBY+gqFSU3hb+2KQb
sCkW+m/XVZBkH8W9Gx2xcVsc3DE6KtXX6V/6sVEoTj3DfDdOcQlD/8Bge4tm
pOwRN/X4fac5iIFgmPO/o6fTFFW+tKFsO6L0IpE1yWbaW/b+ZrU8/5O9deXP
PrfnkXF611hUMraS30YleWD8X2lrCWMkG5ah8Iy4CEL+5wfLZKsvl1WdLe9k
QHvkzetViuatifuzOv7VLN2o1hqoBs00s/7JJy40ZGSs+hXnZAqw33Wv5yBG
XY/f9yCWhM41us+WvC3RAXlEA6lap1Dk4DY++s/aPsPwz4kJgg5lkEyiKQCQ
bx/kdA4Q3n4Px7SRgKC1fUMRCIuEbX7aLb6Jg5KrfiKYtqPOGFoFsXxUQBUJ
p0ZNmveKEc2taHHi41B9Ki+YorhjRQHE8HOQl8FjNJFyYabuoe3QS+Uj3IA7
+PPZGPU9zr4S8S5UXnnplXJvvAnoZLMcg1baE09GznvZLk4Yss7iq7ChGNQ7
iHtnNTSnuC0ykaGzHmqXoBcVVxZFLPuvExZiIft+/9PBDlGzLijHfSIqkq7p
iwpaYF9B9kOq9RnYGFvNsCvOBacM+YIBCPUL3vhC9BheZFHK8m5iDB+TuhlU
TCmd8UXG5H2qGi1l119VGP/jsrFZlkJE+UANzKVRq0/LR0RCnxjnn053F3jS
Q1VV9HKLea3nFhK7yN6ofqBvtPcpl5YhotbkUD7xBRTDwh5PCZwYanSwnMbk
gsHFNJebjASkSW4aGtz0EIulbv+TDJQX0NY+3eK6Ar2G1Ljepuqop1cQuhI3
Je5gWKua7oUj/vCDFADQmDsJV681UGlrQkngAC2WtSncZy1566y/ACWoKne9
Orwaa4UgEwR9fHZLD+7XxxET7SaZHUUqgMVhXpsMsV9eys9207jTp/kdCLE/
nyk2eDUNVMp8IodZ5MEsi9dABAoPk829mZLrYvqr53Q9hjX92n5w9QAx6Byi
Mk0vg7FJGacuUObQ+dXE5QELLVAo6OOiIUWzlejAj7ATkPYT1HV2g7HWF+2v
m+4t1gRlDJzflWA2ztTtBIrf/jlTUk9eYFQuOWI5knEAzIWM64OJcBkS0W0o
PL6eV54Jhnl8ww83lOMr0cwZUMSsedvoJpPoTxEIZnHlzxdYfu2EnUMEQ+J/
bzEfG4VyUfyWoQtbl3vbz+kxqEAuQiOAT+yXaxerUAKKJ740PfErM4aIZblk
aJPkjC4eXCd7zcn6Mc7VsxTso8dozZ0Ijcd/4VRODe+6JM6HdpwE6fKTDbI3
6fNw26hiWvfjyjgGOhe12QP63cRa5t8xfykbi3dB92yGs+LfSHFLLkhO/BxC
/mWRyRotcPhLt9cVesuSWtk2sjLcWDXW9oCo3jEclgi5qqnjxaDCNmLlkyl+
Q9VQCeT7WJLSNFu6KUj0yu3+0QbWf3kZec0muQrbspk9In22G9cwvEYKeyeF
RJ4/WDDk29Imh9UMbDVyuM2VP2CXAOvZEh/NRnnNUw7aFDmjtySyH2yZSC+y
r1EN5smVRh6/xS+84MTcWldeBrCgEPgZgMHd2yF0lPgpro3POJ54C9UhheR1
cy7h4bdf3FiiQHSPC9K8LywXx0OJ5uCTqrbywkCGI27hYrIok3EjHGdTVjWC
edOfY5C+mW65Jg95CvW5YVYX7Pz3dDysV2CRiJSkRnjVqPQmldfeoixGZ4fE
LTPKhaBbDCG7RgYH9zCQlvXdfH6hBupIm9M/SBvLcC5YPULzDx4EVgM475uy
0F6fYB4m1RISVxzCbA3OXMC6SlHt/pP3KhQV9V5MQ/COY2skhSYwER9hlKr9
ljIcLdk4hSd+XZbYDAxueqML3iEDkbot976nVsTH1jV3TjUfKKkCRrvAUmT9
lhg4Oqonr2MzG/39wE7xkNB6mzedLuyCjc0dR91T/059zMva3udaqMOAvvqg
fmaHeRJYqUNO57N1cgALeYuzRKQ1J8ebcUnYCxAz6+Mku7jrn7Q7jFRcjA8G
0g4GLKyNxMD/FNtVWnBPoRgh+YqxIrRCh0+p4zL2/8myAbh14Z6neAjQcBiW
t98Y2RYdiCNi2rIhxixwdF9lZfcnP5AVwcFr/N8Pw+FUrQu65Ks8/92E1Zbh
DDXXyo3m4FPJ1AE8tM56Le5y2l6EV7kh+kbF1ZDfGUolqgV0IB/2uq69vbyl
EcWxt01zV3p116r1r73dm59Fski+JDqu0ftDLtkVfsJ+oE7A6ula0leMq3Lk
Pldva2Dx7fO7RXQMHyKtbgtsM3VWOwBedKpKPd5HMmYDf7xIlIvqKImS8yJi
och9Ej9IbVbl4n3bGhtChnhUVMyl8qKNx6/1Dl3+TH/V5HJ4UimMm2w9B9J3
0Vw3S0z9cv9Sll79lnjO2FMrzzp/Q5Mdbh8jJHbnAhCQDvQ8mBz7wFQqiPnr
gEe5fn3Ssy9INMpXME9Doh2c24PR9Iryq14vaLCRP6zrsoSxTyZdUDsrZNk5
8UWOfW/UDQQ8EPZc+wBp4shukBIX04SKhVVPIu9yZMiG6x2t//DLE0vbBbOq
K33Y2TZWt+Bm+2vZUmb4mA6tDn9CSOUR0eqAxgyZOX/n1yuODgxjMUpNeaE4
uOC1OKShMdBPtJvgeBRcZLkPwmTuEOaFd5UJwpcsJtJ/CQwIMg/xitxrOBm0
PAFxVJb2VkVn5VJlBCdFortQV5Liu+lJ8el1JNyzZa8N0x2FWCIq1thtkV+8
e51+V6JStXyNMPOHWXZykYdM1WT7myqLi5e5SKNDbmX17dDtJs8AFPR06C1f
OP5srQwg2ipMr4S/WrjFSQXgysI6t36l/7/keUYnd/VCCoPwZh5/nQeLwbO5
y91ykYdrLqSttbm+ui3p28bm4oDeYbr3E92SRSx1w7J77ZKvsV+nxCLHfMXn
9n/lEh7MRa4NvR/p0UA7HWWlHz1Bkd5xqstvKDGU1SkH0OOqBhcwb+7YKbGW
RVGobNuKGK+QA5hXPfHvTC5zLWtYxAB29Sy/NqDYS1F947xNvta2N3QZPQ2V
+oC8eTVoHCDG5TOAY+4joTRHpO2lBz/NoH7SGUM1TN+oWrNyHyiuzfTy0kjz
kvxLnPJOvv8oWqDCC5JzIumoMBpv0tbvVEm6llrGSoYj8uhA2l0cskdVijGn
LcMBCGOpJZivVDVVt0romEmKwnH/46CA3BQIRioKfMJ6jGCZpzuRGEbcZ4Cq
oKsLhUo7AajszEa/JtaSMX5ihoYXu5IPZGKMYQqyqA5oLE+kplCxyGGaV0bx
8jIAtp5jd2iIoGphs/EJmY17uEKkQ6kE0F7guz+xf4fk3vZavDNj8bKiTFK4
DrvkUhQi01riOSmlkf52uM74mTEWdTTDgf+byfzXLpRc6tw6hsYV2/L/a+Cg
iX4iQ4Ezn+96BxRQ8cEWepc/LQsdVjgGscP/BOGmVP3FSsgwh2jufdijw/BQ
yz6NFiaIq62iYX39InglNpkTy2/wWxL1dJppGcwhetU1A3farLE4bXCtQVOv
tGTDUyMG3TDfjpiLjaB6qarXy2inpv5Ku/O63s18Rfc0QttmurbttJN7QSuy
B2yqMbE2bn47/YmZ8EXPQ8o8wcSTNsZLA48JZhzzdUdfyzZFEHpc0s7c8s+5
Ksw1PKGxYO/ywGTYFEyaqXre0r/jntbSGnfrSZNg4g1QEy3GusGIEBM2O4JW
F59+PtK8t9HJm3h0EcLt2BIFPigC6fznzrub6m/o7IR91GTnx+XP22WNwIQR
Z+AuU85Tt/aRHXO75ae0PQL5qbf0E0FE7L3ZsSfARd5QGc+kLix9Pr2bnrfb
hkqJ/hJBzfzmypmuYpjHVACYucq39PwijCJRfCrNmWDOCRdU9wrAojRksDbU
06SUT8U5+07JhGZGK/PNSj1qNbKM8M2dDA7fHnDOFk1SH9KfcRNFLxaqGmV7
8MvZcxHifo7qbaGmP5CWvR3qn56zwx+SIVTPOVZN1bHs/Qxdj1FPitiu1OdW
3EakUJgr5ZKGGHF+KT7joW8ICY0V/u9ybbv6kmtJ9fYOTW/D7sd4IVB+C8xa
7AxjEhLBUFnoLbex7sZEIKrp/AQiaCeq9YuzMe0LVXR8FkNdeweYg+I1Fa39
E4eutmNJGCZ7OMnUs4CrjU6DdFUjiSa0WEphQVaPK+mJ/wmUI0dSz3qRmmdc
AXpxhUh2DZXOnBJ/j/H3qJUxghuqD3a3M3y7te3VomNoabesONbL/LNX+xag
z/Cn0cw+pqQkONeWkNq4QWMRcY5PWIkLzkkWmwmitH5YekMqitFaejCZN9Z6
RSLpIkEQG27VrpsO/x5QDA9qkrV4ZD7YYfHu99ZPISVAv/ikk8v1k7cw2h3Y
MVmisq3H16r7cQ7djwPJ0K2K4IeRNmrBOvvKVJ0qF1ZwIlOcdxjWmbw2dbZ3
DRGSgHOmma03wtJJITxQr22voszMAicv96uvEOUr3S4sTh6qKtKfjNdJ3J65
wxB8F43BVeF45HNuzIBcvmat9K7JZmyF26Y9lAnkCFaQxTdnfyf62x9WE6UQ
CIg0bH0Ri2y7PPQKXd2IU3kibfl0r53JX7cqQnuY3VImKMDboym5kX6lhvf3
3KwaXGhQ8PyV84Ah5raXweo2TPum+vQ4xzx3xCn/oIoLdPqTjS5+nMH+dgJt
CpuDbunN7hPAgY8i4+E4RLKiTtTu7eiy0nBDYZK8W76SliecK7fesBGLmMav
w0obftH1h7M8ndaUi/TEgGtDba0gECiIjPfY+jxDUJyEjESvcgi3MCFuI56i
9zBMsjQJ3kq3LhNPMK2ClAiuvzTAIRlqsmrN9nBDBWPvJYJorxYeKcf5zgDE
J4/u2FuYnC7dECGxpKjpJ/A9WJ2MxcR7GqunLrKWaUwMt8sonQa65HXiibk8
UV5kug9JuAZGKW6feXrrCk3+tjZDROrMuIVlTSLGJWc+sCKDhRTiT+Nawruy
FY1CROZ3MHTsitjq6Jg68KDR3d0oEs9Eh0LVmlek3vnv89Posul+ziZ+mVkD
PStwKW/Z2cAiv1Bp9YfwgYcbDsWiHIQvqM9YE5PYT2tEFYxv1QrsmdGw/Dgp
s4u+8Y5DWg+is5tM9bLtwOznec78zKrj1MVFbKBtwLyJ/qQwcME4BsX0Jbzx
/hV+mtKFFzzX8LlQx7dgc0jDbgxumbTUQMR7AN3O/+dOEdT4BNx9LKvp6iN0
uRiFFkTuZsVdRKvf/shmqNJXTI1h3D/MAvPXXYkUpNIrHAPtRVHqGnEO44PT
9GfqYpqHfu5Z+jVRrSJVks3fwYteDDf5krNHU1uFCKZCYjOF9iGVdNSc4ED3
qWb9VWU3V0fTW8XovN6LmiDCkSOjrgUohB0Tulqm+o1WXipu2n5KzaO2HvTi
cumrmq9jzZ2EuMv1T7KxYKaUkVpi8VSLxkeBdrlZcWy1acmh9ipvbn8IZtxW
Klzzr7XVN0Q9crAOo48M9lDFHgiWRnczDwBuf2nzE6y+Kic1Lf4JiXexESHo
RJRnIyOdOTq99Z03BES8ErxJGaa2eYQais8ugyMPHSVrh+wjalEjy01Y9Vh3
GrKZOEEwJWDVdd1sNe+OREWPWnryCWIoeROJ/KgUo5c+AzpmclL3qTmHrsap
UkxArxiQr20Z5QkHyWfCuirOYrDGm42U4uFKH8BfM74pwS4ALwuvgoylc/7B
YY4iP1VpiVgiw/fm+nN44wvKuGIFUlQWUvv60sF/1dlgrH8fjubLcRCOWkr2
bdf/O/ae69YWnQtG9Jun9EEshI6TTTk1jQqGpRuevPXifJIUgMssN/Mu3mxB
Pkv+9sokAhjbyMUD50qVOzw7fu+v3ijSKGh99M7LQoz8AVE/ByvKjizQ7NLB
ENHeIYEnWZTyN5YMUMmq6Tib8FEJ90S59ysg+YxlLPxpxVtwhKBb28Ycduca
BYn+VE9HtpPyPL/Wgfl1kZdiQDaVFLrmW4biGimQNhlYtFsDJtoCtGpy7XOV
2Mgx15Yx6mG315UofXG0ROoIPvDyqfi3IcjM5pCpON6MmtjGkkxA9Dpk6Q6C
v7MRXu+15MjvyVdqzjCrzdhvcI7oOK743MWZ3L4wwKHXe+fzypwHDNnGPUpX
Qk54RtC0ty10eeDZBrR3en/t+PzRJqZHDTM3IhxWy7hefOStjwYJkkWGlcyZ
obN/LLBk48XQq3CDIB/VU6LRfQjaTaKpoullQmRltpSr+im4QMT5RxGuttvM
gJoRHep540U5fRW8Kr9WS7chKlLuw/iRWpzNuIeRXqNEjSSAWQRWDQkvP1ID
0RcJ0Vh4zFnx0b3+RpLIOmMQu5Eb4TSVUY//T+uMtunwYWRF70xFnaGmb5y1
pCVdHEvuW2V+4pciicv49FYpYUpEy8lYlyAHO1AB+hKKCO0lrkquxAhTwJXL
mooituT7xx1TPpsKRL4hWZhAqShqSKVw5YFpi+2LB8HhGl0jELJpAO6gcUBF
WYoEw0FPdYZF1V1cEkzB2TwpJjryuUcvGO1vt9643cY+WeEuNplArM/1Matp
CFHrLRI9We4R4jG2yIhk2pQJgttxYDweh3e4EJ1T42fvZJyqvo9NdzG02FCT
J6Ox6Qz/gr28iXbSpAlyFq/DcbMiuExxcWZG7qYpbfsLrZuVb9jcFg+ekysN
JuNXti48gZPpxnvuqTErMPuiIh7xuI2mk8x+zqb75M+W/eLvzXYwdKYunWqp
VouSzE+vr3XMB1aOtDu2QcCW+lBka0KvIM9240QSrzNdz72Jspw+z80fHA7k
FPOo+K5lfObChuoPCHgB3iVOcUxPi1rbgERlZmqT+phW9Dbzxea4bzcRn7Nq
kVRWDMFDrrT5OQRru8EuDjOHjvFowa2VfS4EGeqXvMNAqNIO7oyGv88Xu40r
tZdMU4bAU82wcvyFy/r8XwtQ484xlsThzqRERz2hcraIFE42+8z+FeCTPYIJ
AYyeTmqiYOGe5BfpNJWJDsEp9CTe9nqdzLsXt89G3w89BHQCWEc6t6XrPpzB
RDxVTSsFcLBsE9IvM60vojBUNTFK6+Akps/R4pEhQUBHma9TqIQYPgcL8G9i
yebcXAVKtjqkLgw24ZUQiHKuPxRiPqhmL1dH2Umh7n71oVmhrgpi/7hzAwAD
vJjoBqeLC69nr9vfl4ppxfp8NxUq/ntN0On8w//B4MCDcZbPPT7j5uVOd4UX
TmdLG8W8WbXWSNRHFToFNjKIU45/VitePikoyWRjOgw68lZYZ+dL3zLfCoR0
qCh6KXtWntaOlXETg/SCd/SmGW/uFn8la0YMZd7PXHAjpdXYisXL9TWAk5vp
EKns7bVQzez3zOC8f6wgql6gzx2shoPdcQUzf2pUJvaHCnaMKa6pXkP6+hFv
r2OOIGFbaFNJJT6DCj3C5iePnY4L73exfOPKfenNC6cDeHOya3ogOxUU00Y/
tZFofyvmLg+OMdFfTUT6psE6TJgOFNPGVL+YSLnBYkJbX6M0+QcehdlPd0uP
R6H5UuLT9CTovDvaimHrvsORz0DQZOB+lWapmzkCFpt3TBNhadURf4qDTpEY
puyjwzDQUwkJO67BfPRQS5CnM2p8xWYT6ZuOIjDGLUPLYx4b4dW2d8LLho9k
P8a9TjI9p6GLSDqIHMa74CmR1wsWy+YopDZvtY+Qe3kDaOKdAsy2hHZPZdQj
sGz+U7tRqkkAcqKc3+QgGX527QGD7vT6B4lX9v3oDaHyEaFS3Ubadupm0K81
JGRwqa81SrOkU3mtPUBAwzibC0DuQYFGD+nY3b5xXK/hvtzj/OcKB1iAAE/w
l3KYI3P1Z3XYY6UpUdY2KPcaeqcOYKGbpHagOiPk7eV0Fu2U3BIjgS05t5iL
lH451Xbbu4eaYoo+4AFHVA6ge2WCHhGog/b1Y9sOC/MaCNELJCyfbKtILohn
sFbuRhbY80RSIkQfgcOeO6KDbGf+u1ERkH6mR5OLb5av9FVAJPPL5wHHaEhU
jyWLGYB9Eyj1n5UqMl/LfXNlmyBGUECVGKtCl8s7KGw5eHBcdOXX46jO0U6X
tpBHiMlMX0DfP397w/Kg+5kpQebfR4HgVProcfFUtosdOGz0YGAQdnvZP7a6
OWOQM/SZI7I2/AZFybXlfrMxt9kVlKhJi+B4XT6zjFi4iKxIDyaz+6Ldl/0v
YglPRU1x3A/LGREf8lAP7sw2Oh8Mupzo/iTUX8kmUKB3jGT7eQUk0PP8oml5
JpihSeqKLcdqTtSi5lk8xJbceUkkGBucuR1j0LTxQmxAgYLHKHDL2Sk37kEX
YfCX91dNk2qVx6/YLaL7QW83SLCqrDEUyeIFQp0xX5pMa1QcmJ/yvuNDtWly
KKtcw1A1WKP+TcVlyx6nI+4GMDirKShUl972Rz4dqADlN22nIWIbtFbUlDTX
8nuNMD0VG0Ns7hQDTskWgZQDcn1xB553nXAYSC+9TTjZ2MoaXFh167v6XB9i
gZzJGRXuTM14vEkIExqdWVTBW1/pY1woN8aKPFbU5q9VBWo+wIc6mPhuaqVJ
lrRWdgaEybiwxBtOdbLLumEwsCVA86C16BmPEjgrgtpO82NrMev0hlGetJvJ
jspkU6hLNJztcD95J6NyKUVJtjM1lcxSnq5YP6iNXROAlY8Ini9/JhwzM/vg
aiJvno9bunU+X1u2rtiVl4sHxNJklJ4BLsK8FrSEjvk/kZR1ryv5qKWDGUsP
OawDafLvaXp6RBt17yd3hbQ/qICZ2csKINoNmNrZfhOcvE0m9gp4//Aaa7e6
GcWDueo/INFgUFp46+NvXD9MNjJzvaHyV2y7YLiSDBi2Mu480epUDJiPy7Y8
pXAbtdTMtzha7qpcSqC5GJdoah4IXLpmWrMWcCDkpIAOPI8z4My13u1F//Xg
7tnHL+Lo7qYyZzf+1uwzBsh+M8mjR7zK0ZpkZdYImHUXIlZgI8hH+/eI78Ey
ZxY9RjSTfwMHmfSlAaff4OkyD07pipyglC85a99zHl/f22DyuG29rIjB/tqr
8tpuRIvN64JPkK5jO5DDXNFpA6FJGU6gQPUx/Mw2pbrfKgfKKEAhvnVihhc7
aBzUteDD6VKxkaPZse2lJHPfjJ4mkBN3d09HuwjD6f0ia+SRkZTIgROOwLyg
nZ7ZaepnIPQBR/q6KL3mUf+HxhIwOOOZCruM+h9NmpPYTJbQTfZRIntP1wch
NxEdbaZ0lEoYX7DKZz0wkuxp8xYfLSvlOdCMqc3/xBQaNeRHjfRnICMfH6Fn
Jzjj7OF+2j+mgMeV1vZL4D/drC8BQG4X7H2xeBWr6s0wH9xJGUHPzzqJWmS4
8h2DyD9q0Ou+YkNUYfJkNlJhrMM/GQc7WwQDKUXCxStzITpiUOprHlKC+UwT
DDz9x6p5KBaV7JvT09hfzmwYz834Ye77Aclqqs1dOazfx+SMcqwapjPIYCRt
K2Kmxy3Lhy9+KOxOTeT396UL/SJXllodC53UmibwphUmz5c7IotcPWmlcIqh
w7bkbcLagy4yWDVbXM5pLa0uSR+dkEej8kIQMfhwjH49pB1Hz8TitER/VMVA
5LrmK5F4+L0uoiCGp2Xl801wx1WTLGcF5vXAhmTkeRmSuaNWqfbjTFXyZ514
FXipg3OFEtCxF4eOJMG+4QNNlC7kNKB18u3lJSx72/3rg++A6SFRt5xD6jgc
ZVV8JnIV+ZGVl5JA8r+Bf7WPZihaqc3bXQ1aNL+Z7oF0CJM34Xc11hE6mAcA
vadOuAtA9MTExUqqrxbKO4PCk23D59eXXdcEV1JqSTV88YYRywDO/Oh1jSKz
z1d/30XrTd+JfEgPuTJpno9f+MCs3mnA8mXh/Qby4ozOAjdmMa2affz5yOqQ
Gx2Oym9yU37Am8fgD0boEgC8AGdPYJIqhBFeXqnOYoRdgrp9c3pEySsRvlYZ
c619q6/XgtdRuahZHAsOcviLBD7UczqkIMTX2/LcBZhXOk4UeUU3ChvA5AwZ
NtM6K5LqdHVI3jnTnnm+5xIlS14P/xmxdv4PHEqrukYbv+7s9OEc8dKTe6Qx
NxlHLgbTVt+y4Qz4xs+X/GSvrSGhos5kZt9ygSsJb0sR0JAhWjTUd3puxMUW
aO2Bynspccf5pazKJX3Zqs0NMaOMlvK6p2qR/Ccr6WlRvajfpiKblIOvharO
McQHrSMa49rJ7K7gL+seKQ0c/b2754rvOeY6CZjruCjyjRQdMJfsjIcoZAxl
WTKg0QFmxU6i4rTMFxueoofgkOVOueGAiDPBPDCiwADvlhOIgdHgx29SHZNz
9wz5bnOINxVyeY+8y3Sy/lpYFjz9W3s2eELojU+skZ5uhBaZYyM3l+Qjjhi0
dt65pVoBj3lIDEJRoe58n0yRF1M8LRcgYZUnoZ6OoCqIWHfklJ+Jsj99UhYm
tJiqM+WRfMLz7TblkmOSRGRZqFUU+7H82Bf/LGB7e4G7ERm3QFP/WKoBaFor
4H1wVKrwqL+9m2yaZ3b6fkHc/Db4lDmXMBed4GfISOeUhO+xObbJDJMTc71J
52c9plkuLLwKgK53DPp8hQe0N7c9O2DLmOAGS2PEXwlXble/Cf+XZVH8WkmS
QJUMC3Qr5RxEsIWYbctfNa4Gve1N7ToXJy7qxRiL1HqNkNC9nJozUKwVFxJa
35GQ/exRkxGMi+Si6jMUK/Kqe5WMQO8J6tLFeD6U62K0HAedM0arhnA7sbet
CF5ZIpT6y7Z81i+eAKjy6tCkKcMrlwpDjRK5iKwMXzQIpndMtvn3ySGBj9rY
h3nUvYDejDAw3Z5cd86hR8J6Ke+QpcMW6wafWS6ggTYlejX4jQJAgHc3DUvV
hU+MmVSUdGWSwJ/GwOIeTzktTBSLXd7e+AC+qNGCO52Jc24hAZkEAy64Af1O
CYtP2w83bvDzZ94s2BX68RVrY68W9w2Pa4pmSVKISntkj103ngrb2UV7B5tq
BB9INSCWbdFYXFKcWwvQxLL9BEHsqJp+7XCr0QnOArc6pysC+IBxokMabck/
ik5xANeVE5ggx7oUntKAT36FPQxdqcWfsOF5N4RZusBOX3pNJLrtWsmAxUvq
YadCnLVVtA5vIA5pyW+4aJ5o9WIMXrSyrF2w/Qx+oyKb7+iboJ6mR+4YG7Af
TKWcPC64agrjNqm4OpIUbyzoVZl1iDdWG/XKt5B0xwMTkk4Q/ER8K0T8OHWD
4zMRfB6FFOE5kfH2HZZGaZ1e7zOF31E2FszSYV0TXdEt6GJNGft2X5K5G4fo
sD/HREJCNiOfj4a2SA7586+h1fcV9FpynetloTxlLOl7pOXzQem421VyO9jN
EfpuD6Hwa++UVYu588ZMYst+EqXvEVtXj7OwwY6G53BGHWWKjHHqos9x3piM
Fna9sA19aSHToNQnWxJjtUStQkZXOW4m6lJMLuba7nuD2lTMoZmB06NoRg9A
Dcb7iPIWBu6Gqx6TOfJnWiI/UIju6voNJ+yD+dLifv5l9izhb7VR3Bs6gC1d
YAO/woQ2I93rVp3iI3xu1loC7ILFK22h24jNfLerCAPPei3Drp6z93RFzoz9
coZZO0oAnemC2nggQI8sKFpwKwGJXxdbVwTDj6+e+PwAOBEv3Qgyasn7g1lL
FdFsjjXycvV1PFWWupgiiBrT0RdBYqgNbRPuV9Cxd316c9eEwpLuG7Q4bUnQ
Xd7bd3/IMCNKCqXixbbOY6krxqdepP2HG8IwmXR1NjroPAzCfWDpaiFg5u8r
vA9JQrbktaYeIEF3huGtafk2M/JRBa3MrYFYsp4cpPbfLF8/cJ5DxG0NlN32
PZav0HGh3RFfjfAWDnnOkKuIF+xYIVNZ4nc81jQ9wEOZmoPjXfqpq2Hl6Hh0
fleFSFqKzw46TYSEE1TVUq0ZNtnwyhQ/ONDG9X0yaRWgB2E9/4Vm+WcmnpxA
Cq/2q1bVRsqtU87GlaT+QCHJ9J8s+vzIKOo9gpNcVW7SFomaD2/b1XB/Xh6h
OyeSgyaBZebck824m4NoQ4CB5e80dc6cDhBGAZr5NTsdNG208PBN7GZH+Kri
AeBbrGqMY4Noz+F08f60SJO+F7lbEAovUIChkuVyJF49gQ6y58SHZaug0Vss
goRvhgXQyvnDwfXXz061MEQt/r8cPzNDMGf7hW1nTil8dM8bGD/VbEvd43VR
z6FmGayn+qxCTnScs+Hf7lcQhCS7glHCyCJYwCYwDc3RMd4sAA0M12ovSBak
C+D6GCoJinfWn+p+vnEZNlVk0qgAHPnxm7ht/fPOG0iMzGc8QGll+I3rPmv0
fB+F5HewknZHX+1P6bDLAXaUlg3LzzgcBKMLK+mIXPagw492OYWeYjO5k6Fc
qnXWU8RgtiFgDs+VkBKy19Z2O8w17VTg1wFx/Px8uIyCnaxT5wwlO0u5CFYZ
QaN+a44G+RvPtWzMQMrt0pAA1h90WXPOO7cmt4cpj6ki5cOGeA3Q8vkQPdss
FcCpXXMfqFkC6W8Hmns9PUUGYYrkI3JH/nC2//n776iSCyUHssBgeAdov61B
B10wDxW7Kif11Co7GT4GBuzuYtzYu4R1J7e5XFJHEihcqMGM7p8+b7Yx1OcT
HjjTuo8EZhK33tS1/di+NOINMLfS2+mxN2XTznfL/w/6zAUThoSXwWg52CJh
BoaT0M6yG8FfKN/xZFUzaI6VnVq/DcsdNc5Kok3U57ZzHMp+OGiEkCxkD2BP
9G45BBx7cjrmajnYxJKZy3awlRm2KzejxBjPW8e/rnQPWkH3ullslhxWKr5l
Gv4GZco0sqNZ2qijj+MtqbVsL+BoyeFaVYxJ+scMysrZ9emxxhmkUrt+iWDf
R5DZ+CgtkSDtoSMM1hKVX9Cq4e0TaED1zqqIAlfbWB2/WFZ3bTJQgHu5q9Mw
vUfKpx0x463BABFgm++yZxBja6oEIRGlwsDKPdWIs52PkPL1igkjGJDnzIpy
8BR9MCLIEKNzmJfb/qced1/9dVVpQqUyLhvPHZBno3O5h2J1j66MMn7WBWcE
a6pLYD/3t9UUgk7IGb0jeJNZd+rjFojz4BWcnOxdwZFQ/08YruCS2gNG5Y+8
wrRlYhUGUlb+RVuZT4+d5Ygo3HW8oqqwdozbfPItcspp4pTyZECq+ddkX4Yk
6gI/KyWSxuQXvBS1zA5MeFyGQdcPbDRVu7+kjfljE3P+SEg1ff/JX+WYTmFD
BEIBKtYb/MhOcQfnXlF3JrNYAO7M3HymRxItMB6ksQfxJO7NFwlA2OdnFxPX
Vc2tdeItwV0OmKUKw6KeT5rwZD+w9p2jKspu5tNXhmwmlfT+BUEh7WULplYD
Wz5/D7ZTVjZ8xm8U3sfOpgyurIhkbPJRJ3dsswc4WNQDLnqZgcihXqGTgCvM
DCZEVWG8Jgq616QQFVt84wWR3vfAcTntsSu7b3YQgUe/x68JkTi8lGNdRLIS
t0KHJ+f1Vav/Xocv2QCipZ2bHLZYSfZdkAwVWNu5vwBCDCPnsqTGQt7/oUFa
iytyThk4gcCoMRjPeOetc+uV3fsJsYA8nP8B/nEWnTvZaKSA2qZjDyr8u/SO
yhXHV8KhMNREN8pHifhzy+vwUVRXLg0yannQTcUS9ymmx9KVY/0zUIL7kdVy
A34WiBFLXuFNjBnbXuAQPvOYULoJYnZh7Fkd8mHABjduZ7Gjt9frCatMewDo
H9rZNzszfw+8QiOfrQeJQtx2V7xIPL6jhNALfeiXRs7vl0tsrV2OGZBVcZ/a
E6mmcyVaSfFVEUNGWC/ksU896N0u3OiYfFidDYjvQ7DLz7DudtmjfQTHJ9t2
lInYi5vP1E7cnNUg/NGe3f3ZWTl+tfLjSDpm2aleglWSFrMsOVjeJFN12aGq
7580JiKgGNJJzMtv1b/VIyNyRMaHPg0OCTpcqjPs897EJ8OiL9t1F3K3HERo
PCJQO4EnoRlAwkV+fiEd4T4jmkBZNCpB2UJwINt8CT4uC5flHbGiwg6OKXjO
S63NrZsZFKzJ0CeOuKT5fGuUa+TJrWK38YQqb74rJ99p/QhuxNgLdsOdICI4
2rwhE51iKE5lHOabPOZBQ9E2Vkna3CfdWc5pQtdAaksJNYuCEF8d0wJIVrpx
V3+LVTUwZJyBJusf54gRRQljjZcJPIvrzXoErLagQp+3/6zAQejEsbPW6/hL
vAFskYS4x83BwNGdIufGeNZnMo7nr7XsESxTwyUUjQhTvKrz6fTgCLZPaNHU
rHsH3sv6yYKUSd5jqy4i2VBZaqlhYjro4p63+ins221dprH/lwT9RJZbvmm4
PDof/Old6rOKMlaiEHmIL7bRgrZ3duf0yckWGrmIP2DQhg6YrvPM51M++blO
Cd2JOpteyIJ72aOo+VZgh2qceaD0ijueHIkOab0kEdAkrgV63IiFbSMicoAQ
e6NRdoV39Gk8zLrkvz15JIwOCY3fTvnLYQVESOi7pqa3ZbfP3SgIT6Vrhcnp
2WIFSA+ugM009gu+KlL+FhOFDP/JXS7O+rAm+gWJPvqSOlln8iJ106N8W0oS
psEJ40KC+qhh4bqaG4ID3sUVFngHJp1OxxiVmD06lRLrJ+YgCMOahscER26O
SJljUIt8DFLi3/GgzxlKB0agkc5tONOMEb4zgC0ohRPyCFt/4ZlVBRSNLIDq
7dnxEuVwHq+ha9/hcEpFH8ietMN0BxK2JTUubsmAJb6fubLuFVaU7MuMcLOV
I0ReWt50HX00df4sbrk5+tsiA7DLlAF6ZmTVlIL2xbaeMxDwSyPj1zVJ51CS
o+dMa5xtEnAPzXcaQY7i1hOVMVLkvIArsDI/ebaSS/sdS85ELVYig1YZyZoB
od0uh5hG7sqY5kLgWhLSgM5O5fnrfUPcz1IUqOjkmsCOztBRafQROSsqH9FN
wxNx1C8uYTALBl6hdowtvrAD7lyu3OT8FMFluQtUFKb+QLMKR9qYh5lmapHQ
8HuSTRyQNj32Ur2El5LL8NpO8cnMf7vtEP4uOz7y4Ydc9u+XXMcOR9MEkFBu
R/7DLBkBV6IAJnSJgjw+BTeZjHixH7/DkuQPhcAf0n7olqWACpEWnnUtLqzr
zteL1OH3XhyysGtccXMK8tZX+f8i6tHDCxgXfKx/nh38Z3BsCB7y3UZX1TPt
CQpEwOH/0srsAZzdO/EGtnTPLy7812ZxBNmQQOuXppqpXfQPXE9knOQiORLz
tYBGRqlHI01kCbXnI7+WSl2siVZEHHw2HHRHgKYWJcaX5Fs2h8KD1wgi8vLr
b0wh8ARlHjJUgyVpl5nBhr3Ie7IGPSYspUYdlE1tsNZe/SQIsjwEE7WMls5C
2AO7T6hYw865P3aHNtOwyaeu98O7aEebY5M4IPM+/g4mwLoAHLrBcakAyjUw
TrldshXT6hpXkTYO6+Vz1avtPz5zkI3dTP8+EttjHJOifSgnG6pbGrt6og3e
DIdood8Hjyvaz3zrEFmj9EWiO4MIPRatSo9NFUcCr4NJTzcNJsxSc0ghqyMs
cqnGxAcUZZ8DUV0S2enxEoedkNIhAuZevovaKboZNruQZz5RdBVazyZLMVMh
QKyp/o+M5R2aAhISyCcKSHOU6aFOCJBCyD7Xw5pYgMvTHkIztRu1yHkk5ub0
CYsB1s17O7S5ISsNjHjdLTfpDU848yNbzg/hULXW4eXYhKvYTxs6gI6U7aZI
GNSetxd3UhU99KlRyB8eoa2lgawv6PfXTL6RncW3DpeFGroh0udfJDuMtEhJ
EUrFdRexZpIBlmCpevO09gwhtHT7c0B6xuZyfItLCU59k8tW0C5KIJxNHjZZ
jNW/AfHpiy18dExbeGkG73o+2x1Wu4+vV7hl2x+Y8JBZpmAF6ymcACtLofCW
3jR55aX3vm/QjU/ICWoTZVsT7wYc20wVtInzN1sQJw7TjGXAIsunZ5VWzUg4
BsUtxXo7GX/OJivHGw+ZFETI12pzxtUfZeEKy4O2Bx7e+d/JIdtQK+xNibSN
tbIHR0vTIZppuG+y/Xv1BmXLgQD3S5hHxSHxEO/ZbW6bLHylT8nKnh9giuoN
HzLNDPhmCYZulXBDdTNo1z94fBho8QES1ctv4sZ9EKDMN//Cm6vx8wkt8Rx/
Au+5DvdUtol3l3zwndeZZySpnDSPf5zgepF+B2is3notMSOnpEH6U1137cOK
XloZf5O3pY4J5z2F0tsRrUBANYdPlPppeIs8GeiowSh8DNTGfqb5ZyGzL5mO
Sx4U8nefQe52HrXFyzqziQ0lRZoSblTF8tjQX4cNaIlco+p1yVWnbfEUrAuS
5K5alMEzSgRD5Enb7Rb21AtlAywycw42Fz9by7p1RDabPkBqaAXpzLCzPzug
Lu2XErXu5QBZTQKW9+9/yoJVD8Fiqck6vaZnJ7iTuTD+/oWjaf45HLlplE0c
gqlHrCTSSkircWQ/+y2avE7lX7sy4Pc3GzuIcp4ZGTa85zdrBZiEkgshriaT
Ii/EeazObV908FAcPFriYydmAaSSN3+bB7r3V+6NfOPRqpl3LVj3JemePqnB
DLtCgbpZb03zYgBk0vqTzq0tzKVbMVeWgceRjrhrxuxqwEIPddGW65IzreI4
TZXWs8NIxb6gn0kKWI+oAVKJcq8xqS1sYf2ZT9T9PovyahlZy/rR3srPrUGL
bC8BLpTfmSYy/Hh50hHdYXCgoh2miQhWxi/dbD2/UpuG64uidxPzbIehpwRV
6sYZR9xr1qxhtPkvlQb3tacFTkc5t1TYVado/DQapewO5KAs7nvhB1Q2Xf7q
8meO21OMhxfTB9byvoE+mG58MaiRAlyYOaLo6aQAYhCxRuh7/3NPvvukZb+I
Dj/+qSmL6Nlz9zKLsHqvpwB+mSpVfwJJN/soCJxHyORf8WH9zuGrHKO7nsZ2
jT4WhhVwT5boAFB5PWX9MTpFqwLAW3JtDp0MSYZaHinnt+Ogv8qzatY4Lsxl
XpSe+pIPD0cR46Puv+XvVWhsOyuKC7VtKMwdmIJzyhjc34pVel57b/+bh6/0
rkGBA2x2I97Cg/+XinIMe1mj5R1JHIZgKSSP66budiqnDGp0qS69Mrro4aCA
RrwTm8rVtAcRKDkJ2CebG9gKVtDIfmN7yqfoflCO9prcOBbixiUgA8sWLEYT
7N2YNL+iZXelMB+cWrUITG4/2nP1K4dyPkayDE/bElIFtjaHhHr1LThdJ58W
/2ns+/Beye2CnMJQkIz9iAklwN62ZXLGYtqOPqBpZuk0Sf07l7m0ws4aBHDk
M7qiHT+z7oLKWCBnKbPyFDjM9gWHjek1rSNX1qP2jHrbj7ikz7FHtORT4tz3
IduJDglILDyObHINtaAk6dt+1MT0qXeREj3zjPsDz5V5WKQ1GaY2AS01dSIO
KGXF3VXJ6o93zlqbWE1ausJ79HvrnhdPDgdsIzg83IQDghs4f5yxpzoPDUnP
mXpkQ1rA81tyMQDM4v8L75rk3r6QWnzppclLnzFnREI3ks0SjTE/3UFTwOM6
Plk+dTrbv2zH5RCGZpU9uan16G1YpB7GnWPtBfftm0lN+vvJzfko1C02tff8
T2r9XzOK2jnji83Bxdhod4d8dRljg3b3wTgS1r3TDI7ZGOqs6bF8rfqHALFe
6sqLKO5sA7YcNYC2gYT/7SmEzTl5vV9dZeUME6TjAglyuuwqmbT+L/bmlmzk
pdrrwqObHFM8kaH736YSPVa5BX1eIBS49bKVf/94YshJkzLTHfh6syJxbzUp
kQ74l3krvu6c93B1vsT7RmzYqNwHJSx0xSH6KTzqMY4y/KSIN9GmrI4WGJOZ
idfNeY0jfEAr/fvM6KQYYwxV9iXS9QRLjJZKtxOdv/PtuMj+L5yNM5nVAn2u
7q6X6XWfREPNIiVJhVXvsUiNcSKGtdA2RdbRqSpdAB2suKSLB0E07fJ0U9FV
Xb7elPXk8K3CluOInOW2HJM/8iGOcLvJl5Xd2xrkES3SjKZXh9Rqg4r/69Zc
Lu5cI1F1SDQGbuNbT4aztquqR52wsmk55EzaDYkiuZBCsvzm+BrDWNQjHFu9
G4yekuR/+GjgWgbQlMAz45P8Kqmkj6l5tAn3f/3Hz/xJWypO/yuwxPROLvHY
seinSt7WGuqpDo6g9MHXwqGlxEj9GZoBkEElaa8v8qe3oGrOe1BAy01mNb1O
WqX78r7/VJynz4pFVghAZ0h5X3CVSsIKi8oQ8O7bBgyqzWT/cG5CeBz45eAI
rcKE4AO2aSCxv5RqHideLaouuXGEuoukKVQXN8OqvZ93qlVmX12elEy22k2q
MaAriYbBzKJA/Gvs1l21WFqrAgksVN3T6tJCsg2HMjItQbIISK9mml/vFW/g
JHDAGrKcWxM7rCQ5ng6qQaCHrzK9GdxOcTZn7AjItW67kmOSFUIgWLTXqdhd
uZUdILeIR7iH2CvmT6m/GTCWPLc30cHxgpmE3wo+98aZdoRx8ngxQgcY2Qkr
OmpYGIMSsnhnheXCk8hyRXJE0xs16eF7x5lSx1FgdPi7/CAtkullPs3zSKod
6sA3stdABEKiavOipgI6jwTOrVVVIX3ZcDQU7aY9z34i8XWuq1fFeGhPNVZf
6HbfTWDoDf6pY1/f3NuiHb12+Vq7vGucl/BB9OjxlI6AbAF5RpRLV3LmDNXH
yjsJhHqudsIPNSqmj6yq1O4odxa/FIh7YJVl2FxGqfqRi/YaITVCkaACtEDZ
+ye15zB4EzgkAWR0s6ypAa6lOAmqjRQdh0QHHtQpDAwDM4Q2DaDBM00DolR9
C8/JRWU+553jtLJMe+riImA0gy0IIHbvTqAS2DPrjI5eq2y+n3TWDZB0nMMu
S8rSS5OfzI6vDYzAOZFaNS9vRzKWkLIqE+5oqWcQ1kb0LHF6p0Pj2v+t8ULM
T5dV8DDJD8iYYkovbZEsCQKqrVtZMpqnkWAgiCI13YSnotNxF6iChm/dKiAr
BJJaK6MboGSS2JYVAxfS93JLLjmnrPKk4+/TUhMh36o71A36mp+sUEn60PJb
+KbbjnfCCP/iHGKE1xdGoLRcP4LMoXrn1ZCo/j+LWc6s+zVCp7lLe8Wk0+8R
e6RgvJjOiapOaFQsydFpDzJdh1O/+5W9r0NoIx35lHWt5xShUbhQF9wwj0Ia
QwIDZyc+FONpGjqAUB9fk1iSrf/9uSRm+7/kIvx8AoA0Z0rQHH7ynR1HUPyq
aMEEXkCQU4q/6+mtF6fXLtfg7LGlwo7Dw8jMSe9nfBG8pNHOCtJaxRU5RsEZ
yPbp9eiiAJ+xsslNyeLs43TwxDSJhynCm+J3HC416aQ0xEQBmp2c8eN71fTd
Sm/r10gvN7uGVg+/lva9737yn6N234Y2ni/feDVWsElJRnwf75nSGcAlA8DA
jmnc+0JGMpH81f1JqpMYpaPbsRgt7aI7R056obHg/sMP9ip5SlWP79WozIKr
F4TuHVYVqsdtJAIWSlux0YVCpUlaEQhuYB7w70WCZD+XcdgdI5KjRDGM84SN
fkbekpsbs/5g2vhxg0mNp7xc24vL7/rmNFz7jRqRLTpo//PWc7G6t9alQ/7u
pjr7hTBMOcQQLWKwZV0SLe4igQ6Eb/CTC/uk50H1JZJuthluEhl4uEasGNmO
ihWl3POUYf5JmXGmiyqt4Bkjpe4sG27pikjcvhuzKv7PlEO4CuNhiE+GsDle
cPZliLz04GKppZbOo/NJaeKS/yTyswCLynftytELh+TGKeaHlatUMLwRsiRC
J+pmsijFRQlGENNKnp3EgNCb2yGdpQnn0Z58WH/Pf1/TbrCgk1bHVUhp71fk
ivkSr9pvuR4LWRsJfwx6/0/qb0/gXn3f8ccjX9zM/JzLRY5R80GA3wQEwLuW
E2ZeoG7/dtELXUJF3evd5SKRgtU21qxe1fFjzgHxld3A+50234x4/5nNKk1S
E2VcjCXooDH0XALXS9R/7oib32P2RpUDfRltLMWegKJsLX6FLqnNcht3LByU
pPEcxMsJkmHlbnjB9q9OOg0+kFE+GrFx2j1VWyZdbLP31519BFNihljCpwjo
hMdAvkU8oKntYCqjHVcbuAD84tULyd92/nT2QwEHIt6dULS4YGc5KqOvx7We
IbO2CtR+3+fnv84QDjiYuDo2Rs61EtgQ4OOQUVKRHT2k+SPhQ6B+23zBfdre
l1hJgzb1teAZQynK6xyrHl629oCREwciZ7YLDzWGAvBb/Tvu8aFqbicUuQ5y
f5a7Y1iQ3knmkfOLkJJhaI+6mwRlw1747q3KYPlWcNwg9jZEHqKi8w/12Orq
DSyNQf6clwZSGTRhLlrkN2IHo2PsJ4BMcvInb/QTQ5ox6i57DmkgFKka4D7Q
HFbBYbMjXwctd8jbehpsyz/RezbRbga6ccrz+RleM/H12BAzh8cs46GK9++X
1yBPPCFbif72M6yCmFKfIlw1QyiVCio7P87aiY8/9qloZS9luvHUgRgAxsrO
2zIPT1CGfcAJbic3zJCXiKG4b8b+4LHnRvvnhDWE2OBcZKWRhj4hMlHQhcO9
lsp79xpB65nv9m2MvhyUSD9pw7Mz20efqKpHVltzS0sqsn3Quqc2rVHOizsV
bXJdhfMC5i3bgP6T1Q53nCQDXf4rgIzySAsHCStcw5bI2OUUBCj/S95ADudO
wUAa9wW8TaLhlsnZoVn0jAXqlrsNtZtVkT15586bvBbxvcAkOEpfQ3P7cipl
Gpe/cZaruV/mG38SQUFWPvHGQMdbN6KnmirafFPtfj3qBsMDN0moBMT4AZEv
gnKPSf6cI3EEiIj94fJWh3mrG38csZ8XOR5vIAFBCFPTkQ8XfvriUhR9VfKJ
YVPN/oQbLpuXDpkLhY3feNnmOKohztVV64gYGdN/7aUm/pBHrkceArAkHdPC
Q9eZjl7IMFUXNJaf3z8VP2Y8vFSrobcXKE0OhFDhNzGOAP5dXDJkWpaKmMHv
5W7IXCpFqFYGBCA3hHx6yPUGNQw8fmihLeobkmbw6lcCEEGVguKfPyShIRA/
xlbcCgpW75rfGjZeZlnOjxy6G5kqGO1+0chE+0HCubif1TUMnokADY0mBfhS
18xLk06zIPk1/ssBhQw+ohs1af1vF0oEv5K+K8qD3xtOVjvfOLuJCRzDiiFH
1/skUOjYz3Ty4VLblXShrWYYXRwcfQKNRVSgFbhigy1CA0M+/8KA0StkDpCX
spQb7wtCjByn1aWLZkMrWEnz5SyRSL+P0Hhnd15BGNi5METJXBkoT6h6rDd7
qUh+GhSRhppiP/LliSL8bp5V2hRxBx36d3FARRBxhOGJxVSmtuZb3EGPrg4X
ZgUNSWzgRQXAvIxVq6i5yL6pqLhen9BZ/j/sfom0dZ0kM5Y+ydUof4WkE4xx
812mEsBibjcGmA1fVRkZvjLjsXfNUt9F7myFZNuJ+GwPw+fQhDFheTC9HQyV
iFF8hg3wSy5SCUQOmAr27/jqhxkE9iog4YpKZF1IaaK5y2szHCqFtDaYkAi2
xND5jbh+paN+mXWC54v1v0j0J9l+vHLQbXVhIIPGKs7FBexHv2Ua67qBnO1i
76+9T5mmYQLiTWkG6rAfnwkK6FO3gmuQqcSFwm6amL9Hjml1ckXaA/hZzN8z
QGtJzb+ORAZlnKJkpGRvnLY5BS99lDgn3d3D7nHmjQU+S9rbqbgKNGek2Vrt
UwXaIBAXzZGy+By5jlgIolkwi7rzLlEpCPe/eQmG9vEPrvZiJYhTqHNH/llj
o+sLqA6x18bnD5DkrYK3xMiuz3EpPfde2S3XDgQCL5CDORj+4wcF1a8anyKN
zdPCU+wjiAl+oBmqmeEYpTY98sESjuNRePXmAtgcgO5tmNCSdpxFB2gpc6hR
zYm7vOHiMOleVUJjwqV2+u2Y8bVYzugc8aemE7/oAR3hkwKZnAQD/Rmm87iF
s53Np8JE1uPNhtrz1I51m07hpeCOG4INhqhsql5NTiAk0YJOtbphEQmVGXGu
BZ4Gvq/I52ZC9nuh/zzNo8JreO0Uhvei6+0mK3V738ednOBDVCicLiXQhcyY
Q2v8tWu6tXNwkiwpEWVL1GHw0NhzQxdwWTFqkH2k3Mm8C+Al+jdqpfp/IWcB
fyt6I/mrkMTwZ3LoxiUe7LRLKTzoZCihYzqjOh1IA3hWaNwqjIKb4chNmpQT
I/xtBM8rUt5nw6064E5zFETBxJFdTG4uEcJxvBH9dmaIvMudp8WJ7eGZjfzn
htBndVP22lTB70V/745TTxgmU2G8YErT6NYKtz8MGdnETluWQJDZ0Z+RLDNe
wwZK4Zjx6l0SztKerFT2sf5oyhxxWb9ZDaJXrSITU9MRa3GivDPx3AhxtFNy
HGg0gRab0LhKY6I8YGf6ttmdO7sOe+M3daJCQDQVbDI2V8w2FNEsHzjQdz73
f+wP+aRy7syOx+PXj6/2hrbHib3vCr0RnD552to5+zUeFN18mN5O1+F5l5fG
8jubcr6k7w7fy2HWi2HxAh7zAmdAIOQ2so9VsKwUbErqaCXmla6RNPNS3zSG
0LxtDkb8Z34uRqw5yhyO4uzdg4pcarZgYoj9HgvMUHTJ1BlRAmkio3HqvIZ6
n2zvEQzZ9yrJFojlf11pX9ZDF8qwVPQfl7W3i/J0DJ3y6kB4wR8NQOAeYbgO
IxF4uGT5tojBqyEtteziwgt/NZJwC6gOAUTyzzy9jtQMw+2WniSQ9PuV2+2O
XjlTs9uFaVNS3Opx9i8In1WrRXk9XORtizmQS9b9wfNjPSIqXlWQUUzbuUc7
PrPYpVu6gZHcFfpshckNO2qRdx8qUV/gNMxKGJDjrRxpJlHAZN//LIRRWNIK
l2ymssWWGEpQsSqDbLYRq5b13gp6SaprELLIpvGI4xVgkvlmHrkCz555oAKk
25cDLTGnjDDJmWyeqXi+FC91Rl9JAMXOAPg8qjbaVIOhrMZ4SDoq4y5HgXCO
Tfgj0IE2NVFo9GG528lJx+ksXIWx66+eZdVeQloj4MWzz3YMHjG4KnZfwgQl
V+9WqD0HaXo8WdOx3s3ZlO+rq9BtzrGLgAdj+3pBdRVYMX/a3KBE3hB3Y/Gg
FAvCyeeJtzT748o4vSm5ub34JzWhCehkpPyA3V+AZC3xcW6qjYe2nf1Fe5uF
AHgpFEt4HffiCXxtGFGbxARgGz5wYJ5LpojDvk+wJavV/zEgJSF3KybuTEnr
1BXMP6ku7xy6PYf0sanQu6yFcmSn/rpBL0SA4iupnCL6HLU3G694kYRw4E5v
iCzfjaZx2QBJq/pRX9RT5KvI2vA6WxOaXN3MUq5f5l/BaZnJ4zsCjpsMRqwN
Wj+X6BCb1KO+wr2BsBqlQy1EWeclu6O6Una+7lWNhvS6mJfecUmd/sSNJVqv
J6Un20KU+WanjdJTsDoT6cqcyquT0XKFDvBbvK60Sc7X+FWbghDKf9EzAOXd
2AkTumL2n6abiLQRS0Ry4Q2+r3rynYJu8nMWV7onnmmBN6NhZ2i8MjBIuu/p
E+3IsFw7ggyD0llTBvFhoA/JbLXVzrx5CKdvqos6VvfglfzBDpe56lPMrwE3
4cs2bpSszDLHBg/gI9WuLfVqBR0a6P4MzRODKsFKTI4E1l3p20RMJhsBRHCR
kXQrZrp47TCyX6xFMdRX3/FvNpkB8b0DKgh4lxgz67L/3QscQRoUqSZBvw8K
5lbPWKvIFdY6R0QvlpZMnrCCo6Q7CGmLBUuy4s3t8+OR3+CgGuM06DRpdwbJ
/Nrzg5GOtHb8kLKg5mOfMxirPm8qLbBdQ1G1OKJwrsmeSEci0SsHhhfbo4Qo
EPCtaRemHrCDjSBivzlLa4Oype4DZ54j4Y0f4/SayF35yC7NcVYW4A/CwDHw
OAUDXm16OrAShivrqF+hTmanoh74FujBaM7htCMquJq0dvqnh2Tp9JZapHXS
9592e9fr/jr0GPlLR1ZGckYYv99lqQG4r48gpUdIY9SJuM1saKZXXzSkcKRE
PrA/te/4Fse4DYPhn63r6nuwnp0qzZp7Z0X/TERd5Kqbv0oTe8/wyk9mbgGK
DyKd+MyaQqUkwfIyDrKcgxZXItbyhfC0Uw8Q43HGIaxWUYXfdVFy3AWREUJB
Ys1o/5xAV49UowrlwvMBi5MPdDztcZtjVHyB/GTiy6+78sAkZENoypU2cKw3
QG4zzgId5mfXMOvg44o+xMEBTYs7YScUi89MEINexla13eV/Go8+xDXvtZN0
wSOvFdv/+slZNHtb3dad9KVxaFYraVGc+OeWTQHlxDp0MIiv3cUUlJLZ/9Uu
tO6cBicc3B9iatRigExPbiYLNmlAUQzVccFg5qh86SKMnJ96dF/WQUkZRGU3
8RYArHMZCtdE9hEa9Qon0C786JD9B46Q2oQvA4xPTFcLP1jiCmAWLdDhCgHy
u8AXf7OySVQiXfl2HSkJ/IzTh/hH38OXKtuHPms5k+svMtDYR8Wpo1BoxgCv
q4dXslOuMWCLFTMyMmjXxOi8aCSEIwW8c4W/3RfI9nwQPPotu1tAzhhFidai
DzUNDzRNYawS7pBAiZ0e7c9zB3MHY9wTd+joXiJcW+JPENzLv1/mcdOqizdd
qe6fdWqk1SAKapLIFOBu32dWniA6uR4IAJDW+pQG+/nqVHFclNP788qTjd5R
UGSx/xmVKmrTtKba6NE7pU1anCvoVO0RAME6KkCdqfJhYluh0nAywxFUrkkp
gOs/4bahlH+HTPBMSSvKKnk3gQrW7WjOAzfwG+n3j0JVDyzFl7bbpoxrSxdf
CAIDIs9AL8eW82IIhtr1jDiBdIi3tQeVrU70cqcKSqH7zf8xZUKhJovyEc5N
3Gh9FeIApzbJuVUOdmgKubSxt+Y5yx4QVyTJ0TmNNJCtUf7PKOsDCNI6h7YF
rmDhVwGRDGv2iLc8MgCZqc1rcRoJ2aZUbx7a99Sbpux5MrUWhnwPLqJtJukX
RTnx5G+zRb8gQGgzPSmFzrjrQawLvqZ7rtFSCHyhlwEip8bUaoswLK3SAWwR
YPo0wNuDaagq/kwVXg9BCoqewpP14xvs86wmfDLQrOaXVvdOPOnYruViJdY+
tAGe6qR95OmbKsWEuyCnEMYHTefCWwXkTPTRqY0VsQ+lCn2uz4FJCxQRvYW4
IouAlFUhFpRFQxq3stcyOFTrwean791gdRnlGs4MGXvMaKwB3uQHN2Ubhz62
xsQ+TU4jEZPFf4jO3VZ8gyCaTcE8A6jxb1xf7FzPwsB9LWmjMpAAsp0Zxw9e
bq+c12iIIC+zzYvmzJOCFNHSAFF528XXatkUIvPKS9vTRGxfpRir14x9mCn5
rMlegUcri3PvOXnjEhJaXnmL/2tSuAg+gDQAPP05d7Cl0cLEIoifGnoVLNGf
TYj2zi3gV/JKlRlkIG+x8L4I7qXn5lmZD5aEm1t6e5CZgidg+rZJgkUhRd97
Hbvb05bsgyjRECo60UdqxIdMdtqJhczlbwLyQe+ZMoAhErzg/IBn3L62Ihif
MzweP4oma7Tj9WZqsl6jiPqOLWU+eHL5263JYU1RKtPWGQQNZEjZK8KxUJos
kBmWqC2XUlKNOj1c7u/doefiRZdozDkHBryuBBOgRHrC5D7UAm+9vP1cK7NU
TV2DkI7MF14eZ0wBxFjxJKQHfkRIiHqSJKCTutUOloiKabYOJ9rK3qkB/A5I
G10B1FJFjd1sJ8t9jhaBECKRGc5f6BXPmvZZLRI4H2vJUJ/W8rZDbnbcAiAb
cYkWRBusEaQvQOP3g9OV/0pMkGrne8M/J6FFOTdhrsPOeVAa8p3Z9wn9Vf/K
m6hRFeIXzEKje7sM7y8V1OonftG4Ek+qhZK4vFqpyY0gyRo0Ez04BBcLZR6O
QvdfIECnwpiGdOlMIpMRD1tVCtfZ2J9FtVpupFGItwed52kF3XEDQNsfpQos
+7oyrnS0rv6YX2GGR7WP04GcGexEwX74+8P/8+RG+DthMvnf70qLp5DfbC/c
Y5/a4bRZBYtPja/kqL2LymiN4loJ83gWKOYWpEHzZ3t3WdjhFypexPWA4pcO
ja7V2WWET8VI1RIIW4BWb0Y31RucjZ4xF+HNtIvyzeZkWySf7QJtxoj4pnRg
+HZtml9gMWCPHYCtVdmENQwMWRbEQWZ6+t26fl2DnLj1VFubi1dZgaL2wzKc
+ofwSYtKMdZ/AAkx4Xtq/kN4PWB5TWeojbo7Be6dv6TcxNflsK2zv5f9GpCH
nj2RjspUaBwIIhgQZefvDy8q0LydopHRtP6wzApseI9NrHBzn/JBOPSnOkPH
GY55QOqbiAsSir312uy2e5XaK2UYSb0/belqLV8KX108v+9cl5p8eItLNJpe
VHF7pW7QryFzBimu9HThUp4POIUlgk4Wrq5eoV09R2K/qcz1jgZYnULSuX0i
faXB1Co5X4EoEmc/kv2WZ4TyogNndp9wsflT7WPsuNYt8anc2jRVf/tEoIJ/
p4JSuwS0Jdf8KWBLHW31H1SHz/tIrXi+clvC3jAg8sGdDXeLo53pyAyhJ84B
tWPbu8PEA3Mn8uQpjWatzeUmpDQHUbLX4+NsahwfD6aq+P/RDndtTpDGY/qN
GNgQHrLEnw2EVExaDHwDlv9zHFfeoRAeZSQdXeMt7RqBAsgN7IitMYZRP+33
yYT/zJueXI/7QBihVGnNlDzC7rGAJq0tTCq0BAfKwlNvq/5FtBQO2QH59TnC
QlSGBEqAaLJb4H7/L65jZvNXRZWkwNcLY+++6q1D1geTUHfmrBZ2+mP9IwEH
8jRVGLSN2vHl/FWen9Dq9hQtC3d9gkAEuWftyquN7iKKZlrUAZYe6dgfYZWi
2BEceJLWyk520ddWGBnudbeleh5YHPOVRC0tj+om+jcYAOoujQTntXkMhkey
USkG/BRjsAW8oU5qEVHbskM1A8voU9v4ehzo/8WSZBJhrZCUGfmTaa+iLX//
S2iXk3JLKzfrQM4M/ti9d7oY46yqPQgn9Rx5rI/PAva0W6NcdfpOtfyaIg+I
9FEmH92eP5tHKc8IPZJ0gc6ere8bT0a7hBIC8lqC/61aJNFhA5Eyr5//RrO6
B0lLsNPo7QnXCB1NSCxUueoSJCWAy+fV27/OSs2kmEZQoqoEEjR+Fm3XKAx1
spReN2Iyhrdqo2w4TERIegL9i988kf0S2c5bvecXMOkKE1eRDNZKvC5kTWDO
BEThbFy7UI5KoJKF9a9qvQTz4TJYMc8NWbpeo+YoyWQDZKax3kLWtSCzItKV
HlM7NBnz5iGeTfjiuabhSNk2FaXgzJRh0KX6xCkU6WC75vKxOfwp5jNES76T
HXmOnwe5MoCbdKCkn4gjUcA2I5ovM0twwVlZKzMEtx5hjfbuwy25qc3OFNwq
s2PGgHgy0iEBQNzsPGd4S1U4si4ElsOTcDNyIFiuhsPvf3VdYNFD+sDZ7Tdi
2XvXYtzd8p+gMVGgeuGI3FVg8r/G0Iht9N8C7WGDI25mKhcz0sjb2qWXQ1b9
YvaTVnZEYo8XrQn5Yn4frNyAyZYqBIzQ47xRmVXW05X2QQOAiO/1FnmK0kfA
4cL15fzkqWDUASmoYj+AoJjQdizCLa2LQMOm8WU3m+i+/NFcqVyT8ljLYO0n
xuwlf1u4TeJdEJiR/aZkBqOk9Ya/5HD1aqlEHE6Us6FY7N9oB37UbCVQPpfI
Ujg09/C7yzi6bTF6aaqckN0CsfXFoPYcmeMa1Xq3EpfTVIkeCXvKGSRlRfmv
SYFEfBI7Iwa0MPK4P0uYpJJTJ3De+T757cNJ5GoG8Or2ZMusbWETrmD3KlEo
wbOgcadOQaW1IitMx0ZMs+RBbgIa3qLLAPMUoQYTV1n4uvqYUaeIGxqvi/y4
grPKcKZgzo1sKFfbsvQMiJFzAUSpX2DYr1MsRLQxvr53VdjxhcI8M5Wf47PN
4X0ZPkm2Vn4PzUr108S3j5IwkW/tZtcz3UST2MYC9U/6EAk3adfqHMxNZp/d
0ZStD0KnhQ3uFcpwQaE5bF7AEUXWDuxa/6SUFX+2JXYR7VOfbq9EDvUkD3DH
eLdcLciJFAMEBH/CH9PFehDVjDzc+QPpWcp6tLOjVKHK9neafIk6eULdBUJN
67MC6ym+6gAx071SrdAZ4D4Sf28J6Ovq4Y8+OI/UjX6wtQFG+RAPdTGiIvyZ
qAZxJYDYiyzOVyDArfiNTdGkl77h/2etHVqj8bbV1Y0ZJlbjyE2OMdYbpZ/v
6SoKTb/sENWbTls1rbcMwLc/W9322wA/E+BjdGolhPaMPwfHDtrQqDcA2h2N
QFbkPCz/5FvI8N0zu606J/qbqOFZo8CXuQgbjhe2TWJ+zShk+VmFQfEyIyfW
5UjdrAOUI3Bqy6vO89fx8WMTZpXEBujXQOcNgeNHhRIJLl2PVE2Dq4QhIss1
fhuQVsRGvxV7fkdRwAV8/NDQRZ1mj+u+Z9SshsgD37YLY686btSt4nYMCQJ9
fSt+Vmu+FdXNPIZNzMBFRiNpwqbl3uXmOWRhjyzLx3esJjh2pbVWDcr/8pE/
2me0IVHpTEqEmmHU3uO8AosVUJJiZ+u/4yQn/nrCqCG/k8XWzll7TreHKVKg
Dg8M/ZB7RA4aolAxAxDVL6PqiXVcCsQv8N+nBzRAWjsX0OnneW9U5FVC18Ra
jyuNW0TmOtUR/9lg1cn+x3wv/v3Y+6hb32zRHT1SAS9cx72BYF6YI9xDbr+d
siM/i31N9AUAtgp/1I5Y/2bY64tq1x8GSZ9Hsi1zn5IDj3UpVPVPstelvPxB
X6KWCk5RrTzSii0+IZUDCH96MkkLhi/c5QKVB/l6IXvfmUrCRKTAdsTkVC2Z
9mtHaZONN1J8HPFjYb04D1W85TiqBkWpDLgVaTYQch5oYeI57vVVFEbauofG
bOgfk58OnNu0WOAmFOTkkBNDnzshlbzGYG7DDRIzuaLyuROF1dFn2wiL94dR
UiZ7cSc9FQjCsluwnI3EkJcKv7f6ZIOFHCJqqqVyNRucID9meiRXXtxS83Zq
H7uMJwH5xWwwAHaHwu983rD3nckuvZLa3PGo9NPCdh7ofzvtAK9n0/w5/syZ
QoYmILMHad/mEejoX6h+YdBMnPo7GBL6kbIZr/EAAXYLNQfVawW60bVaLiFM
XV601ecV9m5FBaGtL0oQKvteR2LCdUh+IPf/G3ZT8SzDCkR5R+VlRS0NweO8
6JgzOJN0KRmq3ifBMe48+4o+mb2I4D3HQ5Chix5BBSgAGc1CtpjO6BXA12ve
AsNPYcO8UC7ovCxjjNptOKOMj+ngGrsUAccp7nw+aYYnHhO4K+hMjgztzq9M
LKr5AOZJgTB6yqug8m3HCp3wLRrzWeMy93FsQJxQvoMgWw7/pNGPJlKG1KED
sjPF2mu9VuNfivc2H9MSV/vjV1OS2OnYEuJ9ZXSBpfRaICYv3MywD6e959cK
GaCyhKEpxUBzG4ngTbf3Vj6mc9NiPIvWwHuIgaA+iLgPR0Cxcvvnw5kdk2kM
DIUFziI55EVLnycdIKHfm4Lh2lt0+cF6jwG+Ax6CJtYt+0uV+Zon+FnfZYnk
e4DpMF0jROgL71VE1Od9g7MNc/63JUjqKbOyzOVxtVkWTFZsA2NII+eyQj3O
nY8ljGSJvM1gE01AeKGGo+EFwgiJhgJwjW7bjBYpI4M5/SVisNRhppb+O6mE
LNRKIAcdd2M+exrFHGZANsh+H0n/MXd69LN1nsynvXHSBgqKaBZYKsu2nqlS
/XPf9xkFlHNyZF4MzyzDigEOZUS++6Nam2gmcU5feBMfu6uqkm+1Fsrh1KAE
eB6ky4pjBX8ejup+4mQenkT/2JP+bCW07QDqBP6fAQfXuBQ1YTpwqqHLPxUM
J/A5W3B+wQ7U9W8GFNJ1KZXzF4PA9lGoG74HAnoIfVQ+gj7mKy8ESe4f4vDc
aOpRx0+guGdeB8+S6ycv061W4hvb0v+8WMN6DnFYjWQobU+UeVkOYe2rRBeq
z896kf2YjohTRh/hECPHU1t3cmESNPkcW9hapPg00whI0+Hh2+4BEAp8CEtw
yMcHvRKpINUErBCtED9tnMMM07jdclIoG826YVER59mz5IaIr3ZH/OkBrGIp
cLCJF7zelDc98ZH19pdUkb5c4q3yL1LlfZBJ8jrCi1BoNgBZ6fGYpV8lp9+y
M4tCE8V8SI1McrNguL5d4VdaVhGQcZPB0JNg8dzbMS5sBDoQrJyZkwZ7ozjO
CypKAJavO+0V5lVpN6fUiYPEfxmFtW31oNOI7Is9goVK0HWYyjOPeQdjWOIZ
d6ZkgvNFIq+t8/J8Lfc59+opAjLxQ6noT78SFg6nschHEmbcVO8DrQPoIpb8
l7LWVU40JJTyGmOs+J2GRAX60aTnNJIJKCvBg7iNrdlxu3az3X2OSjWc+o7B
XzIPKTK8iSLd4VSa9dmKNFCkS8Fto9U/mkED1lGjggrO8WSRWJMI9JuOLDzO
CkTIqrXGwl2QSMMFFYt4yiN+mEvEsAG2Ssqd/cWD5oA4sD76x8pjZAhc62ZA
WqTrxaPn5Xaw7rMOr8Y6o0AJBXmibapAVsGv4ZEKhFokSf/4GlDJ30x3A3Fr
57P9A9K6YwptglSaPKCjVio8HW3Lwci1gbRrpgV81i+pZwDfqWfThlyffZDy
wr928R/OD3eUTq8aYQYQjqdkDuk1JKOqMjTGerJmdi/dCQi6eNYRXFfb7huM
NK67QZL9v2y/L6pyP343IjwQVw1P2yfqPmNsdGDUfjKawLFvvAO5p/W4fFlN
l1yDzlPQ6E+qlkaIWIoBmA8feGfvLwV/wmOlvWfd9VxY4sC4YxBouDWYMTqa
+6Mu57bwTfjD8bpmG2Seg9W5ufM2cQoPzpmfEF+6xkOz2mV7K30+6gyjFrTd
F0XIyFmqz9UU+IWRRcUvIHclz8pwzGEVOHsFlM2cUssmdpsJSZcSrw+vF3yF
IPKt+d0PwDcACqbzA/ao5Lwjjy/JuwndPz4vh0gUu/2rr/kNT88LkEQkJvMA
DzyZhzdJGZDH61DGzA9Q31xe0CUZ4MuZvxm65ZuIZjkpQb7jp7zWIXEolxbC
F09hVX34iNPFyBdLdRg446hEZRF0oTUAdwWmb2Wf/Vh8rlw0u7YBVEN0ODvW
PG/lHeuX3252wYRKWQs1TBOimDWN/lPF5mrgNuRG8hRPTjx0tZNCoH+Z1k0X
CoP2lqW2awl/yc3Qf1DlIH0GGjABaOLMjO/t8im0Swk9aK3jiq05w7JNYqPR
cicY67RrdOwl/hlqZf7pnr5AXbdu0WGnUG/3J7TIEyUWWcWAeBbYnQULW5BK
J336q1hQCv2msWVFI29GtO6IBbRFL0F0b4QmY7HDOcwTGFXQNWMrheUGzq7m
+RVv4Zr9Iw65vlnWi1LC1Z6i7K3k086pLUQ9JwYuSVS5YJOjn4exCVyR21xZ
QG3qZejf+tP55arLN+3bQO3yh5qP1K/nthRkgi4M2iyuuIZeCmow5V9nNwU0
X0qQVGF6uR75cvJmREY/RJS6Ug4+FlnffyfAonbc/A56yCHDN5bCvEmaqfve
isKnYysJOnN0dJeDoNlbFzzqnWRIGifzSNPqoQ8oOUKHN9QqlbdlP/5DNegX
Z8n1XqU+z6n0euIdTRUiUFr2Bl0OmdSLKtzYRSOuzQCCf6pe3GcKpQu00U28
h9qttcST4sL1Vs0Khw1G4BF1hpZcmRXqRAz6nwq7JJQhcafNySbF3iGmJBkk
jXds3/bWzLC8Im3aXCitUMBsF2zCV/rmi1gzvRGR0CaKD5+n92UNfZ+8t3i6
T0ABGT2SPslwxycwsCKFDzQ7JZap8Jkiv5vU+KvTRvXXqVKzPHEpbdF3k2sa
8VVYiT+qM3906UWU+y82qkxYdFtJsjbBnjqAA8tbsRMFDhbR/Lfjxs+Vd+Iq
esqyWb7gkw7uvZmsP+4vb3Wp885FdPZ2eyItMqE9cXk79ZBKad55/wGIUCg5
VgtM2uk2oKOPr0VLpWPRloRmK0ES4Rt6/nxVMBFJtlmlYu/bZfs84/syn7C3
0rt4fZ0B+lyRC1JzgcQgkKin73sSWlrrTCi+x0A7QMZwImZx+dezJ0ZhS7rk
VG9KZb8FofzdcEYdWkS3jH01mmd0wxa4jQZypJeRjf0MVLEdYizOivXDKtTR
ftTDf2a61Lf4UiPO8FtozyRyr3alIexNdGLVlLuEe7H5aGHCas1Ptxl6jSFP
FkBDoQ/rSh8CjotXyEggd4tAikxfIOTXH3/4siYxi04zg8PoIe3mgLhyEk9z
NTTA/Z3phkv+miCx+OQ1rDdlnv5M8/QJLjLxRT7lfUJI0LDpuPNVAS7xKnVr
pm/qSDc5Tpbq/i3wX52IAt+iTCv5Tr+WvEcMMhGp8/oqpXmQHJOQX3tQUM6c
ngyMPQifS5LSgWNf+Du7FxkQBDPOn+bJJXdQHrCKtyhevT1b1iTl1ZTDlrv8
mk2Klr3au8gpV4CdERu8BzPVUMCKwbdcDVnHSMZnM7rjxs+rKpOMXu7EW+I2
kHgRdiavjwLc4HX1OGzvtyJ12g2/FeBIitPrjCCYv6GNmzfwkfpfMHCExjpT
cbF9NFmnXqezAI3IPZxqhgJRXmKQmafk+WfPVppAigURWqbo3Yxxfvl5N5co
KXtaMGMO5Bp69alg6OpAzgL446DK2CNKWgpiFnnX8S3UB6eAcumIZxKg7WrM
m9hB9r08KjJQY5N49j6sV2Gw+wINKHiZcA0hcCUIfCBaIvAQqGIm1an3B6Ah
54HXBb1S0hi6DvPb+V9FsjLwLtWJ5XizkEgt0k7Twh9xcYMnhvAQoq5Y8sVI
jMY8uZHVBjxOwhjCICrTMNxjxknOmNIec9cDR7tYl8qqd62nid43EjdxeBFw
g1hR27OGyFUFvRVxWsyRaZgOSRYOpux/Qm38SmRLWQ8hseK5E0EXg9IY9vCz
GGXmkmCmfzV4iAyK++5i2c8siEj4oDXObrSxCHdRuxEkRGGpQ2AO3FW9GT/N
XgagQT4kOVYWOOT+2fOpwhkhZxj7dLzJkLfPoM6OZYIB25PW2kLZNthri0M7
1kJBhps6a14LuVSYO2GEzMwxwC3yh2vLRF+HyP9hR4usRlBdnyqkx/jHYVcT
bdI2JcZ/4SI9OOxQHa1PueDgdgF1GGnT8qFsLLuuL1wZVikNzf/Aa6swXTZE
e8t8FyJd/j4+U9BAIAzpc5KMr8vurfYhdyP7GqPJGRjJIgUezKsUzRhPwkgO
sKUCP2ZnL5kImlrUGl9SC8ZkoEQ2d+er1GMdH0BMI3qUAlo5jF1O1Ma0WZcb
ilpQcNpuTJBs+bakR4gcscGfIZ8DusdmjsEbEZv/ABNwyhL5Zi8uw8N10ufX
7XMbmjpBHmju6a3ABdTwHWU3p2cRWx8hG9nJ8BSoMjb0ghIADIvFnLbpyvcm
2yavp4ZpygFRwxcsLrzWkLpfbUMXUaV2SlQViID0EtorkNuEdrSu61Jq7UGT
mPkSnLp7PO+JjAg3iJDZr1nI9wqP7UlCa1F3HAf+2pt1roisR90BCKM24hIk
mLY8uTgEeHT+YhU6kExXlweW4BggEzZ7mSI/g835BtLXz731wdv+vPpvUR+G
7KuhQ9iuXFP/F7K+OiEqfgIPRNi3rF2/CLYW0VIRBH0OcSeyZAtoTMeayVxn
uOLX9WQ2ykZxMHs0OPoARzkfa31xabnBDJ9E10h+UPIq6Hi9J9JLhtcj2bcM
LGwF/yp6t84nH3elRcxsxGwR1Dnn4n/ebN7LHQ5Vo70EPZ3+8HEgdvSySKUL
mOSXuR3HpFv7JOTLiKoRsK5D/bJAqYDg5U3Bkv5b4iBkggwaECUnJkb4bMtK
24wN8DSjUt8ZNcip8S0qnN+lTAhDWiQ+999MB5yGTyxlwT3HveXrzusAVdUk
ufcIPCaVm4MSPqrkT0IQ+SCzux3Rj/KNbvXPtpF0+xyfwWKNy21nORgpRSzF
qjDHvEo3OEhKLm/PphEJQR+IHmwkstcGAaGGWWICdeEb3UT2boRoHtD316oZ
1IP3km+loC1KJ8emEk5a/EAH5ro6X+xu6HtL8pdxzcK6FLp4E7iGC0h/svXy
IALBH3e4z5CVyHK4MI9ugK+nGfcrLYmXynQMiCMUJP2uWeYw8Lj8/QSBHtVw
n+i6nwggBvIupOaOqJhtD1M7WdwbCK/d7ApCrArYxHwb6hITZP3zRFxc88Pi
KuyW2SZl4EWBC8+wQlt5HvzGKU9IMM+5/QMpQB7k1YlrX6+pSDhY2qmHDvJW
lj3K/pZHswnsa3oXinnU+neMW0saIJS/vD6Cga4USY2qs9uCI/Q56Lmq0qB5
BmoZkYN5N9LiuM1FcQyJMDPd1GWMlLSOUDq/wbyAOHon4lCW3Qqx/BEEJKB9
LPGsX4A6Mgm5tbJ32VwvvBku0Tdf3sJiyPMI/j6kaFnHpt9QU2e3oIBM4YuN
V4sMOIo+4XZNIMtA+vIPYl2OX43RWW6jWB9YVYIXkI5Slzsm33otuWISYAz3
Ot9HZDAmr3T8sCVYq4liAFso2BVNQjRgEpS0vchwFWyzRkLcBDWsZGbjZ2WO
uoZuDIWALsF9aASJNXWJOQYuoIr6Bi/mG6d4kn4v3A0qMRPhaQlXy1cAtMQo
rwMRlNaPN99fyD3NA6G3N7MNAhXvBCeVkzFUsdUcWldbJVMYZR5rBKJyC7HT
3OuCbYkGG1FW/zrn/KlfIecwjKKb85XtqrvcFmYGsRgRIqcy/Q7wh9v62Hqp
cPYU3N84VT/j8OR4s3TXzSDQIhC7sB/vRxb+a07f2ZP7YsjtwasjXb8tJvn9
HSYBRdqkAPFc2qcRyF0hiEu+ar92PEEfefRUHhFdxrP1JfWwWRzOJRfBaELN
5CryURiEdJW1y/nsnEuCgQG0mAs6vscXkJlkrRkuZnt8Jx96vOjAyXYw75li
vynvIvtJLUwsbTC9ogIQ6zPZKFcNzDUzLdloCwz9U+PMfhjsy/xsf9Ppf07S
33BdW8WODOoA4HdK3V6jchqrEhFWMO0S1tiwwmK7vi8K6xiTG3LWN2Thv6ve
Pb2V6gRy/TZL8lBoAPT3r9oJuFJNLwLUVSjyTVidul0cztnBw/961Ul0uCKo
nniNM6IorXBBrdoYRL8rhSNKkBfJzX7x2b50QZMcnPr6GjIRdEqgsAGxDpVK
jMXc+Q2ukOjcBYdZ13PbUh2OYsMBOphRFuWL4kVLspbGKgOqmgBUZzn3rGjr
6cXyM1s5qcPPjyKsHYMOulw+1ag/pk7n3ZG32ZYy598lc2UIuERD1PHByWCM
yHApNUWNjad6Xm9G5q1enMZ0embF6HgALZt4Mf6UzkGaJYHyB1nXAMfvXBk5
0PDxQ/sWkX7DGOW5kg8AmYZaUO/IoRacYzoLqLYRCghjS03KXe+Wuaznzxtd
b1ohtZPylfJhbWv3ocf1o9ivScpvjYi9dvYGpFbSQNL6G0xLsY+ufVWnEcdN
cRwlk5odnewnhvDMVhDa3+Nu6lwOW02sE2XI+syySJa8CfHkT/3zHs5Fr7eZ
qC5SlG2yXrLysXMdqdOl9LeQRrw3SnTasBnHyGktfbDcrWIYP+AX6I5+EuTp
dngX2SOI7GEMFton6JboPjAiYLKLlETu8j+FC+yGtaPGKhC83KXWyfZM/w/t
sl9cFJcwyXXM4g1ND+YnfdSEez+87Gj/sdTNDlU9nShwOEFOLNX0whqWoDQC
IC9VEyEIlH13a1B++4e4oSeUqTZjH5c9XYXfOie8DHW9w9AIl7B9F9tpVlEq
2AqKhLQTbMItx6Tlc+SB2F7O26AeP37qZMdt+mCar1V9zxWh3vz+P+9WP4KJ
aEZoJBSxok94tbA+6bEl5GrVmCkMISMCc1wkEeiRgLECvwQ0INgE2G7sEl8b
SzhLGS6V/XIFJCWXOmTxO4s3Ix7zSucBxRDlzjqhNAf/lFezHUhiTH7Ew9SB
++rmP8mTxxWs3NrVrhmY3QXTFSPig0AReI3etpWnYoqArVPouepve8cLW9L0
UJzLuiraiRTXR5oQVJchsafSa/c71+Pf+LpGEaRTr+mTnkXGVseWgndh1svd
1FrsCz7WjJnAXo0cY/jyFkFd89qObLov1Zr5QBD7udbH9/OHeyCR09mJiYfV
WajTk+AAUlTp9KSq0H2Q/97AAJjGDuveSCgTpCwSvdjPIx8hu8uAk5Q/S2CV
xzH5M8ZrYq3ihYFHID72Qzc4ZmZbfnJX+oJXy5v2qZ3f1FNEEKJjk6mdayXP
xfDzkPdN0+eLkFbCorMfIBegiPY6XegmmOPJMgFp0a27Lc6vL0FuY3JGplwI
yAuoh5Xc4nabttowqz+X5fRfBhY4Ss+eEyWMwhxVqU4qWLahTADU0v95ALyt
xNFHWsM3GIQ1tFQJrWtdlUDMkBrVKalukRpx1dFZ3sHVyBO0qY6V2xyE8hTe
uCuyzHPmQRKN/JfowjXWZC4wMtMhjdogXQtixBUIDd66rmJX9fVvf98jTfrI
X75y6Igxiu9szOSfNNviX64LxAEUYXyQa0ubuH+DupE0xttXOGksABfq7SQC
Vub4nQ85xnNT7VDjQTQKtYb4fp04UiGKThJnVGO/CVVOe40VfvEeh8vPsJp5
z1HKm14AHrtmXZn9NyTMJUi4bmxlex+HfzgP6HxBocZ+I9IwOborsiJKM9jZ
e5B6MGleUbJX6eY5vYSt5kQtwMYb6dyNxZScznm2C5om1QnBKTTwjZFvWoXw
e5aCcdIIolYpWBUg/xqpa806JLB0XqJwA7Y/vKWWky6YS5WZKJzjyDWLm1cZ
GHXpaHYN0GlYjx7dUPY9uDn+J0J67WuYso5d6Tla9WgN17MJ6tWNHsDvzE7Q
BJudBlPlEFMlgxj+A1lB5u3Dsqmnga5WHOoEcJ8bi/Xpf804E9ZcUiqB42RO
8wwhvIPTuB6dfCXolHAYWW6MH5yL+seBFRV41VBBSusLZnKDGTgdzp0Y9Vwu
DTTp+O1l9IB3u60flahyqHPqt2S0NjjhKCmWZ1Hc8u/1aYoI1EaTI0Mois6z
d6Y/d4pirMUwbYyHiWOiJI6Q+rHKqsN+ybbhWBVMYpCI8OdxaMPOjMrurd5H
muCLRyy2GhRQyQSVssx8ioEVU4RHWN+xsjbbQZPkSm7MF52sxEqZS4BJ7h7Z
Alve6PuTXny1tB3FbMjsCzzt/rktzt7DlDrzuEuzAVJn59Qj8iaDODcDW2ll
Dz8/uBjIKmt1FdGbPsMHKSM6SBfiAy68ZHwWQ2/+Gu4EX2XGdOIjIVPEatgD
wuPbZEPOlUp8MPQ/y2teC9weHdTCJBeYYfzpiHXLMgXt9yLF1zfXKBCYYM2f
qP8wQ4Usf8PinHIJTSZ2iQYlr3Hi7br8wiBA/nT1jUYp79ixsz9nKu+W8wao
hkQwNazp1qNvo7gPSegebMN51eTgBnvZwJZV73AmlkNAah/DNOCUG77tSJbo
CmevRatg3eGWXLvcdXoKP6ZuX76x3F2Dnq9ONfl9oulXymrhmrjcc7tv2pDl
OH9bW/uG6JwE9OqR7YqGXkL4nBrbcd27EMZ7NEEVVCnOEcUK4hG4yuBjBFCs
clYu6W05Ng2NtprXPFv8VBSEpSdBb9HWxAkTA1wm850v/CaoDDQYE1AdUCjc
mRbr20ld3QEMdi1E3lyy5+3H0yjkl1WdpyzCkToPCUHBPwqO41i+M9unjqEt
ir65GdZzZ3BFybnxm12/79FXqMHTDbls5BY8ydOG2hIJtTq19HZDVfMTEV0h
AGbhgL7GlppAxEiItdsUsbrRXze1HrXXJI+l+4ZHFRvVLekbHmy0/Vm+yfq7
XfcISfpYd0lOItXK8budyqE6D7fGeAYxelvbdx/dWDeuoVG0ywkKbeR6JgQR
895pJ+BZ4sZ/0lsMLTLYkGpexP3mXe3UK778w/HEVU3KPpDTDSxHhRQUi32O
b83nVPQGmFifA9/Zkwq65bpCD5RHgut3KOva/svZc7jeYWOfjnrH7tKwraZK
uP/kE/lcPrJVYv4LX9SgThK5L1+p0Bha6qhDT2jbVlDEg7/Qr7mI+6a8KJGm
Si0Z22by5ljYChmdIu7/9EehlmXXlAh6uEJWOX6ot7UXJTvTK8i27bx9dpfi
Z+qVz6GlFgVME4Nbu/XoPXF/XPU9+FUEBeCHUTrhiZWzZPA75lWf4Sklxchz
Syd74EAYepzHEnqjA+2GWPnHUkdPAM9YYIQW05oM0qQeZ6dZnqD1O4rKoMPc
01cO+0WKF2LA5lZWKvkqwt+pA7jVGHkR2x8ZFOvqlxQTzYRZAZ3fcfe+EQqb
a4psnzKBg/Il5F58qaVJTGLX5gucDMHbHCIqsAY8yur3tLwbQoFGdYCB3itw
2NIDYca7OCwud9g6RW4RTKqTIZj5n9nUxA0ZHthQ4l3+hpn2TckWzrDKzC/i
/QC5RwdU4GAfBMNShkcA8gZ3nQP+UeiQLF2S3U48hKrR50uuF3PZbPYCtDKF
u0RzkF33HTNizNv9PiqLmy9uiw7SgdhrTGpQ2SwX/NL/AalNapzbSAovBGKK
rVXsmnnJYRCSTV/t+3vS6woKDX+lPsLsX/Oyo7EJyWh7J1EXqa6/MQ6EL95n
cvs48tNxllfRzXh+p5/0/dCPlifjQIbIcdUZK94Cj4pg7L6vtWTyfZ6pzNkG
qI6Pz8O5qDQip2lMogtjj+dUdxv5TfU82dkxgKbcAIzVs8CuTaHYgQsxYd3k
xSMuXUgsVRmhdmopaZCRh2nLhfNfBoytMaMJUFoUO2QglOw6eAbjnpGRAMyX
+Mihh0CrxpZLVnaPEWZb8zhAvMkvUmhWgFSnE9zPbdt0IOAPgLNbqJ0DgoZx
rFBzw6w2tmN1elMcEuHf/tD7XM8vww4XZR0ErTFvNdFoEFi+dtx7pGJy5U+t
ZzlxIPgUssTMuosN5ie8vYFy8eo9dpfybr8OYR2oREcYR2+21h72fy733yl7
k91nQzusagroj/oUAPAFv29mWZhV9wUwJHEeqGPhvT+vuqqFpaeWEgql38fK
uSEDdv0m5tDHlUSaiEHz27zy2XuPXP6uMir1fNJViwZ89nexRlys1OiyPW86
Lh4cTWpWgfXKVJmANp73aOmsKfqXsoYNdXpWwlXHXjWdpDrPSERihegNqfmV
zLHSmIct7ILhjpnEJgS6OCH/ju8r8Md/6QC/1iqClwnfV8Ctmz+fZrxmCiK0
nCFsGS+lQfSPmAN4eXnNdBUw8HNb4Pszk5r+GsXj23+Ya2LeOD05eONIKvlG
QrhXyYc2N9GVn/y65WVRtbxqcbh3KHHq5eXpTN4Iw9u/BwSo4Zka2mnxOGDg
UVd2goWBB7Pv7Q5qrgW/rqPxXtSA7MbSfqT1+ZDWPJffTg/+3qY4ldlKeidf
Oz6gJ+hCMG2ZvAkuePPQp3DpbKnM2NyOETN1cizYAggdCo/b8pIvlrdDxZ+N
o1R32h33F2bJrNsZAqxMEP9IdB0vmlRWHudPFdQhwxxUwDB8A8STzm28J54f
ky7HPaeOjRIUaMqpCeE+qdb2z80TttC31FgNTNsjE/UXG9fqyiYYz68o4sUO
Xa8Gbgqfuz154CurKsEt06UOL5eXkwC+ONpDY3+kR12/XZhvWuDeLjRFLMvR
OXvtiiAfZGGkUBKT17rUDTHEjdbiHcHpBBaFzuGhvzdO965E4lqbuYHgAQ1M
2nNxiDCgpM2xrucXd0NJSFcSaDeRo6vzYDAQlMS0o7G63yrig7C/Z4ipKRdC
56N0ZTyaIxxfjBJbfD0xrZPQkqEFf4HpF5JOgy+xpNtXZCfnxbwQS4TUlnnz
yWnmKnS5HKW/N99lR4QjBPeVdJ+J4ufbvhtVCgLDZuswzMBB703jrZxqtvur
xnq4QI5G5ZPyT22Dh6wXcWirpJW5arDDU8MK9q0np5a7iaqzBGoxoUp7C6SO
p06amuqZ5D7hlIo+UDTo72pGZNg4f8GQ4FdutKD3EN27tGV5dls1whSqpSKp
yP2L9zJXUJSEpq62FdYCmF556T4catE0U8n0VFLNXYCB55c0jsf455eAa1b+
RtJJXxWfkjCwSIOahlHCTa636ddFtoi24/X6ampT2nRze3Y9WYOAJOOpJS3J
zdvXnTrVFrf7icNuEOskJL833FGIFj6W/8FIluJCn8Qddek3PifNTGIGsgVz
mMCltdoLSuI7BQVGEZXpaJF3oPJJE2/hXBT42rOOKgEsj+JEETXoUM/LCUij
Rpt5nE2jvnLG9yO/IOHOdyjjWgziK5yzc6IexgdyuG4OSGsXLsUU6d7viuVY
lLAM+ewhGuT0U/q/kdi54by1lf8VGOW3MzRVkNo/B4UMk4ye2ZG4RqkJO87Z
05AG3C0PydgGBtsBfEw//2Ada/j1r6p9kI7+X694s/tfu5EuWftL2HVmB/kJ
SrkLWnnDZYiCh94biUz89BWYqBd489Ryf2L2eioXW7iClN4NLUbd2OQOVRqB
z45TVXYk0w/C803uC3csvSnMxU9grVqxC38ckZxb4mWV3Tc+ASJwfXiY8YLw
JMTz982pKu6OShtJbmLzTj85gx4f+wEZHRp7WTKFkQkmCIg94LpkvQVUJCdo
mly6EsUKUTyB05lHTkBoH+ccLltheo9K1S6dBdXWEVyyN0HuBUvHgi4hqhPJ
Fi00n6Z7RLGi7J0PTPRCW3aLt7ifIMf1bAa0dzfm8KeXv0bx7WtnYVs15MDz
dnn1cwOGYS9/5D3WX37lYz/3M3g+95NEZAyQOZBA7WRAE/Uq7Ap5n3kVeDGt
7hnER9xyUhgty5ERZUCFVdbk46RVT2aYGSMu/m2qBtgSOrFfQQmOK0FHHtT+
Wze1uOAPXH7HvwzZO4q3j+yPCkVXMLjlmx8Ot9kpcUOQfGAjHWZB+mZvEwWa
SlJlht1juNCpUW+PMIkYH8U6s5Q0e2ofhIZuh5ZQ5lS+5MEx4zR7iUsnDSsC
CsIMw3oR3SCYbUgRHhf6t957uUCXpqKoR/se5GUKgslQjXIGaceGpaFE/Vyp
bX1T2m6b0btLaOw/C8R1lIwr9jBaZuhyTFQsnDX9dLF7Nba+wwF4PCh5VC6k
7hv6qbeyoEa6C8PoKAVgX3lqsHQ+jUDlI3nqiqHjsZh1qNQ9FS+BrlYOeCua
JV/8iQ7gNBWlrOeMSIuBg5I/XIJTWLTBymi7kNff/ifkKoBq5Okz1DTD2Jyf
5rV5HfgwQK2aOM7/E6H5dW/3tdYUNdjZdZ50Lo44O6JmWsuZ40+1zq5FXcjw
+NEIjlqPxzwsGYpwyZ5A94LyU6BOXwdvNFwW6wYYojIqbnrLIuS8X2omxOOi
gLPvrrXo+rgdlIOu7f3g0Q9w+w5P4LObA52Jz4XBHWVcwsE2LduNm+hqbLXz
xcoB6WAdQiNcqvbemBBugGOjI+2NgjKYo0fqIX+fMbJm3FuZqHvy/sQPEPk4
OXBzxHoL3Z71TWMdoh0oZOQ4paqNI7gZlsYo8IPUax4eNDgsOs6k7rxgGIJr
2ZvBVZ13oY5bIyRshW4jWvcJ3BxH2/K2MBO7X97cLPH2ytD+jpOKPPylTaWG
PD04WQaqpzK8F1R0kWV5thYcv0C10u47hZZMOL2WWY1sJjmArCV7ZJ0Jprhc
Lp9triV2q1v+MOJ/J1cO/9EGdMvi6uJXnzm89BvfKIyKmTPchco8ab/oyC3u
0YFnY6+fEuXxc6IBKkYZpmxd6n10ZyzOhdk36P0nkIoqebZ+NPqKEE7WZVZ+
w/JCn3MwmNtjBTPmOV/JxGuXlSYtS29lWGES03WzsMeIkGBjehN8FW+X5pfN
apAYsXWeMo5UuaAOOKMRIul0ePQLNscQu0LxQn2/FggE43sXwC71BKC7DdP0
W9hu88/f4FMEYZ/qdW5g59X6SJbReGrMOzHp6ptuGx2avKYUDAN+q/IyceGw
IBjSDhMtCOqJz2aS+f1oOdxJ/8WlTPaU9312z8z0ZAnrX+CkVwh1eQokES7H
UMARrkoViMrXdFzPo5zdUne9UDpoBfc+F7Gu+Yu1nXYvpwaCaLLRtIUG9diS
scFUABFEjg7B6WLsaFgnNWwY9d1erNDEUpGfHz+pvvAH4Q+co5YG6uz9sA5G
WkMMuGwv29qat7RW3+lGubYvGzGV4F+eEVDJECtwaety46sRk/uBFBGU0OGj
/c/HbeoJZhC/OYkxGC1pMDVfo2jk/cN1hksyUpgsp0ictrwgVPrbDAG15yxk
cpH4l070nT5ZZbhr4SeET9ZRkjyjpZJpe/oWB5RnGM4wfkseKuSz60sz+iqs
/WqvDGDn+U2ySxgWstyW0y4yTu6mnRUEh7p6dLpNyClL0DTXM0fRDjCueeTh
8sS5UxgQwpT1DKYwpw32epVqp1pekZFpGKrfbBa/zR6X/tmQ48gPm2oC/Zv6
s6mEFhfZBc3fBY4+9fFuScKWRVkTHwebdCg9/XW/z0feTJDJVWwHMLaUSygg
mBX9R9FiEFUNv3RDXnspjM/JRY6sAShx70YmK8fOZ6OPCyawDcDvlAklzwIT
5fjSGR5nA6B9tdVYxJGRP7du+N1xpyg2rC+ZszoNooM9ABNhhCMCYPMDe/Bs
qRH5jSVoQng1hoWWk//YdtFE0RVyhubK1v+b4eFR9VGaU1ah+Gm6QWnYk4S4
N37CfxlAIWEUfozf4FPyXv50fw/mF5tF265bkDTewyEP57UyqzlMXy3fjmU/
FbW5JcGey5ZsfrqiAKaEAZ+4wNzuMUBKA7hztRkt/XzcKtbivRWP7fiyl+Q2
LWsED2vraziBBt8vfbTUJYJgkW5WxEGaRDK+1yZNnwYXJkxDuMyZiIfBYC/9
KQ3c5izyQ3c8ZLMpH+KuKVuYAqrcUh5USwaDHzoBZZR6Hf0BNyV8TwLdW3T2
dFdy/oh0/HnTSSBOGSAFLg4N8yk3RL7CSNIoFxWqeef2vWenKZiJSbtofjnn
9ASla81BAAtCSPH1twa2nRWL6ynsPCCgc2sKD4Vy2Okw1omLbc9s73kStOt+
YpLJ0wvWCBTjNd3EF82CCVYu+loXeY4z0ogPorFf3LHCZnFFOK5+uUwAYmKd
vfxjt/u0KXS7nj/ZigZTzVjspq5DIq/q0cHAhF0vCI/JUIIZ+NNpkqIuRZ0N
zUrT1VpyahpKZJastlFvr2ESPt9JYmkgZQyBj5ANDJ4CzFNs1UzXv8obrQ8b
yhcEWDnWtdFT4rOqIPYECzYEEDJ2n852gyIXT1z3+lf5+KzrvB8tvDB+rQ+2
ochz/31vOssgOGWXpcuinjIX3aNPOEPLrf8sAGkvPvAjIZryj+CwmVSgqvV4
rI6HtIOp3aevx1/ckKBUKyCo8COuajpqPihuLCGNeEiOLx1k9+2V+wcAi6AL
Sa1T5vSahu1OssYHQB+oHK2bwcKKWYZPgbtR4/qbVsXgiJspoPLD94MGkx7/
S3r26oUUvkzwPaO2RFWzKDvNw2p5+HIN7x8a3oyQ1HzQVVFIWGDKnt0AG5Bg
E9RIlLRAtYkhVXmYjvARWbZ3md8Zi/jymHgcOOmn7441YrpCDSfP4e/1r52w
bMsKSXjGyA7k1iT65kP5+LSOXaXaXt63rL0uDZ7QTVWeUr+q5tB5jJZCth/f
5Eod1HdoaVNBouADkHcVHRlKUEBaSc3XJiwO9XqecMU3QmDroxKqdL3PnDbu
GTX9ix+li2W5uFMfaUO+4pABqkyubLUHhbIRLGHMxLqA8ZxnddZ3YnRV9JFr
d2Z6QiCj6DQeT9+CmDQQw7G7CjXLPpaBtkCRPRiUn/Czab7qOPHBmmS7IP5C
keHNWJJT7h1n/qD+LTtP2fQCHJ5+SjljY6HP9xQ3DhIIWXMuq4ykEfFR/M7b
+sCPdrcoLyXgTAmygh067CoIM1bccd0OSP+D81IIufjRKZhiGltTexweVV5j
09sqWtHtpmRr61IAayF0J71Dz0kMRpQsUx4yo9VDejfNLYuTPxSQC130kh4V
F8cz7uPP8WuqHm4xqgDzvJwOXt8bNucJwPfHsedJHhnM0o/KboDTUcgwhWWZ
ckzwwVKdKJNA+Tssqh4+iqefQGJqaCdgTxoVQsnEFweF3TsE82QlDAjms1IE
3p9yq1O4YG3TEO9L2UWKEli8fWxDDpQdjRUNKIwRaO4Nqi5A8fVtkiVoeQ/g
/ykZ+nk3dXQTR5PhnaiUYLagt4qlXQH4QCTwNAcYgQoX/6G6xWyBVT8PIKfd
gfMnfmOct6tnwlZnFe3NrSjSyNimcvg0u0abkEx/nGLFXKRhVe27UwnDlvBq
9swmsMsvRZREyzSro8FJC/WbmDqI8UIMXiZk/bwLKHjzH9jyADWm4c8CfhW4
M0Q1mZuSgqG9YHRBWQwkLWRunuj1u/AWAbmoGb9s8Ff9EvVuT8oQsY7ut827
rE6Aw/mTRrt5BjHZztT5mCkvhSVJC6+Nn/ArYMZRp81pexaQEh0kvlGCyiUK
0bPdJGTCnoGPljMW4H3e8tQk/FedDR6R3pIS3ra9AsD49l8NGanXq2+11Vs+
goFiIGVLPHaFK9Nm7dJyyRL3puJQI1NqfTwn3G1tGoHCVPVb5EdYtyHUfZiV
EBLY9CSZDoxNgOtyGvifV26ao3ve7STGFx5aPZTuRSDxf6pVEZovZObtorPj
Qi9HQbzkBHui0gIeiErY8clWsVKUTTAOFQrFlvZ822u0cqIYxiUG80H3tn0W
h6n8SS4h/8xEmqZCyPaOAkH5N+e+AdgcdQpAUwt2UFD+xWOcgsuHMYHPjUkC
x669TPhqJX3nvT+bYgVxFvQO5MXh2ASDNTvk/9qZolzsiFflga2Qi9EMc0cj
LqcHRh3zAWggBUegsQEIGuSmIzcBrb3otBzrQ8Zf1nCA6fKmlQ97ZCGv/Ffi
QZxzymY+zJRwkz9K1lc+wX1yjfySCHI9wwq1GG/bt3qAuVFvibUK0t4FLWS4
ie1yLVcdj/cGBEQbBK56nYL5+iAinxaCa3RdBibqgYOww/AnJ+uz2GxSFSMl
maUnkLn35CWcAzNJZzi1MbhCi690Co5wy1m8UYnQYzQRiZOCieSmYUjfvr4c
O6oZoSQkJBFxYUF5UgnwypgsldW+PN58JHjop7BI5Fu5x1E6/2npVNT6jH6l
cey1LEBjz+3AbY3wRlHvJTsNEdMjKojugLuB8Wni6dGHb0YhgMmdl6mrSMXI
gyQLGpviMeX/EDllCiQ=

`pragma protect end_protected
