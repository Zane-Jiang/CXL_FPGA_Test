// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Os7OYHtuKjLxo5SltrujDljls/eFPl94layrgODSM1f1PW9MycU2JVWf22OznAJQ
cv9lAtRU/ImRvr9DRt/k3C2lxSMOe93tSd4JncqdJ2wfvBbyyzzHSms0mskI267d
MyC35f/Z2cu+MAYbFa6ui9z2ZfIOQC8FFL5XKT9OpyY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 26592 )
`pragma protect data_block
xdwl6h+NfeAZlA/P0V10YwMVO+SyPpzQCnsZ0VOoOgxz1VYpltQhb5zavSEHWKlh
qfiLM1GRB9TYf0VT19LAqRYKQ3DDCBVBEvQO37bTqQokqccWrfg8XsTu7F4ytOhJ
InucyYV+qVx0FHJsKkiFo7vjFreK/lOyUyLiDnIyBhh4RsaAJ27qfxv/RGmUg7d9
BYF3UMhm9yPH2mjV9LdC/QMnlMQDQ1xhGKnChXDm8xgO7CfbgrZadWoFYdBwsF6r
lCJK53zsbO6AeiVxKbffQhNVc0NMeHmXJmf3sVk92Ikki3H9Wcj8ujw8fBbO5+sj
mxXShJfNapuCp95q3F8pJAhu//mbzB0esUiPLehHGSq6yQfuEDflL5K8xW6MOsvq
nEOjtvQ7YZxjheUlCDapEPJOlgbw86lTeNZClfi8pJs8Z4vA5oCUJTgHye9h9ECo
bmq6vqXXYtkYTcoyCbXdZHUGWFZyFLFAz/jYYPVSIm1ntYpUujAuG9IQxDT6sHom
rNzXx9luGn1n+DlQ+F6WdE6yR+xpD7JTco9a6vqWPEFpMjaWs2upWVgxtZ/rY22N
GHFa2Jmqg3vUBPCI3tzwv44O1EK1u8EIRGPNQ217mA6Wzf2SFORBlPfljQHfqQF0
jpKY+T7wJniAR4HfJlFOHkrv6dqrtCOANETVXlE8VWobnyGJZsPgMtdt/tu/k+Fr
NflGoSg3dYSsmfICC0vApoCm/xPtCePOe12JSWI68uEx9gf8U+He9fqNPHPGlixV
zNIZY2T/Ra3p78rwNvR/wMS3GNEpF7NQ/iZbInZgBI1XJ3hiu/3ojc7drZmBdfx+
mMkxjvsYFTQrUkiFdZMnvDzmmvlUWp9J/QZ1TW1pNFd/rsCqDO4fbLuqVRYWTg3d
jcY1D8vRwAi3usnV0by5x4URdDke46MsdqkQaVN242SvypPsmJUhkP/j0t+LbEyQ
cUiNRK1Qysu2R6da5CCN55pwOt9xgjjsOG2AvPkpJ3tG0jGq4KuAS3BCS9Sdxg23
JHb+xKLyl4PXyKJLZsJUSmjJubD2XOPpeOXVekLm633zAXwgsAguL3lUqbzPWHwr
G1IY8CYO2fdjiJFD/nDChiwptViQFYBvU5hc3z/U9Yk0ZmAmFp90oP3ZsUunq3Wu
f+IpvygefEdgYRmGr4TeHMdMfUmJe1AyTyh5snG/wfrX3H7heuYoh5Un9/1Niwcx
2XMOlNYI4KgxkRfLiA166estEbeo+GjSWf0DLxqhP4MT7lF7tdi+iBhxrxCCGt7V
SJS+Ahs/jubsk05S7TXMbQAwsqYxdDlQYa92FWNVsFHzfTRAtdSMKLJ89y9FpN+B
34pCA7/O9CnLvpPilGsNbV11Wfus68pSD8K+E2jRx5XtVvpUiVky+vLHz5k36XeQ
Cjqazgwf2Kg+9zI7pWGP82mA70iseMsEc4BOhphRiqFveL0Q9OE0v+zELGfxiwQP
q7SNryVH/Rzrc4dG9m5FWRWXb+wlA+a5cDpFbJAue8QMDxi3uuRjeYGko0VV0t32
3b35PLoNgjy5zAWzgVr4q+1z6xgm6J5NWg3EoUkmgegEhqVrpRGJwix3c3Vlmum8
Tc1ttHTpFSbMBtRLhv1vD3PR80m1tmHmZYcLIBEXLK4JR9dsKsgenulZ1oWQeIUN
+fmeV4m7x1ExRD6hriIooBRi9WEtWCuewfMnGj5PgH7NR0Zl4pU/vm2iEaylRyeI
lAKPrc8hr3duEqTDQRgtQO325Nx5gn70EF4Qt4lc+g/zZW9wyp09EcNQ1ZkePF9g
awFJMOYTrKVW5eB7hhUnfkH6ySgzCQ+z94leNW4epni3TZgRfGy9Eq/H7rblvL8e
B9LEL7+kUC0Pro9r5ZKhPCVtD8yW2rY9zVB0+o/npmmJ0JDGl0PszPtbyATbjbQ8
q4UD08p/zqQ9KKZ/HvAJklRvS/Vk7t0NfcTiCk9j53F1o2BCBsnHqn1i5ENSvXQM
tJPDcAarornsb3QHK/TDp5j76gc2sEtPCcxxeWSEyZCABDlQfssWR+a+srWPmxdr
96b8ya3sF0cz/MJ78ipXxu+78+U1R8AxczaoSB5PIjjV5iuewiXdyVeZ61KUdmS0
wuC+YaMh25K3vXBLsBPgUQiDU+UKcmKW5/TJBSJors9MpEvKc2tzYT3kQmlT3nIF
JVB1LUgDMCrngCtEG/vzQU2A1+us9Bh7RavuAfqj/nHQrNBJDaFolrgV9XpP7QOh
ipXZHR+zBmVIrh8czZhHdh+Lo9Q4B1Pt5A1p9gw0n1wKDjyPa30BSgNPbCAu8MSP
LXSC89+nNz1zx3C9idnw2anyq94w07W/+P/iChLian90R/L9+LQfFzC5oBAVnZyt
sntZHMaEeZI4n0m2YeGGW9jm41QgHfDjcwQ2ULtim71nUCP88f0SFk+8I3BXuvnL
IZYSy7THQ8/emFsY3KHAw/hnBwqnWkGphHmvuWtdo6jcdK7Tx8ShWfbZLyhXYDac
GLyKgd8d8P+lsL+Uw0Yi+ZlC0vbmlAaGcUVTgCM45IfGZhiAQUExzUCTAETYyipQ
cjjD6Ybqn3QlHNpY/JyBiPnw/gbp4VEsDCAF4MlQYKnSODddc7+Q9pxCwjIM28aO
GFfP1RAOsgXjsjEM/m3Avqdqjlz4pCowIFDHtNBxPFetiHLHP0po38HCVXn0hFcB
w0ZEi3WSa51LFXvESh99D6UoJtBZgMUAmO1ZwmCk8wHK3xWK8TZERgANaZan3OvM
6Q5AoTA2PajPjxviMs7c0fgqLCDDQpGB4Ciadh4VHoIGk5B0yy5jkNpmNIOP0efF
IjeqNL0yEbh7G0wjWNR73SZ7g/H5Avb9uhwzyUr7oXULOourDYj7Fs48WeK0Z6TI
DRMbUpZ/QwsrEbLZBmRmAZwwi8Kpy2yXpyTqeaseL58fW9tvXBTZn8ub677U7JQK
7vzajiVhPH6KMl1E5OBRjKb4Dx8vdqOF+4fyQjvh3W1GFInhjqWShC4GkuUlEFMM
DbljEQWC0pljf3ceAf21MynWvfbtG6AB9IZz9WrH2k77CPb41RKSU4f5MHw3uzRr
fv1oaveoZRXfO9CxpUunIdLlhKti68aFE3224O4TwCGc3yhYJnLY/iPzzRUihuOE
jxhnL/jTs4JzwS0GAUSW9Jl3kC/o2Ouae2NLFQuUjtHgIlOtKiXvLi/TmJ2PHtpu
xYgcXA1YrGeQwUN9Dw34soiVs0ywmCIdJNVzlkwPcRHx+mPDfdFsGfSjo0peG66S
2LZpplNAo+tZ+tGcMNPYvwn1B5B0j3NfZyRC8d+VdnS1zbIzBBzP1xf2SG2UA2zM
hq4cBnVG1ViKZov89j85ylLWq2UTP22ABbZrCAyvECuDRaFk3xs9dhLzy9s8gwVB
xgRYhX45P+XxY8s5IlJgFw02SoLBOzliBdjFAzyPLaRfVfUH2w0QOWlmTkXJnyJ/
rBRO6gTgsBcbWeURBFBCUJXda7Mdoe6YaAjheTdDXP4gg/HqwPWYQQGg5iNnSN4E
UVEyQH26SFHWtNIP9oVPni26zxnBTLRXdzVya9fJXbidU5WPgrLnq6uIZj6FZegR
SQ4eVqv5WM7KaAWAt9SDCsgaTXcQaV5NqZFLvZOTticFuJdTMSrjkn/z1A9hV/+c
UC+btr8DsVVpGGmiBlSa4DD55qI1i77s22VijsrBQb7ABmLBtsCQZjQZqotrUMdR
inuE63HDDIwCaj9Bof3ryjt6RaZyxYm5N+QMCWfMTKoRvE5ytFQ+F+ueA43AyLMv
qtGRbvXh0i8lJ4W4MBKmS2HstCmR87PgNONHcCtHc8BaWMKarlKLYJVIPiUbwWJS
ISdjyVEn6Tsar6gk4LuUN4nf61BbVAf+IAduCPu/EZISV/TzTZ/ybQe/lzZwNkGC
m6/RF5OAYGjruk3EuqSNSLJ/BEeZzEis3R/35t+LNRt74NsUMWalOqLENNezM0ER
hgmDlZiwX9LFFy/lw6ECOreFV1JTBw8mpl7W3y4Qjdkiliq7TuNsMW/KMyNgvXTa
TfQiJXraVFVM5/HHsaxp9H/zQ8vCSj5O2+SvOl06z6hhe5i06y/Lhqa2+MaDJzng
u26LyjZ25e1M3kuF8yLy/xdTRCiNM9G0F8PrK6aqxlcS/7T+nCGGAG09mhZ8WAmz
INuhazLBtWb9y05GZpgCNB18l5hl1nDefVNQ5YTweEcfysmTzfhoIvHh33L2bz7C
VFS5CM4XvyH/WflM4OlYjZTvhzV5xP+obu1frhdRtYQT9Ur2SeZ07Q+55HGyzYfm
MjdS/BMeVW209a7LJqHJ/bstTMaQvJWV/S/p9vUMYnD9s16aEUey6nusEiDhkOdB
ihNyDEVhOjvhMf1Mki+QuOiUDAuaJ7Phv4wbTb2hirB4BzSecFfylLv3uHO8Zjaw
UE/nd5w1KPGJZ0JJcqv6Nj5ZctwDHl810hxY4u606u81LLFegi1GJQOBuG00cOFW
hVo6uJBjHiOVa3gJaxKF82dboRjGBjaal+Z090BkEKaecPxnisLnKMFntXWcpB/H
/9LoxRea9YuhVSfpJ9vf0q+i1Kzd+VA2DcozPKTjiIFgQq3uC9tqJkgWUDhXuHmB
sOJBTpF8FmuPNsBWlIT1txLLTCwv34baobryDSzNfpW+EeGkGP2I9oHYBF1Pq7X+
Q6GiW5kxlqf2vfphhVIZQUmFr9tDB4LMHNRXg+bWZ12/Yqlc9aNp6FLLsoC0lKvm
eyWKS0bJ8QkE5KHqLxFFZv50W0DBciowYgtlVG68t4VA3c1sUsHBNSEBma/yxPgo
aUCJy35FdnJpp1XnN0aEekR7+HD7efggGjrkSFFVOkn+23rVMKM7PJ83tF6p/4MZ
elZ+hEfvgrTGp8VJZub7oGilGUEpr3+33J3p1F315T6c1vDy9pW0zLNwREW97XLV
hB1MSOTOSth6Di9GZRCC4w8oOuFHHF20Gpwv6f2d9dWn/6nUwu7bjnaItpbOr6hx
41i7Cr/WG0gyV6pXGeIFQFehLIabXeTcb+5gRgmbyidAS9M9G6ABEb464TvU60yx
ULK95WRse85K9iwxYaTplNi+5scC3PMdMK73xhu5x4mOHN2zYrWHyXnrTtEiBbc1
Dwo+7sPN+6+WEsnMMAR73ZwY10FMJkRNhsBVnp9u9rTfWLEEQPMOehtT5s4I5yBf
OI6Ctgk9uqFI3COvWT7uhsI8r0mU/ylcoPlQ/sI7JdptCe0Igz9/uRVo5bjwNfqV
9Cuf0Hd0y9XW8LQfHvFf//dqZLpiLkQXdlyUuLHYRy8ZVJXoVrdT9Ri2PcCngCxN
Ed2yeKDi0LK6M96rJ0dMOxIcymXUXv4zPXglxYvb6BaHEB+L67dA67zq2uiE15y6
zoYLNDV0/JkjSMsGQdOgSaYDL6ljClx78eE71fSVzMbesO2ZhAzJa9Of2KTOgX1L
/35cPSbjzHOl2twP2fVTlolEVx8rNBIOPMlWfe0nRHSsECY/qmt8FCrGphdEIjsF
l0jeBfEKceX9mePDFu6gWNShpFnRKY2eucEmYRG9PZemMd0AsevDvevz3gUd//Vq
AyY+DwqDgLM7Xxhho47FFbdagXsH6N+BcUhlqffPyNvhJkm+uhZiPtaC7jbpoFYH
8kjYJI8mnSGxPjuFomOeyVf30cOaZmctfJhbObl3tmm9ta/bXvlSBGAcoD6AVPUJ
rrD0sc/Y8rJmBq8sEhqweiw3kPOheMfVYucVBHf7XGmWM/1cWfxpyA+IMjpg1TD9
iAx5QA9CJpxUQivQrVFPWAhQ83dEaHwW/0ku0FfqS0TxOTAh8uwQkBnYqeHWiz4H
h85E1Uxzfclb/01iPuBHxyl5YWmYAJgEXWox9pu1i5GNShZCN3m3ki7QmWKE8jq5
3Kjor5z8K6McbX0Ir+t/eukCmQO4gm/wDV79KbgqZZdfG50aOp4JzSJuh4DCNKhH
fXI6NFjlKfsQBX+RmwaLEzBTVNFSr9jHziYGRoc1RkuLAkQRYdcTtkeVQKHLBblf
VZxMDPHbG52T7dSw6RPU0zx2BuJ3GapoZu2RRDI6dq8HXJetcZ16cxV5DtoCltx1
97+tSU1uFuHBISYJdkyPVUfyDT413+Z4lHyzcNrGkBFs7z0kgI6BoiOxmUvIf6k9
s4C/wP6IQoTGPse1xlPDB4m+8aRbWkaTSnqKk049BUSjVYxh/Y5Tm6P6TnZKssGr
fDiUHMosrasnbLPE23BuL1QxRR5pj6zRvDfRSVF4aQmJIHzmFisc3J4x11vsRhmD
e6BzgKUSury2kTdGo5stdLYu5MilieDxH7g9Bx8HTBawl+USKXxCMazUqbVVnT41
LW9VcNQvq1aRGxV/oKYyp0wrAlcyUhskEHI3o+0te75Woz3aTxeFvtLBF0InJSnc
HZ27pp/VrQmt0DlvGPfqiShs1XBHxpqIjpCsqsVxnJda/CANUclP9oe2fv2w9hgQ
IxgQMleaqIuC77Yv2U6D/xiBaObSlTSrwBPu2Owg9NUKsN8yhUGKtZa2azd18Pd2
gSWca7pF5KjbF52wbbzQ2d2EU0OgzKlyYb6huPzTFZR75PONuIAVT1H8xrvaL9pe
NRDapk2dXmdgFAnguELwPdGL6hHLkIznQu8bw6Nab45PiTpvPOELiSUDLXt8HuR3
6PSiaRQRccvJ44pJtayL6JKt7FrBbag5bRKmMcoEs1zDse1dmsqKXgp7iCcdYavc
q6yaQ+G6rsPeq+v0tdYM5mfBGmeJUWVV678jyDjANkm3RaiZscrgpMy2RUTY6uHQ
ZCBSROcq4zhMBoIByuecBdPC2IRxcwZAGzUy22eJM8MHCUtnpWdbCIHCel/w7hYi
Tpq2nmuFBUYEBU5gNQd31YzsSuLuHYqYixAOWyH0/Op7RmH3iOw7r7YpnXOv/BAU
qdmyM/b9rX4O9ldpqc1Ydw5rqur6er1KvfU620Mw4y0jEXv4KdfZ6A19cJTdlsn/
U9ifnhm5wk4t6ypPzaObcv4Yh5aJhyLdmf+YK8Xh8O8eXRbQv3uT181HSCfuCKmZ
0mrUcmt9tLAnMhtfccu1cM29HbS4KD3i0W2/N4nYlghiPMTV1CifFwKh0iwUJw+R
TswC0gHKHPnTlyvH4UFErirrdqH4B6BkHKpGqa7iWAgG+v0neEP8C+O4yRjt/ogd
6yNYx2vNWppdv0I+ixslOjfh7GINco4qaiGOSeORsUL2+Ovs2127KFpHTAoBmyJc
iFzUGk+ynbA5FWH9JaqDhwK7UKHBt27u6MNCh8rHdDvig0LNvIcldjInv4R/1417
2NqTxVjqu/YBrAgB6hh3fNLr9/RRE11Q78zuy8TzPE6jf5n8Bk/sBqzmWcAgeO8J
cBTC3L+7LZG//pBWGvPmv2XFWNocYugF2Q/UgtSlSzp74BSI9UeuzDvm5aTVR6gO
8ADJsjW8Eo3Fd3z9C2FN8ADrZ8h0GaLV+lzAKZm7CZIsZH8/MysHiJqi7jRhstzn
t/77a0sYG4olU1lJCvjeC15gy7hpQ7DE2CZWl9CMeswa536c4hAwnNWufe9Bb5Ys
khIRiu36vT0leSu4pMI8bCRyoNMnxu2JGsFpS0M5QFhz61ACMTlGwL8ej58e8NLF
eHOxtuvckgUnOIM6E7j53UiiHqWOHMQQTp6cKhmTN+Rm8bwn/Z/h8nc24xhoai6b
SbZEoiAsADrK3nRutvLMv27ZXU2Qcc0PyyyRGNUdD/gjTucRWojvk1WRGF99pTmE
JgLRcaUn0+P+8Du7biFcpLEXT73VSvj5Q5LtvTOCH1s1GIfA1cgUdWUnRiN+JAH9
SR80hEIUEm/ZOq7AL7OF1dm37SZXH2gYDuaXxDdIx+2mFRysVmfujgTZWs+93Opy
qXGt7OjRCopCz1oPKK4wg2ucJI+ycInzPUKChWZfDqM6nwhAEH/YmSGYLtty5iGm
ZUAchEWUEe+uroRj6v7oGh5UAGACewZ2/MVzsbrP5f5+mQguGlVKHpirojsKeDgv
LwdA+lPL+xvPVS7uUVgZ0u0bvgOZPNSKzKiOyzUc8Ft5tixY5/gFiW7km/ayYvhS
dmLRevkcynk+b+7mJneI+EhpUlCsc/ll/2lkxMXPLu3vtnyf6qbokeD7hELuRBKb
TTsMDDuPMZS+QOmF4bwefRAzfp90N1Hqm/3rKoYJZAg4GfEZq3e4LpBQDau4+Hh4
H8rkVemNk4nEyBeALY9RHBQH6qKJHulv7SpgeAqDxdTS17lKcmejjmTwtEWTHjUt
+UHxD0zpKWZ/074+io18drEmcIStrny/ahzJQNv7xVIlwHcfJV4b7JHb3Ckwo1+r
Ub0RRp/xB9cFqdCog+GfjCoemlyPBFO0Q8ekaB+nu1/M62ijghZiBAYLIlC4mUE2
eZAqMJEOyZ/4N305HWYv+Q/0sjv+VS6W9AtvhEDfYYLnjFa+3+NHNbYHdr0JPYxd
iqsvcQ8al/w6moDjuIagLR5XnYom2xOHYtVCJB1fatMIyu/od5eblACcaCFCiPYV
0UNuX9NPDeTxMuhKHU6Si3Rs7MCzbH8qVkFaEZkf92kFUN+gm+Wo+UAYqdR2944t
SBd24e6+sSoS0CFXSw9nQMnWhCQb9U38ktBboFFhJb9NmZu8N/2/q0SWdmArs2CV
PoO4IEbYz+Y9lnVuz8TWJlzbJS5ApMKb12FVPRqZf55HbFIwyYmFtSGXsfVts841
GHDxPvu6E//x55pNxXaKLCmajYW6xeSMRJ+VDVjQ6nlkrXfz7H5TDk70uu3kILJt
pdwNemuoW3s+inkM60RlllMdEz5Fm0Wb7Y5wLa5lLUebM8b8oGThGr0X6pkdS2aY
YHVEsjJshwc5HieSPl65besbPjb7u48tD9CglWCIJRVcMZTzDB7Puqq8KBPRMQhb
Ta77lODfQD797LPv9+0ku7PG6TJ8wzUaMs2a31pARg1SDui31bGw7uo+XK2ETWkF
4xURZuOjJyMq5g7BJ6ouOW0r4yIxmZPQpf35zaZ2RKZUcyT7n1OZYnoxHWKusLud
LTu4zxVL6WvDGMB+Tl4oojBwkURPq4bdPDwmYc9jSTwDMc2gn11hj80uDeL+jPQ2
wBMFyGrV342mQsv2m0fPNdBNUm5fJ5CNmMo8CvHlqI7oftmpCdg9RUgDAQnkbW/V
JVcCKetutw3TZ34dRgSm/aoqrSYalRJTA/ZitgXdzoWW0QGsaoYCVq1TjaQi6MVz
ftHHIXTu+/O16WXxAoPksv59IKdI0dxQvSL19hfUn+thBfaCSFLCf8j6UFRqkucd
+95vIKoBhCaP6vL5bqPdF1uw0MGlsVeCjM1XdU6XUTUbNYiaV+iUWUoSaguJeaE9
vlHwkrP4/rJHaM+WzFbQJJRULHGgO5A2sIuJ/vT54dEKLa0sNpO+cULx2a8j3Q8C
B8fVUuBsbKi5MNYIckwNWomUPCQGI5hdvz/UVIpTeZalMcB/hgU4FaxPmvtj0bdv
zqKMwcdHs2RnGNjmSwFWiMR8aI1at0Z2qS3I7yzZsYZ1HRcXRujBc2c4yoxDml9t
4i05sDMaOMGrSIEfUW65LyywnUhgEkaHis+9+DwBPjynL+i17LSWoLPy8sK+WaxN
h2pE+CI5AFSLwtcZGM1vh+YW5mCzS4QWAL40T0Um/tfY9HJ/W2faxfdz16Y28KiI
d2fdb5Hn8GEp6FiCAaOFre5v2rpeZ77A5z6L43+AUC93YmE/g1AXTMRObQckgs5t
IGedxLFmK7OkE8BIv/2uv3rdO1Q4BXk5gnmvceMVhz5U+atzXZNrlWpywtOxOVbi
5vK/cJSLsa8dWlzCVHpxDUdi2+byuX+ovFh+jIQsjuRgljjlL6ydFxPXs7Vv2Mnj
Yeh6MaxGlql1mkHXK+dCo/DLT4hMT/CSMpouEU7/gvdLSlcSLY7uYyH1HUYE1zTC
QXQiVWkEjF2dydAVjY4s0yjVZdxUT5crs5W4x3qNsT29rrmFXUbpfSZOHZG1MIsf
ffAgBxS6LSbl5oVjHQumiXl8juGylZUitpYgvv63zUvYpVnotZaIipyunEagPj5r
ErERvTK1Og+VfmASSpPrDzDzUplIId+qRvRwgyhCQJhg2iJg4UQ+DQqjtAAtjHTo
hvzDG4ZdDjJiVrn2B3fVliHYDNWave7PeappINLwhmbOBI9PaRHZ7IZDUajygYyr
knz/fjONJeWOZJiiAJX/TknCK8hUsM8128WaPnERAylksij48nxcShHfwtqtPNX7
o2U1m64xa8lOE9BCLn0Zd8+vn4rw1BaB+qlg38mxIvhPrtGCixAAzO0DEAgTXk1m
RNk4I0PUM3ipkVugGjEn3mJrZp9CK2BvdzWBXwD0rOB4JpEDU0dtsBXcfbxmgrUj
IpGr7k5iQigB4ItVYANnsOUFLR2Q0XeC3hti3reYL0XaMTbiWMFwSfeU8b6e0z99
B0Hm9d8aBSaNlMvSmGHc/8XuQTcHAEO+druiPxWhpXWqqO0Gt/PlOVwzWhzjZ3B0
mrT6vyNIXFYsfPL76nKOiNql63tiM7+PYupFO3olTshau0zPQS133UwJnyYRR+k4
xPsfDkuB5yBHR/eo2IcDn2vQ5D5KdDr0tNdHns30ekb34AiNr2gBv/p9yrGcLWaS
cRZd2ExorAcXKZiWyFZSXuBxUsEBSCOS7/U/4Odcnim2he3dpgGkrTGj/Rg3Xul8
A7NQhPUH8Hw3KnBm52Elhq6t/4nCBGrJ8d091OSjTMKEF8XbbMhLUi9/5QqcX7aj
htcqLwTFCP+FiTfBeAlBApTeHK49F1dX54ZuZMTf29+8erX2rLfjfS5lK+5AWImi
2jpPoaUHNFSiuzeBbluXjiLb0XIZffGMU3DqUUJQcUih3TZ0yD4fsLRiCyBVui6r
Tr4UkOTqQ1QxZM1NYatsh+yFOci2JfXzR++a/C/8kkirmqfK+PUaygmsP+B8wU7E
As8llyNaLSqdmOOLQEPehZu2UTCq0YYu5wLzG/jronzfB1z0ritSFIdk3U3DzXgZ
+2zBVLDT1100rhITs/rQKfRa3+qiGj6ct1t1u9LxJTEgZgIK+MnKun3nTLVbNnC6
84B2lgxwomM+i3AU4ciA5/OEDuBhIChAHuogKxNErZxfIgpz1OjRSzE4USKwDK++
9qkq/koEatsAmjE2Y+L3kx69FlJbkREaiGZt54o5jBY1AnWdGqonI3YPKykIKs2r
iPJUrkaNd5F1XYGbGxEXO5VpeUMJ5tlIz/fv2cXF1kjU/mPkZqxV16aUlICziLXP
B3IoKTDstybVIdBkvU1aX+cn22rLC8MYpvgoRgw743vZSNK/9/NaUuiw5Gi1n2Ch
8GhaPqUKtydQEqTOLT0sZVQCFhvpVniUQCRJuQfsFs2pG/zNjJO6WJmwRWnUbIw5
uCw9ftnPd97tBWKYvyE4Q20jQw2teN9IrheojbkFVUy+lFe5QqEI2ywXdh+yGEe4
fsRty3qKYFuuw0zlq4yyZKzWCUpljDkjnuJDSO8X7gvzSnUgayr6YnCbm8jC978a
mlsd0Dx6aieWJrr3Sqd/iCGwOmBJ6aKeoY3dsfT/F2fEhf9hJKeCjkp9hyxT7yqg
RqXOxybMdtsOzgZf5GJTpmNOS9oA650fAKDhEaRgEF6LAY7b9XsDIEDODVdl13cW
jaBw6b3WQTaOhDb3J5fSD5/Y/ArXSB8PTmUEWIplFnDLE0cAd5oXKqYLF4D21ek2
K1Smp/B7UoUUpQsoxixGLRjpU9kvuFr6BcjGnMWaPl6lS3h7IpeJoMDE6r444ySq
J6frcuInsVGbdXEbUuHl2B//WdHHQREKhni4HbYwGOtDfR4aHWP7+toX2DVU4MeU
M1TWPQ00XBUVD0b19+bUfcY8FSKjRpuABuw/3bkmQ2Wcbpdqn4yG8KOtpJHZ3TM8
b3HMFziSgwHvmaLbNCFYp/PdRyWrz4y2GwTDfEX6v6vN4sDRHAhn7pesQ2DXpkSI
7uDyiK5vB1ubPsNjaMUJN1SPUIf2W/GbGSXZnSqgACwU0Yui9nvLWH1ak+dTYBPr
hWNy5J1MqYdurFJPL4FA9q0YX7PcLv2G0Jye4va5jEzE2z3MtpcXANRZcqIYTweu
Yt3ey2fXw/SDR3jU6JfDsVh0FYqKX6CDy8CF1y1ynJadPRQ28pYnbTZ8mjvlb1KO
stjUaaf2g4o46esF97mWzm0sd6q7dbYAeTDxkJLkn08+/8NI2JpLkQFn2LzAsJ7h
8fKr8xRspQ4paIl5ntdAaLpJdOFjvJtCqgIVemIUlExD/s6W2twi3A8u2C3lmN+F
o8wMKP6jP7ta8kFb+IOYl0YFYB5ZcJ/RLtk4MmwLW2l42NwzK5haTK5IT5oueJVL
L8GKAHV6izXpp5PHphhWpRwB5IbYfQx5W9c3kYGQQFIbccGMcZ3bTlsz6es8jLrt
w+O8CtiIco84Z74U7MRsMg1Htzg49Ydnq4UJnArx0XdlTN/+ZerFAGpbWSJYMiLf
1vaXEXTEUnN8a5wqgTHMLkHszTkjrNvWYfw83fiDpblfRtsUjPWQt809PjlWO7m4
8LTbBOd5f5+fLdskb/7h2/UXJmQQTe96ukEqv+YsUQJWJVLqbF7ceXeVj1Ujf6+S
2A8Txz0p4rruieHUKCtuFZB+48A8uWbPukLX7ZLG7dgXbZE1t/hipRDvENMUia0S
4yur7+tME7Lokw7CuIrPVKiF6H2Q7pjuoNUmfTk9Q/BmTRP6mL3fsGEvL5Yjn1wI
JDIqUnzJtv4kC0fvpN1rC+zfLEoV3zKBciBRP5dgzWKyF5VfmzajjiRHQfZcgCyR
b+eU/xQaqvHQtZSVdAr+3VGfNvyjj3V9qH6HMQGFN9YrmjE66nVcJ3X38arF/koV
CvC/5ARm9gsjX13rWY9AK5YZBTEb1s3ewJr8tFaZCT3j8HH3ElT6q0O8O1Z1OVAP
baMdft3AdC7x4CuoFHwMfmpV+U+MHztSuMgcjF6+DYs09lNQjW0gjIMlZW9+Gjjn
NQnZPNmQZtil5lCou3bEcSR1LNYwihJ97QsDpLhDoLPCnS+qpsrZsXEYepbIyhDN
hsO1L/hg2n7fZN1FU1iLp+HS5sbKHXwEHdNuGz6iuZ6Y4ciDmin2Jcw/n1uhuY8z
7v5yX/BT3I/bL2xUUVXpK7DXxnp5T0ugawufLftZDV6Xgcz1GxkETCwA+dPmqCUu
jpI+uZdOFZsWTy6+sfgTuRMnl4YQtaQpGRgxPQuK4gW5DqbDJb4Y/uE2ibV8YA3d
AUGcUKpES5PxQ/YSiwom9RyFBWIIHmZ/iW/o3/es/xEBSUAPEhs7KPFHavsH3sEp
gzawXNg7TIiO3J5IgyRuzO18GOgbmbbqpieHxr1sQAWsmWjPjaHq+1bHawjTRWnl
3lKN4t3g/+zBuJACVFTBwu7flqBwIj9WG7JN4h3RBLP/YNzblBOtzP18R2jluEn2
6KXPhNnOB2Xa+F8G84IRRMKYQxQJTH5DlSjW0zJhefKe7raGEwOOdXtWIShIw3gH
5p8My6DT7a8ToT2ILELxJtpnO2NRqj4KUgStqu1hngtjIqYWV4Siac17jERIygfj
hHqJKjO+LslKelUQTAWAA5f931qGpWUd3iIPEIWAG4CJ6AdGtXkbUWSyCYyjL2J4
Ah+dYx5DVQIrqD85TL3IoQWWegZzq8tUq8T+ZhbXxUAg9bIg0FoNAlaFu2AsWJ/P
XTRpujM6Mc5r8LOVfGCw1QF9cWAmGhL7fptU0dAOTH4B6euhSXyUdopYK6JyXJxq
+K7ZQf0iF5WpwcSiukDcNj9eW8DfyyYCz5XcNcA9QbQ+JhpDCAssQvEnE6U8yHjm
BWO8Qg0SMcTzeMYGtPxoQ4vS+n/RB7OSywlWV9fakQ1LBcn+UNtn9jWEV5prOJ4n
AbZ8XW5/jpRRSeZAi7+YUcDKIpKaMq6c1v5MTs5GK3gkfVPUg+k7KMcPpN9+9eDF
9RumroPMeHdvyeLYVmESMXHRwXXNraicmAQx3CgGZMy6VHk4yzIrJZSn6t4F/wSU
1DsZNZxw16hZkqghfHGIinMAYBjS6TmeJAk7xrRp7RRgy7UXuwHo1wxU9cATTj2t
An0J4xa4rlHZ0f2WUyUCOp/V8FYKhbE/Km4Pa1zyaAmD1XJ8BnCVswPCR1CervkD
Jf+NzDcxa2Yx5NIbkRKknlNtgRocJp8Ld+YaXaoCBhG5Tg0kfO/ihBrtKGNDYTRZ
RC8zbG1Y/z561iYafGhfJ1FVrHp8mgEzzywqa2lYA42PcVYhDftKi6L6UXpV+8T/
jNCnMBR2YZ6i2JCRWp4mheQBokXsavlJwFpjz0On5CfoZiEgb40Yi5c+uIeaxH17
uISNseGT7snfyWRT4KxfgSaVhAkZrv0wY9Ay/GFGSUkkCXl7+ToTINBdcbqYpdQD
XL1nYONE7W4qiqTVp1cWEaFB5LDWKhW496tFgtEMDv9q7Aru4D2rVi93ct+mp+UL
Cj6hiL8yaZxnwgx9FAD5NNDtfiJXUsQtXi5+biuia5CR4TGXI3cZzGmenmWWmhKj
5zQYuixhz2Zvyp6iAa0wzwVwYR8s/9d6qDZZnlpWDOH/QbfCpjQ5Vr/MAJJls79H
D/68sFmN2TkMsRt7lWxo3AFMHhgoG2zn0yTmkamQle6A0H0GLs0hnwwG6zxClmQz
4OUkzcRgzi8qvshvVLgKEza5auhDCEtKcDDoBqo1bKBhk0htKJ6rQLGBOLKvk0Ns
RkE2MnJk56mcW1g0xf8R3mbG02OHQGlHtOjQt1sl1uAoCkjMlfGiNdr823PUJi71
/Y/UVNPlMfQrMFdPAcitbQgNTlEDU5StlRz4fPG0u3bEnyFMCvnftNJEd4QJf8D3
4jiudFPVQRxfRYCD0m3sO5ekFV2qPcjx8FibFJDx3V6+ASulHho6GFjoZknY958w
kLoI4HRDFyRP+hk0Cuq9Vl1rvPLYiRcqMaljeoqlwUl9nXKEiZMZnEUCuGoDVp7E
zCoVp16YpGtq646TtS9nNJk5bJpDQcURQd+wcdkr3GGmFBSPm8BpHA2A7tbgESsw
qg5aS2h4L0lDvjfYtqHPFaMA1Wq0jb9+LYmdKs0w5sj4A8LMy2opSOmYNvgR9ZVp
haSOfN5lUh//ZobYQtNvKWBy4ggFhxx6+0hvEpn1CWdR48YIXiv21kKxHPlLSgOm
lp5amYltOldEAJEgV3Qm0aKYu0RgvWNcBlYl6hJPvUTTTZvic41L/+vUNabvMfRT
b6bzwkXY/CoLKAOCUB8K1viYeKMFPo6TS1Hx022c53/VfWCEZS81YVpH8EDSuZFk
MBsrNK6DMK1pQEU1Eh9cA9mVKNBrMzAiLECyEntdFzFQAhRVY8WsCppPTIsEVAJt
BQ+Jv1xibxUcOQRN5qroxKgY27INA0tu2vae1e1dLzbw6zkomqCxYpVrWr3j+HZq
V487UTUDf3r9t5UmcmclKEpye62FiQn2cd60U6A943jPooCw7khzMY3/y30Tni5B
gP05SQP8GXvIF0xx1iO6t1AXpcHuoBqy99j6co06qT76+Pu5z6nXCCZ0m8tUS3sU
w3D54swrQVoF1qjdr8S7ZbcUCBdb8cqkHo/bu1xj46AfgxFkLHHQ3H+A4gcJMoBb
7RNx1U8w9CgtuwYCrfC/ZFuzPwWw2LIdVe5cn1SJkgn4NF8vG3SSfsrf8fKpq+8m
DXzKFWX6MUgMsHjoIXbr90F5yqb1WR949oshrAaTB0BskJ3lbTuEGFv7EXUemIBY
NbDUwB7ExDEU9poR9jPyL9WdpVKE5LubMs6RfI8omtgbXMVdspqtpETbYmG9H/Gg
APeH05jAB2YKTLltWfzb4Yo0QTfd1D+T9+aINDL7RBj+jVoD6Um5rcRqIRur9O1d
Ein6EZCdk/e+9z6UBW+LscuuOg1MiT2IkoCqOs4pZX0/LNaMNKh97kQrvfeTcQLK
rVV+tqo3Ge+G1GKe3Ixp04jE+tFc3lHphV2wAefrCu+KrgzC3KEmodQScAFP8m4t
AuGMpIcBnTkDgG/WB/m4c+eQ+nryvc21ROeoFkTc8WgLNpbvC2ar6WNcznbTxzLi
sjb9tzo/2SSguTyjMQCtr8KgjpoZcG9+bCktJJWR3y4SnxD0BGKGVx/RBsOSwYl5
e2Iur600nqCRlnFBdCxzkgWUSPEIz8s01Xf6ep0Ouyp25iyqrYHxlkekXJ7S4gK0
I+5GHqbCL8ILZF2c/THISWhGZHQM/uOHJxMEs3cJOyKxT/vuEEgkyrjfF1+ZEyOM
RH/k+m1x7T+IhrDvO0KGxKfVefOTQxxKSxx9pe4Gw8JUFkNiAfg/e3c0ZdnLGcc/
6HB25W5R5LVn00PwToM5tfpY2B5ypzpJ6X57jlfIOPbCHeI3RgO5QX2NCtQvo9pi
eH7QzwJ28TSUdorbH37zJwczcEOHXJMJt6wthW/gWqJqoOVmmUbTCpyaWrtVQfaL
9J3c8jIAhE5AAiuNE0+17VnWFl6g+EPbOxH9OmeunXiQPf9XU/2MvTD2DFlo2DwQ
5eKxP/d3BjoYtednNVwFAvTtpVlgwrVJKTJEgDB9vrECB/nkXGg9XL4Iv0kF8f62
HkMfvx5yTkaOHewrDV2KpYv2eJTX6D19SUckvkuNIVfnLNcL0h64r99fQcdp+7eX
wHSNwJq+f2TJOkY2yPzQ1AVqdQ7fTQwWloL15aWBl6zhj4ZIVXMsXmo9tCagfQd5
B9MRvlbIV+oYi4ELxcx6/EluLyLkc41muz4HgRMlQOWsXrz9kjquyG5KtJ3y5cfe
NlMu1ZL1N7V0wxGvTCo3jAYQ0NLxDJkMANXnO9ItADc4A3qV5E2HBm0IwSljr+DT
CPu4XXyyP87ul+Rf9NUM8wwYZGpk8lolWBNIqJgSKlggjhZJnSRpHqNzeMzHmOKG
47tnuB+jl9SejSqmkuEOmS4JfH4zPHulho3tICURr6MsKaZS02PZxGNNx+gp0JuO
epkPhn3nUdkQl7AmwUSOTf8zt828DlQSnQw/LFSKDgg8NbjpzbOwKB7c4lloCTOc
/ZgJoGbCJ9uUf/RdG9/2w8MsejZ9SZDiQkZ6sA2s5VP7697+Y9IGN1l4YTNzNB33
fCW558twmfeEHMiIUxkkHl7n0YFXSnN6592xILTzRyvgpTKhWJlRPdYi4xfvQInE
G69sl5Q/vnmjS/m8X/99d6DpcmSdM4rEtPohfyT8CSZ7LsRDZVfs1QAiOeG7qe4j
A2Rus8MiN3jfIBTYWe8C63LxmWmzxjWMMV/2Imf8/CjtfvAzi8sBoaMxqKT+dvSn
gBEDL0SSwiOfyt0WcYvQizhOro8pCcvN/01xAUN52dI3/Xy90x8aRmZ5bOogNUYp
PX1V88FHl0R66nY4D6cn4lvNUvhUfl2C4PPa6G5a0d8BSDjiHKy/ZxAkvMo3D7QX
Kqxgm87QGfP1H57PcqsOIzw6/pkYrDADHY72CkH9B+uFgbtm7CPuX1GNwKH41p+Y
6ZYCt0z4LnkdLS1mzqx8v4wuzk6GR0QaqCQZFopMTfVptW9C+keQAlVO4r5t+ugJ
/KUZKDRyjORJ+ghUqkvScwDb1E0VfHfVLKRR1a9K4J22CEpeaTIoLxpG+oIWXZlo
9OFZYoTpxOA8wsuRBgVxV6RQhQzQWOjosmy+F61LQFkqE/obzoz9s/cPk+i8V5uk
ScPHF5UKh1SbALc9x/bu1siAGhUWqDWJC8xtStSbJ6wVKpTEUATjfnd0EtqCmyM7
69WWj+hYUns+K7SwOkZIeZtRvQkWjwBfc8W0OdpJBRfQvJZaeMqb8I/xxDP4ms3X
3PaJEiHG2zjq5h+7+31eHSAhvl4VeAlET81zBYY7vYIRjyaaKvGcDfvuuYHB+qLx
JjTlrH+5i5q1LVBXmIq6ihNAXYqm7aki6qAIq5fwRwLK+1V1Z1cRF+0/3dPu7O5y
DVSCgh/PPs8TKKyJlmEPtNs6PsZrrao7E0iSZoHt0luDZUXueutS8YN5+1AYHGpI
5/zwKoIlauFoh5ybT+WVIQ6kbWvWF5ojCEIoUdHoImMhTT/ClAhRcZ0EZERZv6W6
CthqoDbj1jxlnsuyjfyKqN3jYTwy+JpApgnl/cMueos1LIh7qG/kK9zhQlGv7uc/
V2LgY4Q5H7vpSofCKBthWtzRnvffgLpymrho9L7OacfhwuL1/WALQTheMVRHBhJD
EX/42HXD6IkSdAUuUzzZkxECTNVobLP6N7e+s1IaKdS8v0n8FPjo6Dos+lD3UMdD
9SOuIcAcNXTLVUb+crYUALAJOLemrk5FRbsgIpW+1LegvXBREmnnDu1F31MS2Tp9
1ICirujnghsLZQqVsbDv3LVwqliaqiX/DINyDg3t7cWdtMHT9gau1oBkX8dKOEo/
/XDoNNJAja2rowquTgPiUkPDJjUMrkhaQfVD7iSi04aSmUcmmHr8xyuaPj6esdVh
BgWkuyOgX7mLeoQtatX2JdluPX/BmrCLtfnczje7cHAnfCXw1N6LrYTVJ8AGGX+Q
oxU30kH3mYWa8HtAXeWpPhNoGemvIMcVKSMyygCJlSMYDqvysW+JY6t7tktFAmI5
DVnaT+XSumPshYuEzXhFozGpuFthDnMG/StcM+7Uo00ik38cZf5wO8kytE69QdM9
XiQTpxlpEaTmyGlQxH8s4PeEfxBLGO7kAaICSvR0Lh+MUlF5YFcJJRXwWsjY23qe
WrnBK4JbIx/C0DxGlB66bLvWl3pXJ2lGT/NDs4ZytXZ+GwkCI8mPa6lyXmj8gzt+
d7oGDf13gxB25Lu2ehdfe29XgA9eATgcHaJzFBJiYBmlSmR13WvZyL8FrRFjp11b
fNE3j1BwyMz5+EHsxLK64vnnbq9EZiZH0IWbeN4SWo8to6OWvLj0QirJ5R/cb2x3
NJ2OfCDTSzkkxP+3lx72eTd8jigyv6at6lU4DblusocOzgJKCaWQ0yftNcXltm2F
v+I6rfVihgSLtcNDI78/NF99F+ZBnfhgrR9N2nzOMAA6wq3TCmGd/GLV7CDVOHnA
xJiVFkRxmjgxcoItOT1ZCgmn2bBq1dZNDsfwVpvufubX8M2rTDGkxNss+Wh7K66q
I30FdrLAAeBCiJdQqaQ1PnUg9l4jSjfGO2rRkYvGvJlrUAEVVNNeRk5jzYKEyvdg
iB9/bd2W7L2M96l8Ao9vCMkxRuHx0X6lZZg1zfBRp3mzbozAnJjDJLuoDD7aaZcS
/afzXt14dn0RsPbiUDFtvHXkBe+f9hrqoKsFbx+MjEWjesFmjZJLM/8pJw2C7RfL
1rR0xUtwMl8sXfyrEukdgnWC0oKFp2JRxKNbD3Qe0qC1slKCcXjFhOLTxNW2cRtb
4FH3auShW6XkNZ3TKKkSlOQHX79OqRRImst+sdu8WlkGBtIm8zdsC7Dn05QXUv0C
KkyOa5zgMs0SG2W4JiRXo0jvaKOlebsRl4z3ZmKT4MheFpvjZ2Y12sxRDngqpynN
GtEwsIeCAosQ5/5wic4FFdZu2yCvWmFPVFwY7zNfX5QusyC7hV1W3v3LcbMI+hPu
kSSVZKEtg7hlOhySaqjIQDtR7cILhlSP9rNoL79wIxFH/32u/brcA/Y3Sk6pRGmm
G1lFzGi3Sg2gHD+DMaIRjU2KBAV35ev9988Ud5nR2nbr6ZMSEZSqIz5j7QQcflhF
SxlDwmc8AsGezVSc+g+6DbFJIxtWEXDKH6eHl8/T/IZnjUoWnQNIPIbT+2SolEd3
Q3q1sCs9VutbPOJoJE4mrf4NdSiPMx8U98qikEoDG68/hRCKe1PRIji/q42Obige
zhsGzvvZbewAJu/VHCgk1i8uoNhcqaLByltLZzbHBUELvlMeadzh8fmzwqYU+bTx
Sb1oKupsBNYI4COlEHdP8VqfUYIj3iUc7aEimlYGi/mc1Mz3duzpxjOQFKUb0JT3
u+OwbEsHJstED3lvKi3QLSTdREygTFunWGU0vdDAKb0NpODFZ+BBxM4UOff1nuD2
o74KzWOEJLvRGXXAc3AqIs466BJ86Z8/JnF5KyQNk8ssFc4xPeyvk6pZKhzgTcav
5C+9kKsmAaZ39KBO6iWXMkvgCwcmE5s/suTZh7p39EcC0LXaHzPmA/05L+GblL4R
3Y+i0bhLAh5YTBNvfc0yDhoD8XK3rCGcD+yVO+PtWj/BSqq8GtBQc3UMAfsgG8NG
V1zCBc+qkUeFjqyBF9EGhZyGNAg0wRxQKHKXE/CMCvL2zsb+KyYHVMisrU89JcB0
lGyoqApZbIhu7clt5BvUraicsxYGAFtGceecG5bc+AZLfmV4azCjME0dyGMP305U
5n0pvEZslZmthbVDEbY3SjvnFl8tfvc8+hK+1PFkz2L9SKf3rZZtq+CRu2sgcLEK
4QltWw1uIsCw0QE77FDFI6rwZISAi53l+zF48FChkrpDUurRVqSWlh3ybrcim41T
zlh/gLTImJgqceYdPbYi3fv8MUBzgk4mHJRhDeIt8HXomA4l4B09PyQQ0k35porp
tkpiNUpg61w6rv2lHPETvvRSJqtOVSDwzZ4PJAzs6o0W8kBZJX/b5vV02n65j5on
Va+V0zXQ9F8SXFIAUCQd6D1qTDG67iGSrhE5IczJoqhvBHGktu0tMLyRloVOO2of
dwoqJasscSDglmmp33VtF5SMW4HT8uIkidOazgkSnKj9HKDv4Q5c3Z2SKbF0db1u
WXr+65O5sc7Hev8lN9fv32TJZmamFrFqsN/k0fK2BoVrpVAq+KetnJmHzd6TgTz/
Bi9R2uRJ2ALYlzwAszGjR3LH2AkrEwHSAjW4UEDuboLMJg+sDs7kTBUW0Vih51fp
0ckienwRcl9M/AgMs9z+iqpBaK97bT+hpWwYtWJig4u1dohCczTRIstIN7PFV0KW
POZWihZRIFE+yESsDaQCc6+ujrGNDzExjRqCXpSYqRCGm0lBTSG4x+ATs1lDFd7a
sWgcjG/UjFcLG9ou01JfBxg8993V124MVyvUYsvWDQz7Ji7GInOnr2BiIA6uxkce
mR/GuHJKH6GKqYbPoCzZqvrAGxHdsGKmw+wq/fsMXZIw4dnYvwF1WWFF9z5xRpYV
Z5IFHBtKsLp/CrQXVtP5cELt3iftIqomjUpNuXo7hHRwi47X+aW09O0kc7Po/JlW
4qd20Yxx0l1dtEbcR+TtTfz1Gqj5h6NWZ0p2zJbxBx9o8fUpGztRIElPNaWAqAvs
ID+H0z5IhDzl78RLer79iKkWVqrvVjGf2yY7iH3EDrf/VuaQc65jiAsuVYnwYb8L
N0LOA6jjz2ccUnP5zVzkDEaw02DBxm9kvdDBpYX+VSKDMVyg+x9Yx81QKyYxzVf0
nV0eiHPVOwc0tBOkd7YXrvQxDYtEF7x9ydmMjJpq18aXw5h93RIOxt18Ihe1+i3i
A4veePMlaexkFbXDPGC3Fd4s+fbf4BTkZm7AkZtDWF7+8NMkch2irAQdtGDJL0NM
uCaMWDh7KdRXUi3KViYDUSGyZkDsWHNuJ08IxziVU8WDQgHIRmEOY9/vpr3gpYhP
7t3WacANzoE7UJi5ox16S8Qt66We+hZP+cgFqa0szMbI/LgwYVuFIPqFu1CYiuxX
mVF2a8VCWDkKNkAJXfdNLGgFHT+t7kvNrdPlDLnl4KC46LU2Y1Nwq0S+BUDs9nUG
qfuUhl2C3a44AFSjrJZwBwIclpYIOR1K59ceQrE/g5+ZJhMxskNDENJoyE4JwBKF
yS/1mkVZj+I/AT+EWsJUyM5S817DCCBXIih4cMp7CLQAL3C2bIMv/8yj5lH+M203
9MMcfRh9XJOGanUlg6I72ve4TBzc0+0Ilcc6EQOqPxOFOzbpI0IwVfOONBKvyNg2
CfKJ2S9YdDn53wYzbfRBUzLkn9c4UbD81+kFGAavHyK3gtKWfPSResAb6GzlUHqU
ZIYIyPXcpqD0pDtF9dMlxPEQbBoq3KpnM400Sswbkvp8eEihXAJ6p0SqDLZPUKls
9CvRifRKo/1YOueTSPjyvTHO7wZiRqQUVvBAFvxicHa3xKledYjQQQk3AIiGRofn
APyGJ0Y6msEX6nMlHp8E1ry2wAKlNgTJorKZ8IBKceDhsKgq8mUolIz/9O5CiTTt
kzDTNf+AR03TKkImvttKYifm6jAHz+VXismPsx5CahrhmAO2J94sPMU0vA/jCppn
SCkoSqoXw81+J8auVS5XRGrgFNRil0yiU9pabNIEgEgZHM81ufAAdZtXXU7I2Mzy
FNsiWO3/3Y7u5tywyP/VzAboFrNgwgeesAmd6Ng5w1Zrr9d9el+r3ld05hkKXWaI
lwgABqO++YpLs0/IsyqpYu9gMme5DASomfcDwa867CmJVEEDmKO0Ya49bEhxkPLi
c1GmFw0q36/vWxjDH2L2KesS0FZyr7TEQjhvsIEb38MfS+CJMuUSyo/deu6VL2x3
e3VnB48MHtaUZM+y5PGmw517ucpV5wrqBOMJONOUAELilb9XuBt98+XfKyeqzmRl
a6YK/uxzYT3UY1szhv2QcclYyu+FSh+iG7lubNWml9Yu2aQv0m++mktogOEpjgCx
/6yJHuwVIi3ju+dMiIWss0PINaHP1CeYX58YM6afFWZnEIL9anjbK4/fVT7Ey4Zo
habgGyJ+MS4vE3/v/MYhrtfFqaS5cA3373GXYLVhMWn1xSa19NOoEh9HIvN0Siva
b8lKQzXDLoLqeGtQq+Jmcdnemi0d+1uMXrJTWgTO4BBGz+78QnFztePcrQv4hJ7q
Dw6HddBETJKzVpsdgWNxaTCzK5OU30A/RfXAziXl53Wb2Z/wPKROd92xRKmfjQpD
GnRYerC7DmRIvd9GLsr6e2prdAYKCPKSxtavgP7qL6gDwHHZfqYN1O4ncbMsRPh7
BlwZJo1DOnPFYiqVFCJsTBdFggepqAwseFfvjLFvTQqt91ykC9PUmds5WIWyBeL7
8IGExAvvft1KZDu1gyd7NnW7zAhX6LfM17cgnYxr6OyBpc7Fqlk2HF5zeOt/LSMr
jnlbm1uMIbvZx9AG+JMHR+FiTNuZZg6YcYQf0E6/uJ4/ekYDwbxJ+4JvMGcA+YCl
I3j5mOrLzxscVlaVkAugXBEf2NDY90CLAot5WXkNGpnV4F40szBABmOm5dIuVaoW
1czS4RLml0EJKhPA8nAb0fqHeC6srnb+eKGgpX+KBCZickQpAGpmW0mmI6CZwsIu
EHOUJy1ZrrrUpfwefkZdpj/6pKyeAGStE+0uzIp+UWJHIZ3VZKdxWe9gTQHAgRpk
sfgO0rW4vOI5BRFO0wBZdq7WCqT1Rot5Z/uPl9vsQZ567iK/xIPwxmZmA2uMO+iE
ITIV25Jx9i5mFHjA4PPD53iHBjl8bg5g1aouS856hH38uXgRL5dD5RM34FZlmznM
Iw4IUadfyPujM0E9qrR4ANwgI4Rq5IVVRzcP3bQ6a/cFjM7u8OzJuqL1GprCfQ4f
EtEOmBw1M8PNB8tfT5pyt0LkG/UqG5rdd+GyB96ubHmES0TQG5CnzTQLOhJ1eD3i
hk/nU1OJlwZ+T34khsDv7LLnNi+uPvXUUFLJm5h3ogmhIziuFLIbS7ucGhU4HViv
pHZqL1gjlOcULHHA1paftddJZLcgRNapL/XFtrBFLstOKR3utqFsAZhmg2Fvn2vq
fG3Nb3jeNwkKVBrMH4KzsHmzTAvk3rpi+cHsokNKWwXu01Ew8vi/pBzCvR7XwFxN
fBkxB0pk8G46VljLdxoMsI1GDRtGdhBKSOWhxcLiQSfftnLZUw6aYbuHmJXEOM4H
arIv475hgd2OmiLS/OM2qy748CNI8qYUkexxoZ209FikfUEnqvsLL46wTEahfMtE
GNJwO+BOqMSyqe2+bjfqpM/7Nr0JUCBbJUCWMcsxWgiptOkuydv1PEqWjFRdZ+Gx
B9b5Y8/FaGHh52LQXt+TeQkL26c3u1GlKQKg3a4+0N2xAeG5FYHX0ozZsoyeeM1F
FWrjkijkMsbG8ePXnCAsacqhQhBpWfAxpfW7k6eLKQ1ve2tekkJiPIeu+RcUw9wF
grQ0zdXUXB48u7qlLrmjoyTLBlCVngVv5O4lCtt97y1cSBS6GyN4DOiXXuuH0xC6
D0c0FBfLUUsz3gu2pkNOdMaO4hW8XrPBDcnU1JYEITE5QGTLkg0xgf765SpMbItc
3M/uAQTnMP3Twczm1MwCkHpsiAT+tLO1YdQFms3mSBmisXRkmOglLo1RV8/LEsTK
2UpCSk18bn1xpLeKh8tqJAO7MV3G5TqNnYXdGvFh7/jJlyZsk/20a62I5GDC83qL
DfUaqRlEtWrxHRyOSKMLiwsHWTk2ngeyxof2lPngnv/kQHJXxhUXR0AY/aAFkyKR
zLu2aqm79eajeE70qzSehY0zrY7EGLgz39hrVty5kneUebfyYmzbyHdLYdYRp0U8
JwGDWc6Bc3q8HvhMrNIuDWDLD5Assj+WQnZvWj9YAr9RaPUKZ7pJflBvmdqld0mK
fndYQTbQ6Tta0W2jOJrUFXhK2o40NaouYrtQ6MgQoEz16e2vK9LWRpuO9C76xMVK
1cYlV0BpbUI226tNlYH/bDMxwxXa3oeIJ4XWAXCseS2dkkxGTIwEQupcwQh7IiaG
bky4BXjKzQr4H6ol9FReTzl9tjxmzr+3+QxIKxS6hUmlezTqt12LwZ61JtNR6npR
0pqvzaC/HxdRNh3f/a9D1RudpsXUmfLfsFGJSOQqCzQBHOlBSFlSXp6w3WdbQe3C
r9LxmgpOuEv2ar0eXEYJvsS7LGqQqW96SE51V5OexZFrJ9a9mnlhyCYBNyiaFYxl
UtvSseMzmEe2xiBaM1D5Ew8+Sp6nV7CSxtU8kADnMU7eHQwQZ5/lPhSFLxD9nKLK
SNvEa6C0uiDeAkLHfa2IL4NEuOSW7ad9w8TLptVoASnXTTZMYoa3wcv2KaMR+I5U
kB2lUvTeFE3cY2EojehJzx/uPqrJf1lROE9a20YqxsrgLCWfZhjTg4uYtC3f/r+6
eBjPX6AQyYjwaK0C+mUx14q5tc6u7RGzayhFStfZ7CdRxfPmcK9IjP5PGZUfA+Dz
iJqb8v3t2P8rua7GZlEuw0WmVayEOoArlHGeCLrDJzp4OCqC5T9WOj7O+Toy3LjZ
H/0cFYnHkAdZ9rKkZJSvPHqzghHTvEBys6y9OUse4+JZzFkVyPN6fKSjFjLuNewR
Qqb8+QmW00JeS8YaIyWGNxdRFX+w+cMrrPSsyjeATSVtVXv/P4SYmZcNFAff1H5x
c6dXy1hedIb6Zj5RNRfdA+ejvKqKt8/15qY1br0LTIBjteRNSzGwVjXXu13uEdcV
AxQgy/FDyzb7oEmBolmm3UUAWnxekskWLdmlz/RbUzaM3njtHJV8315RtdgtrG7S
jk4sh3s+JL9zXZgGA6yQPoX5u5kkt82fz7McrbsPhT2wy7iA9pU6s85bTtM5+1PU
tWCXL3phmUqafXAski74voCoVbFzOy1vE4tKrjUOu87RlkF0/Fb9KvwXmoTAMP7M
qKpvW6cimAmY0kZEnLxOmozb9wAo2fzefebEmce1rkNUCqQD9eMZkz8BMJaLg7um
Ugld+QUeZX8ORASSBN/116qcZELe8465eofrZej3J7g7etey5qgiLFGkOvP61DOP
DsqFvkuZT5c5X/Keq1dlOo5d8nr1/H1ijNyVoi7+s9OgT6tZ0ZCA6Q2qMJEihLuW
RW/8gYN6OmHu5wHBeziLDzvvvxdHfAiEJA7lxZLS3i6KcUDpUMLKfrTKq9rBaQdc
u/I4x3tTKSiv4tsXVVp95jGdDH0phj1hVos2iKVuVOXrIUz/S/TsaGzzIvBgYjTX
fdCN6bEVzOoc7pw9ObZu1LUiIGYacaNYXcEumktr0JUCx/TjHPCtwyydaAH3bgjR
WBj5JRX2cn+NefsY7EEPW/0PeLtsKE20CBATddvVMXOImUMMHLPkmVm00NgPIxVJ
QPU8UEq8qqKHi7gtHJCSGzL+yqXa/mt/sqvLufENEyKEOKnUgS35AD1lrWXHevk2
1MHbwxXU/Xm7MKU61fYk1L3PIEBAUAWyRDVbcEeFs2IwuzcDUb2rY8RW4nWvM+Ml
tnVl0zJEQiSw+VViV79OYUyxpLCka8MeHnNmtk61sPkYtpmXqvz3eSoHUDzmbDzv
0SgUyhZhEt5IZFwzotD9To1LJvT18XrRiaPA8weT0BgNxZKnIO4cu113oNRRmdIY
k00Q85FrEwnoPYAzeyJVfGxVhJ5ZmxBv0nzFh+ACQt56fFzWFFcreo1gyWjoL21o
28l1OYj+dVkb+BYFRYATwXKzt9SbAlbZu/jx3kcUpUpa4oOIb0Szd3gLEK28l7oO
0ZvlvpaONT9aXj309/SgfNqWKCQApNMUbX5XLtMefnjlg/6FiOd/9bleHA1O4uCU
KaPOxnN3smGkgLhWpSaeOkPJxFH37o8bj+wjH3mH6IaYpga9oodYO/eQTIl20dGr
SnMjNdQW9HPYtWDvMou/WC98oG37SoFgFUhLOJgy80OAj+822cJch4JIzx2CBAyE
aWSstRg3LdBL4jp0v7/TFDh4q7WCx278kjkk+gC282PnvvTuQYu8FTQuLdDbfxEY
EY8+oEpm46WzAQUuCRed3Gy97sluNA/9OA+HWVuSmH/cs7MnF/Fa3TBUsfYHAtL8
FpLV+culHLh20om9PxWRnDcV2+KunLSEPDt7PLnOpQthulRQ9GlG/XJOJs0EVMHN
PNVxwn4yu0197a1LZQSFjtt3OHD/Lp9jXJUTE6OTAlULzNrjqU/6v/xu5XUoKTLz
MVZRMaTm2fzAGC6wSlyugWXiVhdSk6219a4y1smb+M9NfJ9jXb9MqiBHAM9DIp9W
2wtA+CG+cs7ah/GjY/uNqwMXQX77jOWJRzPp/VzcsU4Gi80zojM1jotlFDECwC0d
lJYWyQZ9WAkLeFpTEG4abZkhHXGkyHJVaQtKkZkxP6y45IlQGwmPACFJtfeUbDn3
2jEEOwk5Bb9GO6N8CW6xFbw3c9CfHsKVWCP52b/e9npZntU8+xuV3JKxwjrNW5Be
p/h62TT8r0a6ZkFtn4AwfWPUNhaL41+KMDlkxC44aOo0glMISw2DCwfnZRon/+Z0
9WBIbyxE/zLqvl3BwKppeSD+e0Bnsq1QvA86SmaFqznRuTZQUMHUEvcawm+i2k33
/BZceZTU/OM2MdxEByy8gAf2Yoc0BWz5WM0rtPDdX8qEGkuBDa0E+d5/kS+kRTDq
+LGVCQ7jz6irOhQg3J1FbyUeCdeNVpZZWcnZp84eeBKZ+RCRVo8PsIyzlDAIQzZF
2Zxoqj/SOxcqEe8sHGbNZKGo2IWrqhRHj3SLNXipoJqcbdwH9yWCCODCMWwV5ijL
ZjV0Y14vGFK0S7wu44BpPUNlr+vJR+9MLxquju5tRgdnmJ+4PfzXBWlSIK5e9zHA
u0wXuoFljOOE60yRXA10OfDjZorzAeNhpc7nTOqhn23z2c1GB9WftK9BlNlzpXIp
QksuXECCFB7r+NEQvODNoh1TCJH0anC7rKJYua4igOn9rMp3VSh93dW7+fjstp3/
oN3p3SsGPZxi5vn6yvMqM7uAZkcMX3U6qZA4xgsyLeMuL/ujNxYOrxFvKYj0N79O
tayqd1HEVc+4fttkRp+whpxt6UrtJ0pj3AQxFi94ezvWWEqa0hsBACNF7vuYw73h
kCC+GI24rCcOBkexOPu38YbcBvOBZXngSUezWMj/0opl3PGIYxBPQl+YV92XHsx3
V08by4a4V6cAR1/Irt4bSVSwoaXTJc62z98zQbPpuIZQzh6/9/tQmAQsJlDZNlGm
Pu/jFilq0gqQ460SUReO6qE9mojfYRzsU4Ud3GSFr7IxKVCG6fkCmcy1Ec7o/HyE
+camNt9lFe7uTW1xU6LAODQJS9PUoyrm1PsT81B5z8ePQPbSchnFrDNIHz7J8MYY
KBU3RdzVrVc6kQxztzAxgwWIctcXJWmKFE0ANXX/AFrXZ2zEEu1zzDAQdPy+eJcn
m4qN8TTfxwfgtWyfJF26clzkHfqX50yhM1CUh/fPZ8bgs153zT7LaurXzgWYbSLq
4F8/n7ICjWnNkJnASWX4B3igoKAeRILOePlcIImAFxltaEPV9HdeWlFcnXPdZxiN
pR6nIMJMYWhvecu27CB9Xo/JQq7AQk3E6t5QMCja3vPD567+5GOEcwvKW4ygHWV7
sLO79WqRWBxZ/YNIl+CNivismbhnj8bG4wyEepIu9J34O4ISw5II+CsfKnrDBFBu
+3Jp/3a9SEKLDy/9UFFblFXXzElHJPGAJ7aKz8RsRSVrhACKyx3uM9CuA1wW3sq0
8UFJP5+zhRXxXeE2pO0Ceen4eURXuNdjHK7a3W3yFlu//WmJQADpQNTbCzp1eo7i
UuOIwiMOLTKCwG6wJt3Ybjsu5tNmauW7Cp6J8fnn7mRNScinrFShN9Qqk+jb0C+1
3MA1cBhdHEAIi2Cdi8JinwZ3pU8RYXBnsfB4loOY9+7WO7nlsRDREAWmu++VwCUu
AqeDTXMBN7pAdF00RjHAJEEpewXccyINqCONEOGLJldegWg0jj9ZtMSvsY5aUtsc
b1jc6EdQVx3iynGz2fU9Y/E7nYiN1U3wwQsJQ3aw1p7Bv5zvLwwNS/zA8Pr5xNJB
fgPKF58vblhK7/SljlqnBi6o4/pRRnqmhgK3+pxvbXbhAeMlgzj6SSgzw0vWj52a
S2w78xulzfpScDFGsRE17yMBeu8apYtXccNu2FX6V0uMQGH+aSSZJlF/nbmucrk2
UcYQboPA1KwyI1VanUEZucE73NMeM9mIxIWmYYEPbTqdCvBbYxVFCSkAHbwOgciv
FguxR4ctBKOU+OdyvY8I+1N9DTGUYMTMJv4NSvGgMNKpMf4ZYlRsKAcsfkgkgMGF
GsJg4q+dzU8hWRCocTefUDBQGQaXDD4abFas8ygzSIbuGB7OrlQYuFPsYZ0EIp6W
CvgTths9C19ZenN9gAHUq8dR+7pNa/yJUkCGkoenK7kgQspJ5bquULGhhEDkUhIT
3K3ig0A3Q9VtiIeEqFfn/WdRtzrnWXDPBQ9ibmwIKpPf6EpP+nL7wnLby2AwEEF0
sayfUgHHpYdT05IekyaUtUV6V6EroxzWg16kIa2pLvbrfpC9nKLv1ea/3bJsYZxb
9nSfwe6wOSdHt6+fHw6WUksr+yOi4508VJ6/INi2Bfcd8ZzwcEfEb0v7cxHXRxh4
He93xyAN2AUU3nYbh14XsDpk+eNos453pCB8/9pPIqshAcnAGj+L0Lfo9fTz67e2
hBaB5B58js4h/DuZcCxezUeRHg2LG/5nwJvqOyR9Fh+dojvOHU4e32myryk9NPbm
a1Bev8tTk52JzhaBTCeSTk9fqJ6FMc97iN37GWWicUDK45CGOGJWFzTMamF3T2po
k02eeK+DbweOsG01bBBkpmpletBZsMLQ0T++YEKlHCLD6gTi2zlSptIZgCZPI7Y4
kTUEtjBbDox4X7iUwtq9E+9X1Yih+oBY9Zu/HE1l481zv+rGfE1StwbhHFbY6+Qz
rp7qzk4uEXKtk+08B05UvJf/uJtd5zwLScUXTB61FZSwrw6fsLMnVAB+acxKCLpK
Igt2xBn3mQWe5s5bGs+29ZgethWHnalaUe3rmX15LSVGx1M/5S8Oez08+PvLlIeF
ewMIp2x0mCo8dOxC/sUst+yeEFmMNJe54cTdzUvW6D0C/FfCnupp6G4/yxc0oFrs
ngUwMaYwnQ/VxjvGyP6Znx3x2xX5e2KGTRkfhIU8seZH+T8lU+RHscFa1XVMRHI6
1ob+QyPVIhYhKbIu3n00va/SoNl9Yv34HKaUNRAf/+WtekWdjiCBgqPEZRU9zZVW
hlWcy8/19bFezCoiS272UBW1T/jSqYa40yqakuSym1g7zCJMxHIeUjanz/pARw4+
+aZdKNOexcHMV0GXI2MXqdrxAcTgZCRst5qtkd+5piaZNyFb45ZylRWNWBmv8X5u
4GaSVRaSJaz06SoQXrB9OM46CcEFlaWHF/QWgS5v1mXwxTTU0RM+acEoAZ+TdKlS
h6muwu7WizlPxcfmRXF5wjkhPYSgU8f6LTaHIy/ds2aXzkCqpdcz7kjbXfIfyZru
8R/fb1oYW4doc6F8R1aacJbZOjzto1Xg77++I+mPNNxm/iPHEa//uktzpUmt5bW9
SmeupP9I85eC48e6B9OKQkQoTKyRLSFGqZHX9/AAMK6OAWDYo5G1KxDYjLMAlrU1
rdJ0yLTS4N/q1mxDyQi1aoeo77fjAnojpO9ei3+VlzmeOxLvn43Lx4ZT6gW4R/Fk
uBImgf8k2AhR6Db30IQ44wO18Y2HGZ2F68sE5SYbbyFX5vtCN1NyAqYWyb4/EIT0
2j4SZfBcXOnll0DVIj8Deq4Iw5v2WB0I87E9aV4hcU2PBzseWeui5mxwlenMmaML
mpHD0JGgBisEd+RY4QKs2AGmRHuHWXTl7efG/s7A3qylFnrH0QHizxSQkVJsiLos
9DwRYEwWBPxNiV9Xg9RzMtEJMr5VYlnUv1yxBjvvj+MQFDkn31yp2ippS5wG1h47
+oBc6xIZ+pQ87VR9IIXLCdOkqDrzEQDKFjisrKWfFtQm1fQ4TmegYVE7t6CoaIjs
o+IDz3gr5Hi2203Gm4Dc6g2uEQFOOd4+7n/5GVdyN8BPWSQALpsf/WG+MjyuDnkE
mF6MQuMF6/8/fkk5Bh6gh8riXueQTgbc8R+3y0H+LfSczcdpagpsokDyInNI2Z+7
lWU/7bJUGatINuPO7K95PK69RdhMvL4sBCUREZkMEPnT98yQwsGzanGfPagqt/do
3fjcRAGe8ZUeYE/Qc0aMrd3iXiGfHG/84klO1wom2T8TDAvk1OL+R7Cmrk3ZIlfn
sG3cllXoa4hNHk8MwTdN1gxJV6iAxUr8AasOM5DL7kL96Y+wu30c8ovqkF2eyIY5
k2vZm3lK/dN/EViOjClFkiT7+suevLX7xoo2bm5vN6P1fQcf4rHhufhydm8sD22D
iu1Gda8VWCR5v8ubt5wTNdwdZsgsyffnbS3A6jJQwQnZ/quVaIj6O5VsOTxNHUqI
i9+zriWrJrnwlFrGaeWvMC6SROXQ7VutGkFcCF0ZFuRMDfH3EHipiU2eOkWzuFlo
VabXkTBKVPVhyvvI2rC6qse6BVgR5IUKdIks+N7FhYmPJocGUsgiE04YvYfVfqkG
nZmMfPuNNS23iqj31y0WfTpcUgSKRBYgNSp1ClJVTX2Yj79UJWaKj4Cg8kEA8qAZ
Tw63WUWcYu7tNyoJaTwcToW38MqBLjRfdw17FJwD9iIZBmiTtnkIGflVZg3dj9FB
PM78n1HcvcQuUiJEhHGi0a7e0u2dI9R/m6u9hc5Qtn2QLAIqOosR0Vbkrb8Wt3ZH
s4XP6MdYKhvkpqzATjj2Lc73mrnS8+DDVwPlKYswFSGt0wQiacrPHZSpJXqW6GuT
e7r9Uz86rEo+d2Bv8HcdHR7zJRpSi1Blypo/QfYy0lXukhaT5LN5NtpVpDj/Yrk2
GL/VYUfJOd0mZHEi9bmsEnkm+2WcNIPXr+WB7/9r92N/yKfkR66/yvVNSk73ar3F
ZV4DqrA6HJSdA7Hgo18SzrqtO+hwNfiX6l0UrJmiMgjoDh28tpCZI4GkqH4Wn10i
Whg+bRXLf+xXlW1ztXA/UaD1t9i60p76X1bC3R2R5wMVJtSpmCMvqvlz+QnD32NP
bhPRZ2faydK83WiQMmbf7OENnEZJp3nGpmxG7bTl5hpQjZw3wvASPkXmYVaJLMA8
eyqdpjCEzHMhYdvJGuM9sS59IsAU/IWc1D+8E1jYwMPoqvvcbfQtNVNw5FyS0Q+g
ZWjV+Q7YzY0vTfAAJFBTRd8z/eGuXwTTKz4de8xyouSw0yQri6DbvHWZJ0+u9R1o
KNCZaQvwp1VlZi3N6ij4OpVFOyYTigHcOP1aAngKFrC4BkMpMKD0uQ0k9xm1XeyB
vufVQr7jknEjLf9FG1DiRfoE35IAs4yuDP6Q55etlfD9cHst78XO2vnhO/Hfkmjh
m2GcNjUDOIDofa0YURAhvXFKaSRw6yv/vi5z+LfffNXKzuWl4gjEdtP0xwTH56U5
mc2aKSdSVJ/8mSqB9HCz6QZR/CoKu5Dkk5yboQoIdAnAUD0mmehYQXiffZ1GEQ8C
zxwYggtUufEVT5I+P8uptc45BSCYvC8cJB/NwMGAwCQP/1HbBvU91kyJcTxv7Bhi
iyEWp076N47b/0HDvgXlCwOKhN8ikvEd2msOft0wkBL3nBAr3xKsnQR9wIrLWKJR
nE/8p0Rw1AQAmlZlBYiteuzfJdfwkGISzWm3JzaDZepKNOWPKPoK+rFQn6pNUxYK
3LkwEnTC59eUAnAs6kfekh0Q4yU5yf4riQmKZ6VXpyCEzjHJQgk3/Vdff0dhd/Oj
mkdIHqd9RCqAfrXgpRmOHQgwFq8GFGrW2WBUoEH70Kd5rPNZ2ZIIm36bkU87/S0S
Sh8GUMzWV/GubFRaoJXycW1ughaCGrXuGmXkgvVMiTA2ZglHFNi9SMtt5KBqYyo7
QWEvDatpUYClJOlk3cxFNw9XP1uC2fmM4ogiLPSm866F8WMK8GWxE5d7VWLWZ7l7
3mROsXQojcpApDgI44V+uWx6mfW72nQAiiGdna45ayn7ZkHiHxuc/Y3o5ncHxEAt
wU95kJqXj+XvZgzjvXwao/qHZ5xE4GJYWMq65gGB4NPFct8JN0tm3Ce3xjqX+y6j
wfLVsVbSTNEZPUdIaIJ0pq29+BzwTTiiNaH1ExDr12M+lfW5zi3ZyXVKLCpA7sEQ
HzuOod5ZPMPXGKV2PUq/rOYfppqLsFC8uahm459XRsUMW6RM/a/NVnOoRyU7FOqO
A5aRfTZ9mjFzlJRMM2/eR/HGDTLe7YA8qeSsI3rJVrOZ/2WLpFkgw6p1K5o1HoiQ
gCUMU0G2nTE4Xsre8ZmqpQPdkMXBwjoJ4QygHga39uO+qBbnYdX5s/JIQdeP4h+f
AtXCDfA4Wxm5IKZeUwu6heSf03u17D2HToiirKO4hCp/4giNfDVq4O3rf5XMEYCx
o0D8LGiFXK7RqXp2UIrSwARI8XS3Eu50BlMn2yCGit09o3uzvV+0tg0Ow1ktvBM0
fK5vl5AXtbD+PDVg5CFCGTamkUPP/hbVQBWkDCHje4obOm+GyzwLylYer3E0YfOk
6VoRscjkxWuZTCxEzek3GaM3nQUuBk0nLVV2wLs1klPVj68eY4TZRLnkyHJiEGFA
RDqNQjdXPaW/6ZHKX00+ztlsRh/ioWS/8oFl5uszOKcJ6aCej0K3dfj3ZTZLsm9u
PvfIoxiNjw7Io3OMe6PQznAGlk8GIvnbVMZRdXBacm+Bv2+UuP5acRdiq/XqYXsO
voLLFeAQm/x2slbqEIBVfRynIijThsj8ANuHw3LxTRJgaQ6SgHk2kPB6IgrZ25TL
aQ13GFrSslvVYzUeU5Qxn6JS986eCwmtNgg36cxFC0RcVQi3nYZy3HqJwcN+xtT+
oApeExgAqN3kCcBWbPbEQ8Aaq14dwjgr9poH+BOhMlZxENUcZB7h64Veg40V/8tz
hDUzeyS3LFxT8ZDTGzpQexyNKOcMJ4/TcTi23VCvkGdbV/w/yxHnisnwbWTJckP9
i0BHKac0ab6Bfq4ILy65eH83I+xly2tbx7ZkH1ibW02rdWW7YeQYBbUXauq7+2Yj
I/Ii6HtnsFstYU3Cp0PymFTxyIXP7byYHFK4WX/mCr4r/xlKjJAQtCoi1Gj49EC6
iH/EpR28dvTYzETnPuS9O/sDHLGOh+Xycg4ZnI4qcpqp6mGPP1sFFLDge1VDQpu3
40/uPyQoP5WrzIEVndx1+QR7QxcEEdGcY8px99B/3bAHqGk7EckyGBnIgbKEINiq
04oagGBXJZCoqSMu+8EX/c91nrdUTAwfut5MeXwjRoEHk2H1TcTzz8RH5OT2c4AT
ZQn+txEWj50+U+QeoJkJO+jE2MQW8fVMpdfrz0A2Bg59KcD5xGdyfWPlzGV0aYcu
6JEZiAU6q4OhZV4F/PFxDPBYekLg6weFHnXFTEhMlYJ6AGNb95pNoa5B4GHUyFbq
y3teYio0GfubsJb71JzL0DlMCpOSItEm88SfTF1gngt7RxHo54JgDpX8MUclrEBH
xB/bulOX9ELAhl6qJfiJ/E3vvGU6t8lP9WnbRVk5L7gHY1jYmtTEJkkne2K+sLHv
5yV8o07+y+sMFB2QYAksamLuCz9QAXG6s6hN5W0owo2+m0ciOkBt6B9+f9o2ownH
UlV3byyzohocFFx7P+4BM4LcS+efLpIJBmZ3XGBpHuEyMQyQj3aW2CRS63m2ciA5
VqFMUvmQlgB0/seaSWmYZg3z5Ep3FNHHuwrgVLoZIpTqpYsBHxvcT38GAkgOsBWy
8odS96dUlau8QzaOB4qwiehVMcndM28t6Yan9yNn1DVwUMbA8n56xRQrr92I1uUw
RWWUOJIxb4AomxwXgJx4fBNfvi5yT6qNLsjVEIHAlFKP/QpaWv2L40CMMYt2Cz0+
pVwwWxeZFngRExuiN67PSuxpwSWHJ3V9Ugv2TOKYea2fZJ09g3dXpqhL3eGc9m65
1v81F4dWSGbGwenywJjKKzZxV01vBRLNczYAkDpCeQqp1LqKmAQ+37lxWcCPneYj
VU7bxRJ01k7u0lK8C3+YB9o6VbszdjMc1za+w1YIrnoQnwx8L8kpYv2aNGdVALKF
jN+2yexHux+zN4dm85a+k1UhekvoJkSj2q0lPGxSHrRjgLgNfsbJtkSTTPsntWuS
Dpqgmubu5TLAlZ57/xGIkOZchFBnY1z6alXu8CSGyDotob1mxICMgJFlrfrEcykF
LzHPMjJgyQOeSyygSLDP6wHnyetZKJzXL1ATI1um9gs6AczdNW4OobHHv52SXoki
IAA/wPikCE7+OEDmsaRVhh5S05lYiIVIE6ub4vTropu4H7UnIQaLRLh6RgVajD7C
POX9sdLSIJ4nG0Jy+0uXvkB+TlYoQXKyCjrnUkK3yZaAjx4gtmw+FKfcweJvavvf
BPpxtszkgTgpJtzpQ16eg7PByKloTc+H1BMqFA0r9FBtvBhOJhSvMXQxvdv7E1dR
s0CuF/kJ7xx/elrAvB/NrU5B7flh/GUTjCpwVDSLMegshxQcVAwB7TV7wJ+jS2+d
JANc8i1P+mvweI9ka5ZXEPr0qVRyHeKQIhbxHgCFIq4DJ+I9langpWYqDksmXoJ3
k1STsyGNwAqfTOij/5xRVgXzblSR9r6VenW3Mj3pZe3byNEx/dsdN4dusCyGPcDv
Jg1EtWwlbZFCKaGCeJQAqEqmnm19VHmV3Uv6qB8lnzIKP+gmLzAuHcNlmYbGhfwc
nh8RtIyI+RoyFoXfhsj4y/qF05U/5irpzusz9SIYGe+SSnVK5gDm59b/8kguU+V2
KBz9M/116wtrc4TXfQTRyVxaElqH/dZlcbh+lKDFvE1TNiVTByw2OjSz2xYyC6A8

`pragma protect end_protected
