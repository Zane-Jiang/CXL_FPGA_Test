`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
fGIuZEoBQI/7XDEQZPRXJksNt8eNK1iWatsqGvO0MTjiFu6+rUaVsfyoGlKUcqTr
0qmFG7Ec/kJaxD5RidYNFWp4ovVx/hRiHZ2UBopp4cgQb2yIXKqs08M0vj0VP3WN
5DctDWRGCT89PHK3qmU1VarbEX/gpqaXdiohia/tBkQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 59872), data_block
s4AxRkv+1fP/YkhYercjotiNyPdlv7N/kTJdkzKF8dhiT+OmTUe74eP+SRdAzXaL
JgE7hiAaofCfkaW3jjPrBaY9iejfxsUYS6EFTxX5c9jnos/JrazdptH1svG/90DM
CU0yYlmpiCNFYWaZfxpLjuOOJnqdvd97/FMOvLCfsfaSq5D0kzzrgwoaNmtaVHmm
KuQrdbrDsOOC8RpeNS122dj0WfANngmEcycuKXV8j1yErLIEZnIip+USi81pPBbN
ku1WaFdgxysIR08uJzch94AYfj23YK/gPSKHtxBPrMC2sdSHiFfy8e0KGATYHeK0
jLNr0CHFwwOBIAt6f+iBi0Th+QbOi6l/x6drboncke4oas0TaHXBp3AZrqY6kX2O
8JKs0W96nm+e8CoDpsorPGFlxJxr9g1Fg3fkfnm8wA0tU93qKuMgW1KnsR9zgR3B
CdLF1OWWZNJlLJ0PgVcFaaubGOVNXNM36JgUrQGouCHJIx1OE06YYIkVJpFWN1w8
ZPGafcDyYq1Iym3H2W+nkECLgoWVe+p40mO3sNXT3wNTLDf14yddQ12tBovdnW4o
FyuQ9QO61XxMq7Pw3VGbqLo0NqNRVqMNlstFmIHBiY6B15wQhA22VSouq3Cuxwep
5abHTuyFjFMtEuqxIkF0vAvR68nwl/NvVClsPmqB6a/0iG4hCBuTAVsHF651BjNk
x1+Aoz6BTHSKVaeeKMPAGIFAw6hfxjgdkJTFzTIRXSzWV4YJ3awunEsfDsHEsZpA
PnsszAFyF2wXQQic5jfUl5PoJSBbVuoQyEkmSQOx3u8Qx44lcrhdOBbEy+NvUyv/
SYzHdFj6SWmHAg/XLEhrYq8m3ADvLNxNpbSF7vsQFOlDKHOuxp3w24nvTXJAFur2
1Pl8OCWictwXzSGuR8/rQiEmd9ZthZLWyPw/XJKo3U10xNNVqawGjHHi8e2OrJve
zmgfq497DUXzcK1Q0YbOMtHz4faROiTDzvlRgAXV79p4gt+HogrGFtButc5GxRBE
kf6nwtQjLlgvLhtj8mvfLoIH8cchviiy6qKJrUN1U17xbPfd1PSUGiz7WqnAwaez
voJ99fkBMiIB6PPbXFmAH5+ZW+fhILv0E0Du7SVZNFSYoG+mtUznA2Kw1fAyQ/kf
G8pcoQsAwDAASDy7UR9W9sLQUAiGH1s7AlsvmUi02xko30ljEfLo3hlZUQSXSe7h
S0ewtFr/bkAwBDgXZ02mo7eFDk4ZcOVdw1oFRSOVh05U8ezXTMTtt23tLT5e7Huk
WZNinMIERhxdoWvVoYxZvjFFjHdmuIMLtE1dQ65TqhDDuSK60EjAN9Lqhb67fx2Z
lVgOEMb1hh8KvsdrFEZYxVZikD4FWR1PfeY4cwmYYBdnAZVqkxnjx8yHpPAGPuSW
HEma6umRDNLMX0Dtx18GtR9tSHkW1cozzl7UiaeEAGNlE622z6/Gism64ThAqhMQ
m9expsfJBW4x70EQtX+R4kEZ9gjfaI7G71C7Y+SDkvH4rOsRxZFVfmjaLQa+rMYw
gGnVruA8TCHVkNHHdwcIPQ94d5h2FRTRo+g5c7g8SOiTHfDP3ILblYBg9cJ2X6Ri
Ne0K/4c8kbHPPBhSduA14LyhfkMxvJDT7ezLSBRy76bwmEEwh9YST84YInSuYnX1
wFi+8B67kukI+KN3BUk4kNIwnewTYP74JeYHl00CdcIQRK/fZewbe+oV0l0q0jBV
3vV5adEE/ul4ItFjjJAy7K1Hu+BMx8BiwvZ2tYVN+gAk7R3QBajBUyRaDTmOoyX9
qVXZLYjV0zn7rf6qB3QzVx1Ad8oH3Kg0Z0ILBvnCIICnPstdqGDDjR1tbqG3VLYn
tVZtk/4D87NbC3iKJpAj280JDt0aseYRZr5J9FOIYGSaesElq1/5k5TYT+SPRh2h
MyvtI/aLEEbkTiYNj6MJAy2MvZyRxAclIU5Ca9c80M3X2pjTWw1t8eGO103Yaf9p
7oJipXTe9ks9VVa+AkccKUMFzhp8QE1XxxvHCPmX2pHe8RA1BdbpG7L+7W3v+fLv
SLhnFylaP8PZYSJdLwkFMvO0zeo4qvFOOIlwf24lQ1ryW7l1fIt1Szyz1HQTYDWK
yUzs4C1reGvwcNikrbQEnWPKzg5s8Nf20Z4YhQ0bH1IorxBzl3l/GqF+chmVLeCH
9BL+/aivxjr/hAEGv+obitnSgc+vgkQBsLwOSU8hwaIB2uMiArfdD1uidzJqnI7y
XqA/nZPSVyRV/J7udttdvwXsouO9nIdR4ArmHulXwIM0K49lUdOg+3VL/vkEiUgy
FUqpjeP3A8tgNquVnKrakLXLaKLoXaVZQbO1AouxE9wo4JGfF51wRMwgrj9gRf0v
CQRzCiDtC2vw/g8HVMLvvDQ6vj/PqqI38rtvWh8qcmgRX/7cQwvhY2vEqedflrQ0
gIYAHtr1YNM0FCGX+GmA680s1aqV1oS4YH8VFCzeWhbeORw0CXmPi+0Dcz3U0OAq
I1Bm6WDI8flRYM7sT7y4vCw5xI0oMZjzdZzeC+BAfW5ckiQKkVkm26jzWNTW336n
HME0xjQLuNynpouLNnfkELRElrq1SdFV75p+vInt9QU3FVx+tcgtgIWEsEWS867G
KasGps8Fdi7Ja9yTcPOp1XjbT1v7oSyzLDjatyBNTfNLQ7d23ePpV4A7R2G5zPk6
/CYu0BHYpPxUGIDGho7Xwf1HM4KQtSpvO0RVyfVo8AN/0SyWls125FeMgTTb8St1
dHIndULeXOqKIXFewsAAb0sVkDQsi0fpTzhCObJL0aEMmXTi1V6TObvulemkKlqj
HLcxnJIxPgiGccDh5YiuCb6jkx8YjcpmxKIHE/gWSD5YQNXFYmQk3XXsQcp9F1iL
9n3nGEQEsvo9i/+GZ0/dkAH1qSXLbwIxbBwCNZGOYIlO2NxDOq6fTDTPcdlM5E48
eylsIkmdQp0dK98O3PfZolvauqOkYSllbBtuS+I93o0vUalnDFix9SfPybm8HSd4
MSe8c3iGdlOeERQq4BHK/bFC2NlnqxDRddyZMdNrSiBVHXYlxVwsDosVovRAqD9g
3pR/K9bes/tsHpkkNmbyr3Ug8qXZDvuTod5GOWLnhWBIQfkEDk5exhyLKdXsfDeY
i7XAUNm3aw65jAEDac4XZcMDkQD347x5seOXZ16i3aJr4CoZ/lVHNqZl1iIgkF9y
UetCdSeo4MtYgCEFmOgLsQMoIdN+OFwAqlINImFtE5e7FennjhvQ2KcHZuKzMOTl
cb2HW0oGKtkAj1HISyyEt4lv+pjagv6X50LMme41E/K1tR3vLDShV3+VM7MB5bUz
iYh/JW9MfKYmlvGLHPphpSvu9eVMcP0YXrVRPqqJKZrVUOeRBOCyyTMalxYrC2do
yp7Qtg0kJQN0e9wMtEAozf0WrPWzKlJrBTcsH6e0FhW7V7HGvyszHhyiLaQrYvut
gHGlvIS9wyw5r2fmmDBcTpprR7Nb7AhhOaIbJXxNO2dj2goyuVB7G9IaPPz88sdJ
ERO/ZfCs822Bf7hoeWE4de6fUkeYYDksDodCtwI4fmVqyk9f9ZFHa450YvdiiEHX
bb32kWucTBMNbPxz8SwQ1sIzqPGJaSPxVt79bEKvpEPUJZzNR8PY57vucjAMKDnt
D2xtGtF367v2q2pxJbxSSFy0g7WMTGwVJXHQ3jWQBV8qgqvFBzQ1xi3XntE/LOS5
r2S0cVFtm7+HkjVm+h9vjMnXBtsEN7zbHJ8f6ekyYTjaxSG7OM41H79WsJkeIeIt
QFDRNp3Unj/NnHgVcMW4WUdT2ujdY7k2CHXTAB4xFf9TkcgNildaDuZXyhOs6c7s
Pp6/MNvU2cNzwkLOM0tlLK7SO6AT+4ihmOSC1O38jKz5S37g9/jUR50GQ/RlUCk1
fE16TcO9VXOI/xhO0lEvK33+Xb3qwrVtOHSJWJ5KZQnArM2TExmTgYvYPuwn1gpZ
ObxMM96Iil79eoP2SHCScAyNzfSMEGOqxll7p6Ecv+Jc5YwHHf2MDzYp5eh0svmy
LSa9++3TgUxmRhBdLPi/prDKOXglWOwag6i8GI/Uyu0a9crnnSbZiGdbckbtXuoF
2QNzYZKzJLzyNxFIYExCqI2joZOejLpNzz4AJ0+7y2b8gJhSIt49xnMGDlHIuKp4
jgLdsVpIYtm0g1BMdhU+Xc0Nlwl29h4XNdPgDfe7Xik4akZHMbiBJnvOJVjWZQGD
MGsDCYlowKRfIWJt796/u9w766ueXWouthw/wzCGegN4QBywLDrOU/IUPHPOngrB
Jjm3UgVtfz56NxtvTa/k2HL0/iJ4FdHu6ARCBA8iEMkzog0/vJFgfAhivvS0Ktt+
jXuTGbMORwLj1ZD6iubPEYuTuruWqCoDGIaLlpOLjtx95jQBy9J6bEIBWvIPC1Lr
UDehBBk8mfqOEZywjZjD7H3bmpWDzfoD3gZBdU13W3LBkiaAXssJd9jWvI6bH6Ia
/zHLTY/woGYuSZyqV4uNaDA2EsQ7bfJlKSo/SjTEMtyLJ3P7R6Ihm4XXQAZTwv/j
fechmv19ViIHTKDFBzWcTQpte1mi1iwELwlQ4WLXfA598hLtEZG2aweIPVvQl319
TW5FnU2c8m0JgF1wN0bBdr+LoUhwKULqPc8+DbOWwmssnm3mcCYXBkD0jmu+7IqW
3t3Wj6Nd/5nWtmasomeYnZ9XustCts7b3SWegYn5ezebBUjLu3V05pDK9bkbKSMW
/u0C/dT/tCtcN4PGI9Ke9L483peDfDZY9kb0nHBsQjZuydHJsRGdkR5QDuc0Fv7Z
cx4mnCOZZVpwCcQ1WOF2fzugAhT8gj1g3obQIhX5Z2qL4nI5o4J1WfdExJlp35vX
9e0/TJaXy3CS9zeiQUVh9+hCDqLD4jq+k5yWhOBlsvjau4XbcoFCmoCMus4o///n
7TXiSS4946WrCstTTGvbS9NTpVlNd/uJvoF5jsh/rTa7H9foGBraboQJSH6ROPHv
SV1fKFeeKMnWa5JWfFxJOFbepb1Wqw4xtCW4/52RXdMuYybTNA33wHKAjie3J7KI
b7y0TAx67vW48Skg3yY+o4qe5sgbEyLmlLF9a2AhabhoD9rhY2iwCMd/HMfzUeDO
AiqbOx6SdykHvRLEhP6JiVPPsPa8nHioN7mZf/TiCQve/Fp+rmL1ouzbhFVfna3S
w9jndDrAq9ks01/BLuzCvGvCKTvh2wWcCSZODY3Sb4WsrDzfQMNVjLLRSAMAI00g
VaEn8Wpr55PlTXWeIBiDv+1TQthfXKeq1jT+GXdjRNASz74I1nnAXsVXDr2hOabT
0zPZ0nTD0Q3fMFYaR82NWURMjIGb0BuNm21MjpybOC1InYg2R79OepyJLtIeSWoj
58JGyKIIlBkgs+0L8d/rK8k3f41mCgycInEq3LjaVCJTCI8RsP12+kEq9U/fOxkN
pW+aRvNAJFVQF/vJEq9At9497MnLYEvsZQHbz/naBkxKgLuAXXSvLpflsSwQ6+hw
SxxRPgk1Ze79v4EAIOV+5tYDOIu7nvQt3YL8AMqd2WXM5/Tv29shwoOwHOIHUnWx
P/hpD6gOTsfKTSv6cPPUQnXPZofzYNoMhdYunWWPJ7imv0VzpDSqHU6KzT8Wlxx1
dEi0n2+bzItcg9qy+KMGAST7HIcOmVv2E0Un7bkYUPKe5UA4eEhDxbnwIrViCCjM
eeF0bs6GjSLEdS3YADpc444xYQc1Ydrv4zrb2QkHjdxTq0XA2UEb0U6+Rn4edTN9
tU4KfHhSkPIEM4Ehv4OQvbNfl41doRadgum6YigQwVrs516AkWaOiOqTfo6xr+8u
dnG1L8ky2GuqmN5ffhT/K0jAkxgtO40rVfT7cmfeaegYnrZ+oNWGxF7S/Z43NYz9
/o4PDNoZG3N3TgnN1+UnxvzuvVLXqcC+vVNVIgkkZcxVK44FNPCfvJnDuo7/8qCL
EJ5x2Ks+vy/ETyzCAIAxnsdi9GYgJRX7s1qG4AliP1/rO+Z5TDIKJVK58LIimXZ3
jf2LGup3mhaLtIIGYCxD38y4rVOMdpj1zqZyagphVIhRKpHq1Yp404AvDN/qA5Py
8vGRApTol9uSOxasu0DSaKaeFX17OhzVNFKftnqy7XEa+IBtmokDemAX4bSZRfWt
VjijvPJ+T8wJbGdIipm1u/6J+V4PzHew9/lensMx+L0Qas0l659H53aL9FbAFH2A
Vo3I+uYg7o4MxpQK5LQm4hok27wCyUlYejzX7WxOf4FM7CIeOhyQkwwbVghzsF6k
9t2zw0yANDtpV50WEf+RokyG135lt8rbJ/WwMYjEyY1M6ksk/Hv1HmnYwhggsnSJ
9oAha6pHHXCIc94QBzCI/9+EjYCSKf0sklT+5rn5omIuw5DL3et9em2m71Vl9C9w
TZvT6HXq8sZnLYnmTV6teX9N2kn52R6+UflcuxPQerToQF3OH17tMKKSY3Wo/3lZ
bmDo7o1xMZBe3K8i+FL62xgzVcemyhxWimEU4ydvGUYzm5R2nlATZyUs16I2227M
LmE0J6lNeGlJpJlgAKR+JUaN85B8eZdYZLe1ilvHIl65wd9iL/mqmnk9UsMLPS2p
9TuSJUu63Z7fNCXd5BLadPDdCZJqLpR8vs1C227jzbA/hEGpypF7MG/BoPqhvlkZ
46jv0gYMTHcRUSMLUe0al3GDQDJHbyHHxk44+EiLIdRIPku5LIbdWRTixrM3si16
INBJzZkBzlCxUnoEhIWYFTxzGleri7lZvNg+m5Pm4UTrWV/YHULJ67X8t3y7rzaz
mLMLdTlwBAtKrt2IF0CBtVBffBshqeWdazoKkbpaHxZmO8NViV3rOTUMPtvTvabO
EKatuzEI0bcGyGW1p6ZQYlHfTr/DMsLcy6YJfeR4KaYFQlpattrEdm8piLvyl+Qe
ajY0O6JDee87lFOtMepyZzp0SGqtiAUnTa5HXOUPvoa+tEAeLXdO7NuQjsRiBrIw
/ne965IdzmWHtakmVZrVkZz8k2uZ106VRvUTm5YIgB21Om9D0GQvug0zcCfUvjxa
kTVsqQENyBu1K/FoWLV6sZmNyn7vXPNaZcBH1kfmvHm0K92FCnA7hbgZHMcbBrZT
s6pd9haqW3pdG7JnmoGh2TNTB90lH/74OBNK53zPTiawnJeBiPtAlVjvqswEMb3J
nmEYd4H0oo1J4fxM8CzATRj69N6BkPlhJ5xIZh5r7/AohEfT32ZNDWfjYVHnFNnN
NTj6wYaD1bdwJFjuvYN2wNjDeLGbZJDLme+CQf/LVS+2XV2mIGKBis1vMSlPFJN4
kSBs9UsAZqMEYX4JXtzglePjAZHdtBhLpuQoqSoCkC5Wm0RLEnY2Sivxfhcbhszb
zTYp7+iU5D19/aNx58h1/A7VKb0qKSnV1gFYFgzZ3y8GBGSf+7pfl1Hax5BRg4Eh
DKk8+dil8wH4du5A9CYI46CUbMv0nTmn4nfbklXgvvhZtiWtwG691T18YD0ztSXe
XKQ7cpG4pcPP+l8D5iPLawe3woO8maT70CUmlUiOeg4Y3jPUbZwtRRUeWuirYVEw
W7xZmfaMzcoK4xk7bHvLF3aFT3KPKmQT6okuYaYpdWHWe10FxvOkApAKUePepodF
ZkoyiEYN2qCW4p5Yog4rUtZgX4UFaHmRlKKSMVgYZuXcnCMMlbPiN0XEH6JEVcMB
Aqj6uhjVZR0w0Rui+3ttoBx+qQgr5KFTkgl9qOug92XHvbSqQC8+7YwQB4DMfQQO
64WFTwdbOrubV2yZ5v9Z1/8Q9OOOndwVYl7OOWaotOGRSFZDBtaAlvSWZEmugwAv
oAqKrMkMDz19rEXeNVOoQNRyawSjFwxUCf2jHH3g0Ed61AascgSWB+1izz4888JE
RiR0DV+IOcNZNg0qLDK0L1RtWm7Z4ZnqmE53ESrZvHAfDC1zUu/NKAPtm/AKxDDJ
Di/XUA5fmqp7iCPecsHkXN5ZJiv6QIOo+uhNeIwJugAUbvTBxruqRbTqMODofGHv
1gYxqY3vCdPJ53AcipxCnP7fqUUrBraVJ94y9Cn/ppXPxgbUaqIYqUEQEPk7nxQd
nHxndZGYmKvSEyZGBcBM4Zv9emWOISG9E+6kqZLuBt6FoeUFKseDv+fdF4kdNQF1
qb0RhXUj1srcKuAzD0SdmMIyYKBfR7woeLW1y/kPYQqXgV+3sRf9oWkMWPUEy2Ft
RzrTnQRRQPmdY+EHFTgAokD1KEojheXaVjHRSVcxpBJNqcIrklVsHy1db7/RDDkC
aC8DBLIpluoL5GlL28bJWi5xMUcABzdYEdNmNXpzr1pQ2kOwXLSLvCa7rnIYx9Kf
gCjudcvCbmUCCndtut+7XdZ60wqpAUUdd6k973eLjsxRUL6bCot/uJnVzpJkMXXw
+Tt5s5zvlbtfz+7TvKOjwOfReFTsi9yfc+U4fopaWKPWFPgzwvLL6kDo87WusI9Y
mLYaK2J0lO85CpkLKQz//ZE1/z8ou+XGpiCuaeGtx43JGR82U7PVR7yzBxW5AQPv
lZoD1mFewq9yogFSlk6q9FAtYnRNRlb36UD2I8Ufkgp5vdSEnNYlaRiue+yFG/eN
jMGRM7csNKwwzDVipd/Buez4qGHE2zWfYf0PjpCxwA/wYDb47YosidUQuh+dGQYD
hO5lAzBnKh1a+D3c4tQTIO18x5J8Fj0NF4hkwIIQ/dPgUXEd61SYsUEAZZ41K7On
0eEbkMhirjx8NJWatE99PviKFqHRI5JbjHZpNVh5K+tcEJ5OYNnXtYwj5aORT35w
fm3wQs6pd1X8+6mgxIfHB4Irrf6tGtThhQS+w1JbWpPIyJH6ke9KWJQjhDvb9RWh
lOzTiWJZm2O8oKGiTSia6W308OFYVXzQi6qp0jU0859xLIfN2gk/tpR1Nrm+dW6k
F5JTht0ai/R6khM6J9nTSVZxMXgBymhAsvocbQ3Q+aCgEnP9glQuzAMiW7X+VoyJ
WCwYssQUMB58csReeygNGo/NwjjJfPSrFSVrMthJDhinYVdZ92cl9NcmaZ4XBgG8
mA89JudAAYQQEt/FIS/ojVookie/QrNt+t+oG57PhMCFIasHIpVQyVVI28WrQ470
2oSrAVtAnJ/3nZEIdiRFABgLiOO6ydQ/BZDJzoTfg2d9mB0sP69FvXUX5ayTG2rK
7d3xcRwXmqC4AVG2ifLq7UPiqUP1kNjjgrrAc34j1V/Nlz5f360kcdQceQdD9qmP
E871aDhCO1o+69SpfNYohATtF/qZyDvqr3sNlx97C0o7sbDhJBnYXoUOqelgTXK/
AyJQR+qTLTfvaBscF8YkDj/UushJsq0p+bYZSmWWJPx1fLVDbHFuWX7iZHR2vsJJ
cuJM4fo/FQZx0aMRr4IRKyj/aVSCzGZlRi3u1btsSOpu1eCMsUDO/1JAo11mpKVg
Biiok9ONW1aDBEYc5hYRE8kK55c2CqcoICK9szRO6Jqn7/HzDJuEqYk/0AXxUbVo
um0vfvcPFToltvfA8lBr0V2AqPR6gCBxi8Jf93oRY81Hz82q5180BsqmeB0dQNV+
sPSjE96hWebFjvh27g6tS2zE/9FmmzwAqpDzbw99baRTiVg3DoDXwBv4MSk234kK
bOC2Lrbsgtg+lKJH/toXwF2UqT6sWtrzCbo2RvGhRGNN6uw4eI2ZJE/WnnVV4U9s
GOlAZR8kuqug10H1P9BeRrawHv7ibxP4pYeFZhV2woNX7mOeIN0L4QffEJhFFyXM
fSjePEG/vvaC/msK8KuOqs+vJtXLxrQ+7KlQF+Dyu81nhlqsx+bqSQrYnJMmfEEx
NbXRhv5838YKAQV3Xz3yBbXP2lc/fcphRUMcgg19YsjzeiATdT3IuRUyVMZVDOLw
P540iiJ0b1Td0LO/kwdZNzifnSieWU8UXS8nTQ2XoAhja5e2fd/rX/e72iQDvBOr
gjjkrMYN5uVe26XChZfTTWlPRpHogNuP7Cjzpz2UgoNSQ8DGMSR96H7LTaD3i0DX
NU2PBkEyUf6kogQ1qIwzOXkQ5Gi7UqPEEZVczm2fsKEZnA1w4lHtjX4v40YcH5Et
79afU2caVcikVH1Z+W8LHMxqPNVpkza302EehauNWOME9nbDx2Vosv/I4GL+porI
U4Qvnie1pK+2n7FkVC++Ctt5vcMtyG/FM+aZ/6z3R3ZKb85Til76mU8T7l9UdfwZ
ueeSxEg9zsKun0ZuEgI20dhJYI2GzeiMep0tuKTijOdAa0e1XPV9YIbx8Idx8d8j
sx+vjc/96p3BHP6cV+8Fdvqg+PMpU+McQgYgN3czMxxPIiXzfqxnAvK+a0dJhBk5
BAkaJmz/cmjN4E7hqZkwA3lthh00gyeVrOgmNz0QUaYuUeDjRBLAPLI89oMz5mTo
qxARv2ddpQWr9kYPvXJNQSopfijfuvzOxNgbRS3cWD9kULq6JWRfZ9zhVpNOul6V
RqD5Wj8UvDCJBdixbk6OXgNxKMod/4XfHCCeL4jbIvXSrqM3dAImknddtXqhYfmp
kAvQJVqZODfdXIHKpWJBg641pvXaqK0T/MVzQ6nSJT3w+mlf6N+uK6sRvqsR426E
83S8r4IkPMLPUyo0iptfdWqhdRrAEbxk80Nz+rfv8Ly0XSBF5dRQf+0x9gIri1wC
Q6pmbwtYydtP8E3zIAMIQSQFlEfvuib4FjUhYxsaJGYD4iPT0jswM6BCFfWG1sr4
qypKDVypkjHsDNodkZMaNOkAfK044bTG2XrMI+pz8MnTB56AUw94rLwZG+kewf/o
/0e/w3kVITh3lELW60amUmLxSIMV5+Pyb5hsR92+I1Bh0n2g2BrHvLyHoDF9i4lW
C5nKYUtDLtBKt181WNCm1tra6kL9NSQsatQqvxIAeZMkP6nH450Lj3IubVMpUwq+
9bHfgnY4bnaAnS47DFzbaALSJOfBUpuhB9fgdkTRVteWZQZeWhnBOBJo2SlP1VkN
DukoxeT5ozkeqnPEBPzFnk/SQk9fMJGVy8owEhEf7sDizl8gHu/Z1LCtab05WlR1
NlgQ+oBVuvJ8IOB9l6CJ/Tp/mphnpk3s0Me8gqL1QLN8RKvGEJUAo6odLNSangoM
MArjLd7sldsIgju1dbdRGY7KjKyw+YgmrGJ8MDF0A3ogsvXnngJ5cyK6HyNPJ2W1
qEOcxDahSgkIMUsvt54eWX61bFFtKTRrh2K19wq06qdXQm4QHyp2rH4Vm/mUeJ6z
JwXsXxQfXL6I2ZzYAyKxtYt7bFxxSbXWrHpCxt1TBoc9ou9TyDGQFzD+42IbJY+D
pQg4FTgIxlejE3G64QJnNei838Q4Od3VexE6dC/p23L7DyIcr9DnlpUPMfJPxnya
uLTs8nGp/onFTBZ1cwNECrn213gQ+n74MuDztAqjRX9UaNrm3NOv2mhLxjk+wNhs
YmQmi9BgwTQiIaeXZRcA9nOJtrtnZ0bi+6A1f1BTWQi8ylHG42cid40n7tJES3SX
u1bDvVfe3xlU73sU9/gCZXV7yYqXcZGFNBURCY8USjebJlMkhmtD+dfTPododqkh
0/UYATRT2ZhVZKd/Si0yh+R8/LHmHyAVwsu330keBigKYSxJoaLxyZ2afqExxAdy
GaWOcxhBA31ED5y7kcPd9SFCsSB1cSEp9KRPjIsL9LShwCg4ciqb2lQSYhzaKnpx
Pnx7CONNgCLW1HxMiH4PlJYHHsqbc2+MiNFzWxKhiCv4El0wlVvDOk6j62oz9ei7
bdavqoE2UEHSS6mxPqinA2PB5D19MaYWRZeFXoaJ6QmSJUvC9lzxfk9Nm7yL+JhW
naNddOrEoyE4B6wfleaUKSfLRJKPqpgY0peeXAVQ8/D7jjhQkMQtNvISJnhJMTNd
01cQedFqgtLmC71pqA97D6RSCQl9uI6sb+0pW2uX3MGd2FdMpNev4s4/przWozd9
IznqiBerhFFwUu5S8FVPq3QmupRV9ZxLQSUD6BaYTZPSZD/HJgrUsa1eh/lImAXX
PUrLHGDFx8Mjji+1+U7jPJGVYTI4zLmU6F3R3qufBEq61Cpg8SObeHn3egY5gOa/
sKzr+fwMDxJbKGpq91f+v+qW6+IUdCboOQbvJUH7NFAx0wQlTOWJC+nG/78o1JnS
lma9Vl/ZLRzGoT6Pm6VCRUsyrkkz7TxLI/DQe7bhb3UID91DjR0R3HwaF0cWt1X2
Kth3t9VEs2Vg8cW1s3SB60UvTnKtE+DkgewMcQduXa4LsI8O8hHg1rBZzlWJFu18
QYRxMCITse9KgDlm+lWuvEjkCkAAZXXl/7nVWACXg2t2ShFZRYcGwScyN5sh8j3G
6KClFCr5f37D1a4SBsb3Bh34Mf7znap/Lq3y3VJ5Gw5scFoSipKGlaKE/5v1eTl8
deXVK+RJX1YrEx9isbV+d8taBczp7inWyBVm/0b9uqKsz4lZAcw8Urb/Oi9zihVh
UBptum83ZdVFNEum10D1wVL6jZTRPN6R0VJqIgM2rqSPjUWYHkRyvFFjtViMUyQH
XMp7MnwZORk/AZDqaMbtt5v0EsMkwoBPU4bkG6AUbtic/PeFyPVq2ut1viiKB2fG
/Y49azKhgx0I5d+PHJemmI8JUZ0ghI/kYfojNcVMb2F6H3FT3BaKpZIa3ZbzvfBI
nF6LvKWwrPysNU1QVsgD0quUnXfG7jObMjY06WK17yfaF1RuhPv65Oy0/iBuAZpL
zCIjhbFyURPH2ZHwUNlpGhDGw00v3++UF0UAijNMZ/+lYD/YJXaMXdAFQP83PbiK
A0NJtHB1FPq07kM4pC0JLxYN+CtX3j8lIyPHwK4jpfHMRFzvDomRTYSDuSDfgkNl
pbYJddLi+QABK8dKEZFux+vAYu7KVbdjQnPo/oWFYOgFEAkFldjClEZCViPEzRa8
lkjnMcX/bOqVfBcR7qyDnAhmXBW8+ho6yzMPtnjCOjFUW/m8nqvDB3GWYvd9Nb77
SSyopocR9xNW30W8Umg/c8cE3vOSZQUa4D7kpZwRHaYXFsDmsYqV0CPiOEYoQ1Ti
FktEN2D8wEUVHfi5jCNzRojOfJIpR40sLl8AZKKRzp/uXgQi8Kzc8j7rez3B3fpD
vVwmfhE14bu5tq6HCQ8h+kzMsLz2iZugTI/ZhxT3uXRbEhNUsiilBuppQ35fX4s7
gq6FHbJmCq6wBGndtBp1tdkn5t9CgU4VNuEb0k+ivzsjMCoRaDTnMsxhkTW1cgH+
K603Gy91ktCMNEG/XrvdSi5GKwaKP0RrXVm53L2J85KoyYh0VPOHbmDUfVvP3xBT
vHvo1NxiCcxtuVUaHpZEmLjmC1cr4OPX5YilDOBK592izXyhNQYDsrlBrpZlCPU0
fdexv6doG/hC6ORca25qEAtIK7zoPowVCdabtNa0ZqZRqhwMtRoT1Kl7JcUAgppT
zPimrcZ5UsVyuPV8ZPCm3sFVjI2FP+HEACrcyaASnbGHu1GitrouvYcFUWuygvmF
Yy6T7jEmHbtJSrHCC5jGlPi8LSzg+xT73wZZkP/j7Q5Vs4OANry8+wAWs8j9zggN
QS9tGcgg/m1BEu9rCzvBfS5e2CNz7OFhoSSjFS9NCsWS7P5H0uTgiCBUEP8kXlRV
LWbqIRFV3l1c480u44fKO+b9s91SU/EW6/+co4kmM/wyFJT1YzOV6IxsuKzmNyLu
oGAmh9UATlRbnQ07894ESFDlQnJYQyCN/JUUOwhLS3GNLMQ7oC5QSpwChsYK9TqJ
E9UlhjPDWCGIea3woWzXlQfTeVEoVnbUSUcAiUYS4JWTclU1eFwijs8GZSQ0YPx1
J0Ig4eXbkGfAtqawJBD/gPzL2Dx7X5PdmG3foEMVAFnNjQ/+arwXOdsrERotghmk
0PT3gQnArbE+6HfOGFQBDEHM5DE+XhJ+YCHEQ5PLbT7RauDvDu83MlVphyQsasvj
zXE8UxmBSq+ndAEXVMVStyGiidRdCoPET/w1zltwRNTqu0vppxigiSHbBDtXw52R
N7eRnDoycouBs1Dsnv1jgDiuXp1RDDGMSnFt6VGqJmN12qSkCx+IhIqfyisPYcVz
NA3QrnD/ZG3lNXxQGYtfl92rZioLzkycvN9hCWsaMCjbRPdSNrGx9xtIfTh4ZHDZ
UoqSVo/87Bs1cjdkXDLNgqmW8uTmmFbvlu62yZjILLulfius5eqp1w5OJSfsPt7w
ZaJcdMYtiyFXeuu3OEy+wYdHCv70jh2r5tt/9BnuNtkGIl7kh6QSr+v7CIoS4hy6
hQhfwyuRjf70xhlyHx+G2yIGb2eA3RuZyhq8ga+S+YAGpRd0okh/+Vg5Cf6/OTgq
4TAFN7PPLg3ScqqWwXXPOQrQD6UhHZguyEowCm8jVHh8KW7TWDvF3sOD37GMQ/fY
AztqmTfknMeddbheSwqwAAQRYYjv6BwWtxMFPtvRn3BOA3RK+SBkMwwNUxFODUik
eNql1T4nfKIcEyjbH3A96oJCn/0MppvH4zQt+/11XEug5LIocqmmEK1WHaeD3KcC
qLggGXgYqSqyjZR1msdJpneapXHpYer9RQq9b57YPzIsBwJTA0f0qvvrf1UW0vfk
F+HSiuWcTxsPcmn+KbYRj0LJtwjxkj6h8JpLbXCzMTFkER5kFxRLm+i8vlx3ka/n
rUbBu8EJLJ/siFdnooZJpnni9i9SZNXtQcukieUKdAJ0x1kqqqwHMzvisrjw1mmI
K96/WNtxF1Dq1nLiQDu8oibXwlHLN06yQfx3Z2baMPLJLV/jvCQVvRqzreemXgTE
FrcFrxUAFiYgi/cZQfhQ41l9LXyyfC9zdoxbStAQsgn0ULLVgFGYOhu2R/uXD8mt
Ilbn6pmMIo0lryKhlCp8d1D1o0DCPm9ZRWLtnki57lDByTEsEIiPAnBrEaAZ65Qq
P3/KhgSO7LlU8EB7yzhRmL6knfXA70eIVcgGAfgUvbtVGh8emQjaTsgEXnBw7y47
1WcSjjojibrEby2jxu4iwBLMw1kiLnityozk2QT3A8V62V2hW58CwUkEJB89Q/vM
y1fg/8MRY5bzH8Vz5oCZENMFyaavnGUkPPHtn1W3lY9cOAGiKWmt2OYI/xhhdiu+
3ryAMWrjboVun7JbOwr03ARKynAzE/f+uZ+/agfm7Ot8ac7YhsJ5iZWHd13gwe0A
twGcrxXTRSPZhmPE3NelFvSklHn6D2e/CpAIfCvHAMTQGfQLeOH4U7Nt2NDgXYel
pDWwH7GwT1FWiM/cM21H1bOMpRv3tlsVmBPDhWLjtOs3fPTk9DVy28PdcbjNtuZM
CIfOdv/QW+tTxlHjRYAsJZ74SeAS85vfx9cWta7ctZtdaoOKWWrYirniIeKQx93j
o7hXvYElzC5RJy+hDw28U82plvl08yr2SdjUw9lYod0AR9konIgDRJIJBiWTzTWD
plhAqdPHA38bLbenBcdckYF2JgXPNv39jolwsBs0RShOjLmExmVTblzM09wDCyUr
qqONz7AodHsKRWYsVj5K5umjKI1rbw2u0hZ+eqHPoBoNyBP4dlWyA8OBynZGONio
DcudvCZL9TXKBi+N/UB0z1Qqrnclrz1jRDaUBh4issPKI+HAxRg6Wr+DmzoXhYFA
RHfdkcsU18o4myGZNCR6GKZoxBF9/LJN7MBatgjdMcuzkl2nhaGJaPU07x28NPFp
uzWtuIPmJ+j5nF51Fhcpt965nhRnfnOGEeFADpYJIzmwSuSprRdJixL3AK2i5sLh
DXfvGvPVChyTKzR71UgvzK/s3B4MQCx40/V8nARUdvMU5WxJmLYZXq3m5DwBguFN
yIgDu6fRqVPr00hmBOAYjWQ5V7leFzbaylOWnr2ofI/XwQuPMQxVhBxV5LnpZF3f
27UgM2i40ZZ7p8HzhIbGYprYNEYBwnjF1/eI6B+GyoOkKrn+NDnB+YjajZgREuGS
MEj7nHumVXMDEJoUWSvD7/GeSBNAqZA9GOT+7PhsvzmKDmF1QqhPmHJ0gBcHHLtA
ChNjw7ous/ufVvEgdqbRimMD6lBA59DOiG9Krgt6aidDDcuFJgGTiv+F+7E3IBb7
4DWytNG86uaUdbLrtbU2zd4sSmIuvAF5fUp2+n3oh43RqOzGjA5QRQ0jvzA6RZfi
IM/uqCgYJ+q2Dhd4LZ1wLdKUDWWh1RovfMyooxbYTmvpU3Kryhm7WkI4OIgflLLz
tVbCWyG43xHpcVCcPlev+HkJDVLu5alKE6mGtbt8CvHnxfs5qAHRTKhpfiQ9zd/i
2B2neUWjvItZZPTIR0mjpmbisf5JCm4BcjzRwnESZ4DiwTWMXR82EpbG5Cws8reB
NTGBKiXPzCammqXIiedHM6YAhJCOp0NaL7476Y72zDNPwDzyFlQCAH5g8i75o7Qy
9JOLlXLyzuC1gKHD0cG7ZVy5LyUvN35tfLwYhSdm8SxgJb/JHSJomh15yP5qO0sq
cjAUCbNLs+RmvhRsJhEIBzqoDKxj45amTly+TrV48hGIWKGcT9ZQrazQaNk3k2KD
nznlC4Rc4CCkzefp/AFXq8ZJ+N3zE5woQrqcumJh5+ZrUemIuYCu5Ah5EUedEH9P
pSwIg9hCs8ZkuZA+N3eQ89e6pqpWFcm1/w3pV0y2aRT5lR5KQahNR0koWRr4MJRC
WMYdST32wbhydShQt5noURwVhhEv9k2K5z5/4MGrkOHOyKyzo4hJ5pqisxyhXB2F
VYFs/AWNBycGTq3Hw8mRsw4bnTg9QdbKuhye3a3TxvxE/9x4881CYFSvs6mt15p8
WPNNqGZlKX3nGcwtw8qtFs2lqrufTqzRmlh9dl4bj+ib11IJWGzDczmrhGfwzXqB
qcgvRoauCb8B7gD2VyI0ST+pCEVnO1NJHO2efKRhfjXnSetiXULpbCp9ULE9DSWH
wB+p5jNP+n4/y+W+00UMpcw3/nXYOFO7wH9HJ6nOvinafwaYSLQoJ7gT9NCmS+XU
qEMdmocGAQ3s+pwm//G/dr9v/Gal9QkCYujELO3zknhkfC/kJp/elGmAF70JOVia
jLnr5meaSmFxg6BVTjYuBXp4UB8J64tdUSMWf4DDZknsSCQvjbqc/TfrbTBtmG5Q
3T9KD3jcOwFAC/DWBS/yHemhQpWYswrsnGBtgYFFVGTnr8NjfSS6ZU5h7tmMpV+v
H/Fx9PIwx9VmwLuR48LD4uKsN2KWtm9C6KSHX/h1ptdVRHZxKdNqtL8oysYTePcO
xB4jU7pAuIx9PI0ylZ0cTrN0nogRYTzczIObh0FNYcioDRw3vmsrLu4xg/UPEYaZ
W/NUmE1fwrjPN27FdgfVAKaoaqV/tsWMbheNXUlkXf4Wc0tSPenF+7lSgWsy5uWy
zcYgmj8tshH0aNEvHzQuUMmKAklEEHj8tWOvKcPkj1YHjnXiSueF/f8SIL3S7q+T
nEl6ieoa0bR0Yivu2svZVXwayZlY3MFfAmzVbcCVxhppUWniE2cmu1+a9mymCSOZ
Z1tBjPMLyt+yZR2oFCh+OTidHoyw02FW+Gjo6Qsuca+UdkHZbGv501aqlTUumon7
8k/gPQeXDAI6ewfZjL1B9Nm2hob2m+wnfxnnteQqhUJcmQmVinOqEQ2RZusZ/ige
YPAszWl8juM1u4dtzqnjsM4TiaUENEelGBk+Vs0Rj7vgzCfI5LM8RJt+NBLJhe+l
m6wt/3SdmIAcI35QIbrbYb9ZLIy70UP4EcQyFsCsLLq9JqUfz3F9QpNL16Ymww9x
YsbfoEJNusqbku3q0H6yoc/HuMuzm3m3Oz2d6dbqPmSiKOj0aH49N4obb/uYwv1/
/7HmtR9rlWs71Q66uo27I8v96LeKTTLShuVjItG9Ib+Jv6wXcM4ZaK4NkXpDvY/Y
JmEcZBoJN49WXfWqKSlozbO/h5B0ZsbEyJeSspR+48o97nF1YdZ2UFBn6V2I+E6P
xhRfFZTb+A+B5qomF0G56f7XP+5Io8L2QvUzuKlug5lV53+nKAUDV5Q0GxCXgCw/
5+qXEMF1Mzs38nKjFIkRMPeRfCHUd46t2JC+Ngme4u29CI00ET4IQ66fd2JNPVgh
iLeOFNE1Tg9ilFB/TpRFt98w9ofN1uBQ7yTbAgydPzTrtpnGG187QUdWWpc/jE7T
Xr5BEUKGKP5G4FR9CaNocYr3+oX4cSV4laus9kAPXOtmRioW7D3xwa0fiO+Dn9GK
+wIbJVFMrAqEDSd6NhDYgq+p08N+N97w6KP9bJBPWJyArMekfDEEVgIlV2awwRn9
VRDr0DykSyvsKMqdof5PaeJ4pWR0KBlrgrr1GxKE48x4ystq6clSb27ErfC1vgYh
c8knBxGWsup5HnLXYWaOGE8QtQMjnuKsPp4AW9pJDwDbnLzsRmyo3eA31FN6n46p
74fg1d7io4sIS+MzCUfvgKsMZPBnuSWyyK+8OWmiCK7oADKo4KOVNR7/gsaPTShs
ykeiyKBqoqzt5WwyQTgxWvmoZNkRxncLl3SRVWrkHE/tsdl/dTZv5L6ZMp2PYi0A
fr1ofGuUoR42kA87mf8FUN64eU0DR8+8ATZvYyto5FDOsjlbh5UOGrI3jzRrUYTT
/XsXyMvxUfqICfu9XHm//HBsaPk0dDP2CJ1cjz9LEBo/urwQQTr7V0IdU9UT+QIJ
gdyAGNyllRVOKs5p9p0ny996VHufTbUrpEp2O728CHGHH+5aSaoR26KbWMaDyHD3
LWRFs+39ccgwMbI8UQ4pvY9UCTz1AT8VdmfnPyPYeyRgFxJ348Vwe4iUCKDD4nWv
9NoDWZAfkMxVFf00XcfI3X/VpjLgRkZkX1lFHvIAq91Ib7z4eOAJqzCISgOyxaYZ
o+qTktRbe0QqWGjXWvRvuT7kMs0SqNjMiAuMCo1ZhZxvH8tEJvW9CGlWfx4aJdmc
OwE4CnNuKfhOIllpCLbip6j40orM9oFMTvpS9/eB6fr0Pf/F/E1MLLMT83VkVJNJ
UO0zfQ6J1BISjXbsrbX6O2qtRth9JeZHmPQGJLl6GPzbVpbIaHO+bxwcrfE1JhYu
ZdFN8ktc1dMwuDZcv8ghrRMlsUVleOo9mvC2nzCSMKH8H+BS6LRivtu3KnqaGiyu
51vLtbZLnfScL9gNVf2YqgpaLwFhfFNOteSQOH9synMavUX0kpJjmYNWgd4wHazQ
40nwgKhNk8y5ay8XKMAwGJgYT8MqKjl40F2bT7DY2t0anLXZxJg+BltAX46mcsb4
QOTe1YcUrRFfItfkqi7dq/WM8s2nXgqZQ9YBNdiJ8vxu2tWBoHo7mXMQFm5MUxU9
LJzYM6sJ6JkS19bApbHct/17xxyuh65vH4odbTlkgHcFPaZXa9LPznC9M/Svk4ty
w9eYlf14ChZRxbnsILTDhbEor3zmfikXMzcQpbQBbaj3umPmQ5r1eTPLQ9ub70Jv
c9NXY7QgRW8hmQwsWUdCQiuzFW3OFPyX+BSYSZmQF8E0Z7zfHmp+9lLylLOM9UwY
ZDayPOtB3hHIKOvFmK8X3gklX3DYhGr71aSoKg7j4rUWftJ/3Ckmwt9JUJhAqzsl
QhCHPVRP7XI/mPMNy7am1f61JUr2XlfLtMR7eO8BTSQPdNp8L0zjo3OMNTsQvZjv
YleqGWUQ2Lz86eOYXajA/YztUVptwveaYdzWFS5E8MXRnQxdU/eOw2rBB+jp9QPr
PHxLL2IRVWteng0PINUC0BJUlVNF3EJlhLTyUieE7rp2uSBSwjGvXVKE/Lu0W4Dn
YYJbc3EBqGx/fmGrWe3CwWWgO8I7EuqHCr0V4Ku+DNJnGA7C/wT2qGKRScw6hhHw
u29FDZwMIMTd0e/HZpqfnMLWNxdb+JC9VX0Act79glF3kaFviCzuOUPmi598/Xvr
xHW6QD5h5sO2BMT30qmbu98P4vxdoHTjE5WgzEWUBJakbwpWXsS5Ouv9TlbB/X+d
m7H73FRoW7BQMswVqJWSl+ENH4FsMb0WpSy14DpfNUlGkn9myG9+f8l7Atfc55Ub
I1ljSnEc/EfEieEvcZl9vC1T4a2xzjEd20e6wMRocv18Zee4XSS34AxFIWZSamNV
whm9z/X6MiNuGEQU8e09dG7x0opjQvQ+0bYci+7w2QlZoqS+rlHXJpQqbU5tELMq
lfZ0d3A9vKk02x/Z58c1TlMPIoRhBCnLulPpa6Ec/veZ42l05LzaPzMkGylAzk0+
pDx6fcML6ZmE8XPDmCXWimOCfbHTSlWuT1mXRkoyQo35rGxRyMaF0ETP4fqK7MH9
+uC3p03t/OpvbAOBUAXv47higfdZkRBf8kCJKicJ2cJqNkTL2EISrJXBJbnSLs1t
9HRH8IgJCFQmtjNOtI7Grfyl3UtfgX8h2Zdw33MR4EZ0ZuS8eOCJgL7oYFASBC/I
z+M1yfu6u9t31N+EWDiV4qnWp7n2UcfTWRnUsKUCFzV/3C+PPMmhoPDddEXjTEsT
TpETHaCX8VDWRPx1fr+aIcBC6EssAdfrxI6Jk0FUWxcrJmZfeL0LJQKrqcnVvmiB
1HRxUOovf/Q0dJHeooE3MrcemxCj2x1KlycttzNxPdYY94YPg7mtQchgbNIE3yrP
Fx82MKgHKWGO/D2Lnm59rst5Cp3gd8aLysvE5SdW7u5yRugWIUDstVikTSVQvi/i
q/+BZspMnQX5wxXnHMCYUgZsTnyq7XEAb30PAX+t3WRID8HivfHfPZZk6FBvnU0E
s++J7B6OhDvXsPxVr68tvl5mEA66lum/ZK/IXDaFUiM+PbVjeb3O+lAJgpKYqNvn
sSk2pmOxs8s7tSriNhDUrtoOdpeBUEvfYPXz2MbiyYw4QYdsVYlO4dV9atwwehrb
1sBXRE/ISlrHA4WIgTyqmDxxsKO2UvDIFtMAk8bbnHd91M05yUSbzxaNMT/BScbq
ScrTaJ0Ut8Z6bMHgQTTRNI+P9gVJS8EtPS23HDml//A0Pyu89iE8lnXPDEqqAQ0t
fQuS2JLzDsyb3hZn7rU9a/k5tFfYQweQxx6dhwaOcbeYhKsQhhYbu1gpTMHRCYjh
GIc2YIONfXH16/LlbWaXyAG4Jt6aA5fr90n99uTenQxFpxeQaVsabayxEryliAJc
gF+xJTvtRmR0yQqcpf2QGFRaFweXd5e925+puWCyfTmi7l49Ize2C15yy3Hzwt/t
EoimVwUX1F2LZTXfHfZCLOwBcsi2MBdiUPcVv8K3FysNEaVEpgUF7eUe0LpEkAfJ
RbMrJVVRfvHsMgIV6J/jeTLkzhSZM4OUDvvIPZnLAdIY5rNE7NfjCvz7T5OrFLHh
n++fs+n40LsIFQLi8cNPTX1KkELf+LOsz6NYTPKVvd2Fdu/gBXVYqakUXupKeKlo
nC1+OsBZKL00BKfBeu8eIX7AeXC029vGDwQzBPNAe5XV3vMVoFYEE6ZdyJU7JHgp
LQpRyvpZbNIgUx6YyeW6OPOEf3OJCPnyPLNOekgqKEv/l7ra+LrEW/2Gcphy6Rrg
Tz3jVSDzmdagD92gy+k0VfG0ntwTKP8DYIHBGS16QYqizFCtW5afnNrFsC4/8XIo
7Hun8PznX+KENsj8RfmHKPRAcQFfng0s9C/Gvm3yR0VtIyxPU4OMTi0BIsZoPhTF
gBRhD6i09LLPoa2L9S3kDLBoGSvMZnRvnfWWhwEF7bHse28CFSjaomlMyM5ddLtn
j96KkMbmU4Yb6Mi+p8JXjNLNHa6UIQaZHD+IrIV/7ReDNkOpKM9H5qfnPw8XuGuh
Bvo3GKGaeaj/gAmlet0Ro/XOlBsIcQTEgLHgE6xzlAMK3qrWDXdOPslvKWfnDwFC
2MqTbuXlXjVlZ3oK+WvwK5LPCZWJvXb4wSrPahHzvbPhXuh743RGtNnuQBQe/sFL
bEOnFsSzM1Y9WrC65O5Ki4OrRUyr/YARa0jZRpBCaMyR2ppSO2MTt3eI2kWhhujn
PSABVZtE7M7jq0M4xoU+airMss8k4x9de4JdTZByvJr+E9r5EXGBBxdRSj14GzPg
Lkp5Jf0rvTK/6z0ZPEckqNqDVEF+DARyGIZ1L1yW3KXpwO9zeAm0PKUo8ufLIVGU
MKHMWiabmqcgrItP4vL291IP8kUk2B6ywe9QOIlmaM7HyTBZdRDebUR9lgsC1kQN
oiBgUI9NvCY3a8dUbzgPYxLgck3XaZxSgfv2WPWE4LgvtiCNwBDo7eTTvJvRKLwH
4U+Lmc65OxkTGrTxuetYZLmDyvwTjUNkuKuISDWlP9E6W20v9Iyoubx1Zjd20Z6y
jaiIgq3UgC/pI415Brq0gbZPc97mbfqnktIBDbofO6o9U5IyyRFwba3BBY7DJtou
VuyVN5EFSQfMzhzLwET3Ac9EaH5nyWGbpszO/vRrf/CC915mIwSNx4brvLWzPSIB
b4t5+7e+brm5mb0Fm81aJ1dvyF1x429W90+UDrZa5I5HUH8RYbkPiV+sjjJtikoV
9UK9D2UhQp9dhk2hXTkwTUON1G0v/nVoOgXd4gTxXRiMvlCuFw+2l2hgzeBvVvQD
yDcQB2xGQcL8LoUVnPqIxl41T7sdpmZLxqwMiTxjcXHmniZkBs1T9Zu8tYOySLTn
IQlV/eSWiCS0z9+j4yYz43FxnXcKmIZnHhDEHrGRlLtOoWElpzU0ZWaWmQEYpqd/
qIx8RzZZhxlPBm0hYm8v+Y/G5C8TFy29ie6hZAYsqmwp//PU/9YnagSCFz3xT+Ik
uBBzv9DtpF9GKLeH1e5llI82ySzuvnEXvE1sm68q+gzOgdijaJDwCyPWxxVaveuW
4SE1BwPJgQExNd9GjFbctVCuvKqrm0nug0WMYP1ql+RRvh+4PjBHcxy3YPmN+zX4
LxNM4/9j49/T4RuuZxtZwaF5JR2hgpmXYP+Phiu+GM5eqYzZWCldUP3IOoWEHJz2
6kqEe+81cDTqquzE6Pa2wkd7wTHUK/2GlyA4vtHGDogycG+WjBIfCg4UZ8wUUBWw
gnPagOEfpoTRVp9HZLQo6VkJ7ktUGAH8pRnzInTRGcIc0UJ4Q4FN2qgjfeMQAQTC
ng6RNByU5R2uj8kRdl2tni34zJl9comfZsqeHjo8QXHWMblKMggPw5WI37e4kMli
1hTL6gdTIWJAH5j5jZoRVTdjiN8wqD1VID7pIsku7ynLGXgsOPA7PeaXs7Y2pf02
dFaLYluLpgeblw3FKb80ksogW/i9NetvZCjdKvRQO7kVpTkj/c5gKsZ899yL8vBZ
O4VjGlCkctYael6rHj7lWQz/K/uXCA44PHPh8DLANS4xc9rWXsao1mjCxNeySO1p
IU2M0EtN2nkGYF+gmlo6DVBluQeBQ4+M6E0MF3Sn/kaMt4EVHC6FYsGJsxxg/ThK
ovGbo9e5rkBXC438bbHXyCAK7uOjX0hSTTMZW64y2sMIpjZ9+10qNW+iQWqU3gZk
lqBl3ThlwudqDs+qVaA1L1ie5cWRwss6pfmbWlBKLVmjcYAp14Mnh6QeZwwWTCFA
XRjRLinlyY1JAxjLFiRdxPVA2c/5S0RRWEx8DaESivt446szDLDl3G9NtHQqQ+HC
dGbx0Fn37ugOrH6jpSFVSVgayROLUFTGv+i5dSznSCFgJwEBNoyzfmPwzuTIJd5o
xM+mSoXVTAoyVg05Cqb/imPYf/ybVv9vkabFBR9flFQzm5xtXH3VBYq4khzZjdSP
NWyWUwlYFR7b48fSKYIk8ocs+sNaeh+8yMNdQDDjWfZccprbeYmVfjkblzjUqJrW
rXsnF3uIhaWUc15bWFvHTG3eAVslnpE/mAmsOLIN8pairM+nL+MZkOZxV9PXD9ux
qRFKdKsyx2hjD0Teu4O1orbhZOJZojtQdYu7HgiC7ReutLYReJ5l6YBQJVqiJz4y
D79cRjvzPh5ganEDs22d+YFSjSD2cJY5vJ7cMHg4ClYtP3VAgIuDrhNfevL+2mdU
aMGOugLU4C1MyqFqycX9NO+XlPelHqfLsAdh6ew6buntxRAawr81sPV00s1T0Q+e
BgQ49JjA4iGlEF4eukqr21Tn2qQxstcsc75bDuCP/WOJl/YPDWg9Y/nyzlLSX0CY
vInzmYpGtCmef33S7RRq2FFkprCGhSDXL2ZCVNhjuVSpPx3E7+Fri729apJbw4zb
nTpv/77a/5XzxY8Ahkq5qFomAihp+C9mheQY1bmMrYU3WolYKeVzX7XO4xeJm/ql
CwUQT+ZsQ8+YC6aDUo5ASrkvnwa0gDNET4unY0OVKrwLT3cPEPZA1La9Kd61Cpiz
m2iGkL9cXCUx5M+vYtsnbsTMg8Ud3bH5yuIasuVtNQSAXFKpW13DGKl1TMWR8W+c
sXyOAi5LojzYLdEyEI0EOh/DOX+kpnHzH7Dr5xcZaOUAe6gCvKSzkpVC2h7OQAy8
hy/e8O2MF95BeQlKO/POdMSZmCkyRRR9R7g6Mfx08pmjtRCCLC3id70OMw/Lz6MS
j/F1Z6j4Wc9uo5U74HpD+iILeKxJ3SxNofYKBuuBFhMnBHGYLnvoZcFPyp+1cQhy
gmg+eGaPgERiZkH+F/pr3J1TZrMzu7jnyRTeu/CWjQHLcS2HBYKmkcAZUFZVykM1
CDQR1G2sPkOM6g+vhEKnOOYCvyQIBGAP4yvdVc8FUHE3wQuM0w2NAatfu4x+JmVE
ckRkYomcPFJS9WLg51XLPyj7SLfkdISQjmaUK2KHi5B2gEAkQlh1cqZX2OBlCA4g
rTtjOQC+efwxuz4cIhiY3/8ri3nKqCu9/xll+OplsUW8MZam2kIhwzdiVlEtNDck
DrpD5OkafO0y+AvPhHxurtxrtrSqhCVCMK8vWYspq82L4CBZJx2olgwYEhsVvsFb
M6c9Co0Hwc3J2zWDwQlYstwXpLEnuaCVqey1kv3/wQ8TUSXlyNaRf2iiS6FlbpuI
L8IUXoN+MiGRn4otDbwjYszuG+VryxsGK8XtyfI6LeWZCX/SzrrcURYHAAAEAGB8
bvKN7dHkyNBezbwAaSC5IjyyozEWx2Ft14gjxoAiEqz2BKDQxt97GKL4SKkI6BSk
HBPlIQihT0vMvc9Syn1C30O/KxAgHkJeMLX+v5G9rgGb30ow7YlOTDdaO36wCrNQ
GLbX83K1tGAT12FAkzSJlB8cvOdAGbBGGQOBfecHBXVhCBZANbcM739FEJYWBZGc
xKa9Tfpi/XPCOaqaVsZxXGcWuFrdU+YdAVPf2Vz02I89nIko6SAgt/cbJcl4jmua
A0xOKQjcG/7zJ/7Mc1Kj7nRKJ0L9OITdXqX7oedccGa37Cj0Rn0mstrB7nCknp2a
jjSPd7TGacFMJk0w6x0Kql6QkqR9N5sDg7UJGf/cV2YT1J74kq+2IGjD0K+Ot+pc
Kk6wVlUqpiZfylj33rjSGM1IJM3I8p1kqCbjf1a2g9zekCNAy8CLAs4tK3jx27CZ
8xwO+rAQhu+C0yD7yNXCQNq+JHm0ANoJOJdVGPC8dkNIo93BqFsw1mowoqWAnNUi
gqkPanuHte41fNyGG/wHYYvvVN6NKrHe3Kkbn4x7Mn9M7t+zsPgTdwrAJLhJcQmr
F2wQchyZpMBt48DLXPPc+bHXkZu+oQ2fjFasUKHjYbcaGpvR2iuJdDN1QX65fXRy
5OQeJqmRvtZ5UH63rlCNc/8LvirWl6B9loscSCYin45Nw5hQyFdXD4vDHcaCHrRo
GYaVwbII1hxYlqUbsudYTUSsjg+kNdrJaZAhLkfVuSY32TJdvFTrvnv0Y/2eDh26
NCsPrc9kFU6qW8hX46HMPyeyzw0WgUuZeX2CTI50XjIeuup/6EKC1nLIth/soc1F
MM3W1tvPOj+cYyi83NLEfq6It7DfnDe0yfugq1KBuE5cRfeD7LezIJH+0ht8EqB8
pIQVWcUSj7lRPq2RZ+w6o6jO9x8Ie3KZYTlkw+9aX0ERajNVvcGIUVfY7/CsT7NN
vdPthsm7XLQIhzlhLWAsNo0MaIAQS8v/BR9sv/0dcNLluHXkyT6LnQ4AzA0du/QP
wS/YZNgJi1Y158sn4fE8AOCKFyeVvSfMHvtzIjc9Qo0fT27iymYqwe/gIHPp5XLk
9MH1o/ZP42RzcOvq5iDYEtkRuLBSMYsXzJRc92i/vjpkxICasWPyo0ocSxDCQKfl
NkIaPJTBk5hZ65c1oeWJNxt90S2B9gjYikitYG3hN59GYCh1ctlDby52txo7qExQ
oIximMR0DT224HMOuBQFVSNIFDnhVxLP8dqlrjj1Ipbi4zyiqSkq4JcI7iTsDYV8
aNP8WXfCRm0mu/MBIJxdS5Cp73FLY/TeVLB+0NSDrniIv4OXqtFyP33FzrUKV/Y7
N/NLhTGjrH2oiLZFMe3HKbK9s3ttr2LTQV3NkSeN7jwnInBpgEsrn+iQ5QNtRehA
75fq0xBXBdxoN6qrSs2hayzmHFWbXJG59Y8PAsn3HwzVRawQ9/szHGFSdtRuIhSP
ldeJEGtT2+BzegZdN097WqjK8Wl3y77rrfRO+NbEF5Ll7s371cZqc9c8m0q54zsb
oq7ltdI+lBZ0qlkUWeM18N14CrdRXhvESERb5l8jGOgePHuyQsBBlxH7eLKWZ6JY
gjVQZhAAx0Y5AV8maFXjIIAB7xiai4Z9nF1H0+TKfu/ynHEUqX7Q3lov2hJbUMJD
n6ZN8/imKCa9LqYZ2Fkd9ErewizUTgmNk0NzjILkVW+1YgQ45A0vU1ZZE/1vyVpe
RN11nhLR/BdELZM1QdFpsXJAD1ixWVG2iuuFPODxgFDleHHp695+DjL9AX+hN95t
+lAWmL46CpuUdykJLnwNI1j1lEiIAsfTI+sB3Mpi4FTMkVMGBmwvpFmP26uZXrCu
gG/TT8dOrEMuWBwQeQOIYZ18YhGIlhH3BthrvRdH7cwZRBFjrDSD91Rr3wkNP7/K
2/51EdrA6Tg41Paw3u6v+y+s0KNKn27FkxKzuZ2yBTYJLpO7iwX/VvBd2CUQhq2w
hVe90nWKW/kz0tZuHZ9e+fFox6Oi5MbqiYqUy67NaG4e7u23D68MlegmA05pTTUT
nH0pdL+nlsA65Gxng78FXpOF5iBbeYhPyQwj/eI3idlkz4G31BW4tQH2xG7SPdx9
cAr//Brq83H7IbkRu4tNPpjsDPn+UPXVHTuPPuNnvBl/LBhwVwQedf7AW0ioLuYr
VeWWxPp+DCsBt3t0HpQ11ue+EbzNYFhtD4/sYSM3KZgwBOSprA/dbx556UyzLZnc
qmuEVfb71DGgmqnPLo8ssnkwT0gDFPxrfvba39Z51KP2l8kem4X/j1dR6a+vZNj/
yByxPPrduRHyKbR9wBg62ozdmHmeIdyASrkpmbji5kj3K2vJg02bMRC2I58Xxlyl
e1JU9hZnFDQKlVD2FJedUbSzVbdrAoZ4wkzhg7rYtEa4vfS6tHxGufOsdjHkU0SU
3+TqFSFDnma/meQXFIvUUJYHh7a3RFuj9KVKa93zQA+CLvQRabAkdNsSl6bHRen8
1oaZrcVlYvzivL0FtggCQJoiNaE7KotoGPGxcQO1MsDI73cBpAWvtVnTWceJ50yv
tS4gA+6V9EB4UyMU9wtfGN9DHRpSgVsreIVVq780MnxD8aurkD0yPlUSOhf2QN5e
PCZ94QtRG+WxMBq7CVAjYIt2/v2wZ3OexuJOmzZtkCA+IfGKXANj6/9gP+kDnyDe
YssUE+lL3TTtc8EDJkrkCgFRJNHONTTRWrw/TA1clQZNAP7uv2ejGa55bfoqsCFc
dBQvtdiMNGYuner234YxLvnKHzHvv+Hpj9YL+EoFAV6GAoQ2sXhr0GgKz7Ha/tMB
fxxw4SMZj+jdSp0Wnew8QCh2ZrwLrinClYXbDMzTfw/N/kxNLXn1Xb7pc/mWmVuv
qIc7OG8TYl8M7iS+Anw3+ITK9ei+xwACqZ5SWkP9WAfhtLtNMZ+GiH+vfsRWDvGd
0XwtJivdzOKimhutwP9m1FA9+XMb6w5TyiOJp5ZU0p92GxvqNXFd1mPvFc52tfL3
OjE3ri3drOGyY7aXWIpq9vx1/MwZTWJu48clEA2kadA8Dny60mqj0tkcVWEWZNmN
zW7YipnaWfYwHF/iMny2Jyh3W3l7Yw7ACaKB4koWTnL5QsuWlIPEraurTuHbEXTr
MsH87b7eGNc7eLpxJpAp4xjiExybLyTxgKYKOMNehi5ZCtzaB6/pOiLJxk96PUQj
brb+m3cXorz15CnzfVdQndTm0PsiBYZolCV7HFD/UGE6Bm8ndm4pqHKyb8fL3UXt
tnyeWzCjYQe2LusOgREG5Qmt3AT51FfRr1uDOwztNl2ym8INo2EEGvlG7aFx3sxa
ogud9mdQttrhZoZLdYVYIZ6MPkY3c0108zgk9zsPXeaV1USY5qM9Zc9DCaBVcSL6
UdJSY2AZpYK5Vp9GoW21uP54g0LQmfCNrMHcPhQswCHIPirQzLHU16yaH+JEuqvT
f+ypIZkUqezpk5+nz75DXEBCuq1xZ9BMt4kXhBSJrmQdW2bDpWyqKhTjAtqCXxQc
6o/MM8gMqSRnOEEdBCHNgy6qe75B4kCTrg6nOyp1uGnqCkg+3FeW6COHXXtlWtZs
eokLk2kbcrbi5ldWJPgvM3h4NdssBmHKcstypJnQBHHH9e3ds7GHTHbgPrKYfo/H
6Q8JiMFYH3q1+GxrJKm+N32MVoNxsYrye2dp1DngtNZo4LmP7BNoMaJGlF0A7RFr
aZkMNkcMynNgJm5K6su4Dl0t7uoFhllcS6Im2P9GhW9cj/PnR12nwASbGVJgySvq
WstOrCvXth6GRpkNfl35TIbJC1cSKb3ZoqFkZdO7RKt6OOum+pGe5EaAIjNa8/d1
1hDvI0eZi5NYBgpqhEmAarsshOl2OLCv5DTAk2ftpLYJg8VwuQO6SDUIg82LPAjf
R2dflo5vHamiFRfhY4QEFr6LJ8DJoa0yQE88lIEyeIEf6I/jFKfbjrdfcAODUiJg
R2PVsV4QCPmVkNzhLWmAYf/EnsKs0rw6P2ox2uCh2Yyc1MAyD7PUJOsUJ4bNmEe8
W8VNOIQoQ9JIvEyNJDuXM1wPl2CSelMU22g80bDivdbQHoSvey/a/gwnQq/X/9PN
E6Sfz0a8Mx89t52lArogusEdtNf5zNpa+vArprYmYzhXrufEygGChV0TBoJPYIfu
y6y8+OJrx/4IhyS2eGC/eNGdiHBew5X4TIHI20n1c5aZRuNMltfn0ydEOzklKP5W
/CKwOQ/nDG2RdBN1WTK46PU0/QnWTJB0S4twULCf2oK0fEt7RWAD+CrvDQ7wwuTc
zPMbrZaW3+hoRobGCvKxPn4sUXytoH4F1K9H9urAA2hacY8YW+SweoDY2jNscrOw
Ln+AHHLCRrZmNUpKxMOjansyHXkZRWNI3wsOsmWbqHOQsSNIyAtXzT2zgjN/68VY
db/bKC8je3y9ZdsCC3aKBR3W2WJ5Z7xJ/SDbQl6RBmzmzn/a6fZxY5Qz+yQWUq25
WZlAug+F2IqWZRCNAY2claxozSVH/RZKzAIDekRJhEcMpp7TyG1jLdkHP2fuQnSW
PUD2qnMZHtKVseh9ItRM5j81TOyfVmYy4+tMy82Jhg8cd8NHeCv86DqpuJDoZXB5
UIydhlfJJ+qRACAMMr/k9mpnyvqxqmRPNsx3WCSlhZZo6JjudhSp42ySFa4HGRuh
WZoCHx76UtHHZMk7NYCzuP67KyBcujIHmcXR4eSPU4ELRDWHNBKkao+F/rw6L80Z
44bfzR6mN5BeYuUmTTPN4cFuNuyRWdcrttCdUTMoiCN6gtDnPMIBHRsA8lmlOZPd
MpCIKKsTBH+6EAuIc85xTQ4lUeJl+bfTu0MURy+GwOXIQcPbSUCoqAeXXqeGHMI6
6Ss3m7cq0sq1Ov5AZ9z37GGtmCq9yPUmjxHrc4C75RkHveGm/t/o42HpTtwXD6Ke
ujOlN8QCX3ooNhG5OGAlV+j+uiSMxzcaH9MWBGzruxfhOBDQcefwWKsWi9HcUSSY
mMa/8At6kEJSe038zqw45O/4XV0rMXiz3Kl3uPbG9eeiWzOlwOSMYZ5nLfralihS
C5AMP64a0kON9y6yoDrKVTFsTDAQQrcjixd6gENP3gzwdlpzHy8OeRFRGfMbNssL
CnKioAI3GIxw4bSSTiN3z55wB94pPwSEW1wHSX8rRcmmOVmnTGxf5w9DYy/XURm7
s2XAiuztEaoTztjmWnPAMKbCbeIEUOnYGnDmMeRlcQuUPO/6sdTcRGG2cTn1P6ee
YCqgCEnbcdLbT0vqhO3kesxDiLtW5IrNP8PIGODZWaT6AkXd9Cc188WNFr3gka2s
qP3LzP4amDUPZ8+5mRjFM/CaCl3jSj5S7zAgUF3qvVJjd1QDrhy8h1bB2z+OQDbV
9qsQPL3eDxmlofkjJtd6/NnViFRnUObsvV/LyKSwCUdt3x6dNPAf0F+oDxdFaqsP
uXMWWQVGXTciqJy55zBFp+as11ppNbX5bXrPjCsBEm5k4K711A41GuF2ARsR416l
PXXYyJzmsnSowySHibeBfSc/Re2sSIaTpXLbo4ZhjujpQF1gk9zUkaXJyqyGcWdw
mstBJ7ylzWUmVjbnABzbfW5tHwtoXGvZkhrh71yfPpsh4wfcP2Lif9vVFlvyZJhf
0mMLrTQd6X6syr3VJJTJ2OMLGtFdhZnbmFaO/14Z9Krqgg87wBTsaCvfz/U8vHbV
F1N1QzyDXMQoreVYQ/pHQvO9eG+VgIQP10Rnp9nIUu865eCA2D6aEIZXPVKuLR/c
kBq21nUGeS0giEqWDDpAh5dn6DUG26jCnsmyzNY0pMeG+JQCL7X7Zm7KAUPeye/y
jMqkUiHnl1sGCT30VWENOavpL5tHxdVl+u+tuPNADINs2bqyUmfQKqwFkjtoT5uh
gsa0iK825b6mMW24YWFqxpalwX96nKCpSRycwalIy+c/xDJfXN08OQ2qS6EfGF4i
42DiNpSUvfNGloM5BXKmA2jSwBRli/4V/C78XpEflNrWUN02OipyOgUk3RvLM2HV
5hGxuTKc+MqwYtqy9B55Svnh5PZS5ax85B+IlPh6r6dzXddJHFVAq6VKVMK+ShkX
pIs8OAmFEVR3smqgnBafBGQkxZQ7MbwSVnKv7uJZg2vFVXHYByik7unFBlbxfUy5
tHBVUpbwKjd7kN2TcMQk/mzK/bDs+DI+s0wtNvyqNPn1qaKpnOSQIbnu+QlRlvW6
X8FMBaoULiVy9ihBa99RwFXorZmepOXVmnO5ZobW9AZICxper5rVB8ra9XIju9AG
iwzeY6uPkuCcjgKHHcIQluXI6IB9NoFk5GlQsXmT7YAXD21F1fmIqiJQQqS3C91i
9IPddaCC3DU1yz4+QKx1Rxym5djgel/hjHKV4E8zH9OsttBLJ1YU7907BM+1QneJ
prPb484LuJD9v35ByFn9NCAN+/6wnwvN8Vh/G/dTpqfDa+KMwYykyAmVBOu7snB5
s/84NJqlMYuElOAPMxlSDPnpK6B52ZpAA+8VqO4M6+Lcd+tnsRRlsUvnMLqtg3BP
x2k5+lIn/SY7qoFkgpcizsA7YayKPE9lqqoMcrem7Qe/ESEn4FMjAKDZsj/iE5qT
FYTJlda7r0Yjt0uIt+/TQSxb552+2wI1wf9MLapfRR8v13izOi9m4YWb8m8lzqF1
+QNExIo47V3nNG0yaUHQ9v9qz+EjVnGT3lAq5/Nws0w9Y1o0bFbsFZBU00Yx4t3k
rWl+FDWugEXVPWh4r78PADmolzspFrQcAujqLMYazJr9d4TpFimGUcCyjW9ss7TV
n1od4uC1tonV6QEE5DSFECeW9+K088gyd22i/1g2ngpbWMCUq/Hwbc7PFtAs4SSK
AbH/2npkX/wpBmrHJoJjvYQ3y4H+Y5QGaHivBQfk+jTlzzRWjdWEQK822t9iBlls
JXQzdi5mSPeK9hOFzSHvgACTsD4N8oHx9E965h0Hms2515SRAhHpd3ULM4vy/BHk
KVyRe1/+5ExKJyZ+h1y9KuCrGiW1BkVGpJqqjlo5zMXhgm0wHBKtI1Wx8TEatfmT
WYn1t5P/Qd+yBnBdPrUVPJdbwLs1g5EEINdanjCxPYUaslJoncy5BfhVWCCPqstj
e3GOTYXicCRGPgFcgiwOTkHOE8/xxeXzpWOvIZGQNtrzWGKFz6E7Rw+OsoW9C9mn
ueWl+EMpLgCKcrs5axoqIavNu5e62BRyJ0tKrSL2tjq/T2gloGhcE61e0PJDsIOr
7wuIBDFVLTjzwO19YrCWGwk8u0zUueIDQr+p4zATQ+xPr/OKge0PVzPqCPiw4bo2
KHr8GMVvxbIBWRslLMJ/BZUMs4evcfhnOUosKWSNl+y95q8Z/D2lsH7m7u6Dra6/
Uti76xFby83E8cbSOQ3dO1xQCWR1isO+vlfMXkP6dWDUOyiM3+UU5btjymNP+0bR
kGvmai/pgtfzMlRDl503zBzcJ+DEsrM7p4I5RMne8aCVKsTzfNOO/JEH4+DoquIZ
riMo+Hom7p61ShdpxR1Bi4U+xoT4tPLHnqHp9XBpI25cdiJwVRLDjW2t3Mcz/8YK
6jsbumiB4tymswJX7+ELnkvLGyOeGPPdfV1uajRLZfPOxT7BRThRuwLowjI8k7LX
mZWNye4vgL9y1p/vQXwjov62jHGG+qbR8Q5/NsW+SdV7bh1EIPMX7OFeyvw0iZqY
JSVwX0wGxYVw5thhyXRbuLsAsDqz/7NTqfX/7u/lbBH8p+28wQMGvlp1w62j7qe/
fHbiMYY/kldPCIsx/v9wrBDHRQMva+IL/EhvSV4hIKcqm01L4UK9NgMz4eWZ/EWP
sAs6FP5WyzOa6aJ3XSdI0FISU4hyrOhfQqIeXfskoDsxsS9lsYng16nstXCIqm27
SCxo+d/uWe4A0gYBrpfMw0wR3zr2bdSjeXeuXUicxPDR/n+eimJOFBmQc4BKyv4s
ielzE6utID1KCe1qI1rxFzFOZGgMj2mekBFxXtMEgva4sXD5cnSXHZeCk8YCgnN6
CHzR5u11YgY0DUVqhxUyE4kQtsFAUapc8IY6MGaoXMIzQvqm/IutUFqCN8f8HHa5
XFhCsakIqP35/ad3sZgjMRYJYBSrGLnGQ/dlfPug+p8NFOjIV3ZJ5349ctPkU5t9
IkdZogTF9MxhmBqgGudPj57aucfHnX0KGZcMkvsAWxynxLrZ08TBViCE94Nx8j6x
DYafg6jWzKNEGrgoNlH8M4gIYbYPni0so8vlqv+KLlcj/iojLU6P5axCjZeptNDo
c4tAlA1M8ZQxyG/SYiEInz3mR5nPTWEO+DRQwKFBkkkbttf9Rvj++foDmuQATgic
LhRin8sDi0KVxMHvl3cFw0atMdrxLeONiP6E5erOCyxWSN5qfis2Xgol16Ba23xU
8uagxRAcUyzC8fM+Nn2ZoadAyJ16BjBYaWkeiSGbtSweH+bmwnezTbLc61GEe69Y
ki+XzczsRzquQjfbhdiXSmq4h56I5N0//giyTaM+Mg+CwJEEwRTKP7VOghzx9l+m
KO240I6vdGczHA4qAlAz/klk/1q4meqSSF9kQa44vDy6RaX8jpjXvoHWGlEV7dS6
YSk1LZ3J3xf0PR5xlEHVgFpS76hzCkcoeQ2hOv4Fp1qUtoYOuLFmDeGKmoepOCNz
c6y+SQJ/Wivnc9cxlrIEKumrn5i3nnVbioOe4AMd7ZAUZb0PBnxNjX+RC74ONtph
7N7xFsSNAxxO9PJMpiOXFkF2f1QYA3oqra4P9II+TCAAzNAhM9KYyAax6AiSWVbb
xzL5uhOGk0GGu/B4kXwn9Xxjl+2slRfM0zBfqmbI9QrYVOVtQV2zH1N95SWd8QmV
pkR+Rj2cvKoeRGXpXCb2RPiX9i/t4ea1gTKj5fI1S0+T6skOC4dQdVf2B7hEPTfh
yQCh5bI2vx0UWQPf1cysh3bHmTS0HeO21QrwhOnin57a327rhkj8UNYuwx2Isxlx
7ep7+S3SXKZVeYjpzsKHrI2N8R9pqkjxMKvRoyQo0HlB482MgVRdQkyJSg0OEBBr
7buLOIYHuA07nYtFNh+JsHaGgrd0YSjyRWzjH7DFO59LMebyf/sxHXXQv2i14cgu
P2/WenKy8o3QZOXIKZLP2v3Y1uP0UYfx66XtTMiVbHiZKK85vIlrDMQG8qU1r92N
W74XjYQKgKLH/+f5/OVeoVUUgLXz/tDIA5ofQxGOAYvnvFKjblaKeDCpQ8Kq6Lls
5LO8ShomWp2vZMM8vh4ahTy/iK0pRAW6VT8PMcvUocamaE7wle7cmvQLLJg8qNGs
UMwF8Yg2bEpxl470qZyfVru9q97KWr7eY3LG76Kh4zvfYXjJKG1gIXYp6YDTDEu1
pqT4LUzQ+bAEWz4+vB0oKmKShRyi4svJHQTg9hlprttiDxq3iTLXxOuYx8/tu39Y
WjzQyhmbxjSZ8SNEDBEECSuUQrAz0Dim3oKHSfXfM0EWtxMZMsBZUn3numGP1K5z
/uLW4VnNenudMn97Zff//mtl2cWhAkEYZ9WeHsEEEVHrAGJPDOclGV4HKSXj/aAC
JMHR8qqFAnYjGI03VaEMgEPQvuLzDHL0Q6grcKSXdFTRTjTDE2lOokUNVCflMb1l
c/OhrClHtW18ToRUf9VtVwG8fLKcM54D1QsyKX1fyuPSP3wQFfJLB4oiZgQmLt7Z
cDA7bRgVCQb4QPHcZ//L6g12UQkKGe5VuxzI8Gg8J9qUXPAqv6zHRXwIVy2jF5+f
2Cekqcdp7SOWik4NSULQ2TfRt1f5/NRf+sVZxoT/hz/JLk19ODfcFXKVCRoFW/zt
GT2DIgiHP/RaIKEOVq1HN/UNHeO0KKYUCnAwoNwbJNu0eUDS/6kI3USbjJbQ988P
GSp0yKgvm+g4t5tuIckWOqqZx/leAo2GFpTFkAviPATzv7IbJt8o75patxWe2OA+
cTNhZQCRwXyS0cCrV3e1ScrIGkqtnFZUg67u8Jfebc8yyCnpBH2Zas+BBYierdff
Ogo9alI/2sIe7Z+7UqXkgVwG29Yftzeu2xtibloerM8PZW89sr/oAwhp4G6Ux4nG
PznA5YGr9fi1pWHIFSzY30YVDYY69YpaWbowXWIJ1q7GWUai57cawDFlJOmJYLXi
7hMzOqv5Su/m5446A2C02ibBllmWIgyayS29OAN5puxayXsodPyQHWu8VWw2ygxd
ncY1veBY1Gv8aHHzBH4KlCWh5qOA6dfiQ8zBc9zFu4/4fo0eA69BpRRGlJgAeVJv
Gjjuy3gVFsxHGuKkOPzASUfBke1zNuJFRfQH+Ja2uRNWsF0a5Q297eOtcqe5Zpd+
DKCCNVEMvxQJHyhyGOmZ4HimNPOJG97jAJXDtqxklc9NwStVEquYJ354EBucIFyP
U9bnd3/Gm6k9POeoIA8e9TlpV/Agbrb4pDP3eDwtJJ2Pz7696eKKTz6BIx1xOP9p
Z3ytJtjBTZfdnyJZAKd9hSbDprrRS98OXWsdK4608mlKAthUgwxnfN5kDX5xSOOQ
sVbg2sjiX9CcyENXIIG/UYoXZppBvj8tusg0+x5/qTNaFC82Yf1ENq0sY+FKWbg9
FOLzpbr+O2D9/6yUYnKOKoC5F9seBjuw2fT6csqrrWWH7o1o89yj3gDiml2aMlBG
HpdhfhUak0XMfy0O6GEYAYugic6nZVw7ayziaUO3BOzQZl00OplJPeu66GOAvEqn
skYtx1sFaNKwHGfue41+BUpG4d23rsuCvdYl3cY6WklLeLT6tLi2eI037AXWlyt9
UZ+AlS+jKU1qGCCEKyEpshk84+CUFA0CgmdZOxZVQOcINPt4hVXi4FJ//7xXOsgS
lVk/5ID7QAkepdeCMQmuTF1mMbU6jHvqMFE8yP/qZ9uFyTPJ0NHfTVOaZA/eCk4+
L/KjQyZRkonmB66CDoHTt1RbIjnO8QoOLxo1lDja93RMwZLj4ySbPGmoNiH4eJEK
cHNGF8VyCeXNFBTxff4//TznxbSFhpd3o6fCLFG+FSFwQTlMbVsfUNMMo+1J6LLf
VAwHtFhJox5Q17aO3y5gd7h9H/5K9/ghZRkZZ7OLgnKfwa9q+Oeg2iRFqSHkxDae
aA5PEoiFrkbwA6aPHceX5+wtn45zb89ShFAw+DN7BoIWaQPQ1+Vbh398ezdhnpRZ
kmmKOZCbro9DdSaxzHBJYGvYi3uGl7fDm9jmtj6Ev1t7t0uWrvEUYCk981bKdY2W
E4Ci9qicTRM0tSj02VwI30RzGPs4b7l8ESrGwEC556b8JN8AuawBcnslbQpDlYXq
TH6YxCKSCRegli0YoJ4bxgDjFf5RWtgl2jM3DdKrksiGiZqXTvd8Old8fqSw4Qiu
Igio+mZLp+JYmZal6J0BNxyKNau+qrbdrFd3q1imDULyWTpzwOjyvKPrne+rptx9
Yis0qaNoiX7ubR2z9n4WC4DAb6LVSJ4tvFM8/2b3fqwenRdaAaMYeO+18FEPWsRE
m3SGlG/DAyAIjVxitCn17BzZMqJkJbHV2e/y+r+X5iPdUBt1UJQH32vAJuPug591
s+WJzAxpi79yFI2F4c3VyCA8YOTOowYy2PxXexvyRtci/Od+Tn5eyHiAh0rP41EY
pIrC+0oAkk/3ouIWmQrk3nHFzKUem1fmOEOPEAMDd7lIhaquCoo4K3Uuv+l9G9eG
XP6PofHvWkiDlKQ+xhlgcJCoyyRepULqpSsrZ3GQ2BJY8Lv6IGC6/4tcGA2hQxZW
ZBLiPeAcIHQU2p8dXlWCphClF41R/woJzU7kA+GZDZL8DYpruZ+ydAdrKCV3sARw
Lk58s4JL4ugwJS0aVVxkmlsza0KbvzVveh0haE6Trb6VkBmjvDWkMdgxhnrJ0rCb
2OMT3CSCZFyTZ/wkDQurPhnJEiHRygWnbAqyBYYtkaBgXMPHoac+xNlhPKduJhc0
XsB/NKnIupOogT0hwSZsXbzGyws6Lbdb1OsiEoxNVVNuaoBQoJ2l/+uNFJgHK5L4
Xa2P6Oc7/i3Fi6Ey96m4FDauXvy6n6rbvvsLCQE6WfCOJ4nmOj5p+2lW6aOYak8t
SkYDJGcb0iM4UJxZG4MV9V0eeuBcnqlL4I0xgztRx/3eQApazVDvn3r8pyJdUZb2
o2W8U3YS4cAbu5TmbYbzy+VKroaOm0DwycXJ8pJfCwElJVPKBQaAmAnWJOCc6DJK
qp8waIadJG+ub6oB/y/kTBiSP3qkphEc2jPUK0tDYIEm8Cjs+/91MHQuxTdOWhpT
ySfm5gjtZjtH4kGUvuBC48GxQMx/EW8TqqxVKfKKbQAo972CDTVl+1LSId/GdWwx
tyVaEhzNKtLatNsZUy3T4RQSDzOQ/ERKO3wIrgixx4hMnGDfqO2kJCX6iWw8el3D
Rc9yTl2f/Vy3An7H6hyKN0lVUrv+zaQbKyab0IEvU2dTuWqE/4XaCjXVk4NWW6zC
pNY+Xg3fydwel0H4q97EFM8DQIcUk/HoEZSjtmmj5eNG6bg7sAIYd9SPggR4M/ae
Don02wG1j9U5lzf5q9V2oVrrOENRY5EKoHKp/E507iUu7335yewoPp7zkyvsHoKV
gXltBZuGnRwN73eCVHFFnsnHUTRcdlVIOmd9IkZYxDmQEzcZL74UCRvpV0v+TcJz
6QwjTSRJaThP3UL6MAxXF+go2dpr4DPZHNzODevWf/GcCA7MwC9ktl+Dg7X7awby
0WrTepSEd7L3SRyHbvc8Fufwsh9Jfn0YCH0sWhAQj32893XrXoxyQKd8ZTf//PNn
lAsfBN5Pfov0XBFhc28WMWD5nQBmoO4u55KYiTTdduAtsVuyfnUCE6x3N421RD28
YBrfGFWkE49R1iLyhydFUEbA8Q68gLhawd48zrB/jPl3BN7GMN+gOfdCxX6kUx+j
7bvgxod2xiN4xgQbVsCeDB9QYOlAHp+GT2hkzDeJ3ERFr5brEf1ykUOMirgT6VSd
NTFaPaUYXFmSezkYedr7G+Od9BBaIaPW50jntdycT6bCvyDY9/Hae6VpaAyUceJe
mHuEZggxbNWwjA0ALzh/skiV49igJfbxkOnekmEThlIdVfUXeuWp0YGoYyzhQPIY
bhGurmEmRqvDpYMwSTQTiUFclpDEEedDbHteWivroOIWswbjBVzHPbGpuIxcAJdZ
sgpiVp3Q/Np5DV2OT9OuPagjUsu53bS2TNIFVcmy5SzhPWCiuTbqOf3LFGojpoLF
zeMNrFSGYLxiNiPSF9F3O/hTAeJSuFCBNIldFHQ5jvaf/VmKHlDit1E3hf0oio9B
Qzkeq3fOnXby2vymfRvgFVi+a3J6L0rMzAdLShO0lC1QgkhIIlQfLkCqmnuaf3tF
O3zyfmeOnmbPnVd65y9JwlnKRCHTRHmivMrfw+ADCfr3wY2+34YvN2CJnTalzhF+
YU++iuuFASS30D138NYS2qXJO0MbcghXZfzc9TDCn0PdSeFZlLcZYt1n2IuYGVyw
fXiOUkRLdBXhqQ3BuAyVe9GiikQtW3ZD2mMm7mEiMZFnY+5Nb6Y38KGDh1dxHQbQ
kpz1CM2MkFjGxBYyzlt6WlGJWC9nmCquc/GKONOc2dB2gm55ZlQHEGz1taKP/e7S
82y3Wjclg4bECwFo54pEol+5DVvO+dpj7MXptvb9uKeyQUhFtOZd/d7CNxDcTRlJ
tbu7/EsUC6zzcnl7+i4Jy84keR/J3IB5/FWRtU/vkuNmYaYc4j+sRByuOmkWp/Uf
zzRWdD/xd07XoRcZA4WmMTTV+J7WEXkj6SdF0F2PDaWQlwx3LaAxw+F9mj18S0jv
jcNXIdq0X9Xs+7IpC+qzELB74mOHo6gULzXROn1/Z+MHe5wr0n6ukG/Sbv75GEu2
p/uhgAhgp++HxBzVp82/UB9UJK+HozqC0WiCsuY8XJ+BwUd3F5LYYjPu82SQb11z
OaBbjNQn9tsBQiktLr2/0Lty+T/TBt77T7+zHH+Z0mODgOPeD3lOsYqSPqKwkIiS
srKJ/TOfruckLdsY86HG9HyQNZ0PkYaQDr9ZtPB53h9cd67zlBBMnDxTtk4jkR0I
tBPVMANU4NFjH/lTySAOdONNWfsPpZyHpPSB5TSh6G7nYNrdnxaady8QvS1f4QoH
UY1KkblzKqsOnItMOX4Uz22rIsV4ocOYJPYvZYFl0PyAJFp819OryOx6MGy4yps3
gbTF0JWScbgP2PjouGLouF204MU5HzAd/PyU37ek2uUTdQJiqGhK8CggcDz0rlPV
0M2m4hNGjRvZq3FJVb5jsl2YDg87DH1j4mCt6QqDwk9SQoYsz3V3YcMo83rLzWll
wkiU6RjkPVEAH5UltUTqOwlNCCP5S61AwrnMMuA/zQOqG8eLuAUPhcMCH5Ahneh9
slIzt7hnM4ap10lr6avjxuJIR9/cWNZ5KfRSgyV0Eek2HCRo1gs8mCv/FPPlOOwJ
QkY9SGxVfPyRXEOPWYIShE3E7VQJ3cQBPzeb3dtJY9Yolll0efkhgYffBnWeFSNF
k1KLciQj4GyniRK9WSpLA+MehB8BFB2NaRLiZ4JFemkEn58fJ1Mgi2uTeIBXDdon
bO0E7mz1gwuL7bH8hytasaTv5PvD5mIWC+2YmX3gAamDIj7XnK67sDBpX/OII185
kAEbXSJTuqtxF7Km09wHjqajif8QFtP/qDTiNFO+VBIZreLHdtDlIk1aBXLyZBQb
t115nRTGw5EuEV6IWAZGU+wdbkFIqtCb9E1GSRMT5pG4InGqy9yGbWqvknKtaZkG
QHj3t+1WY+WbArziU41LOlfBVjdw+IeLPdn1YvfbNcu3td0wKddq2UvPYJ5Kj8W4
a0HvNkaL1wsBJTNUKwCVHlhJfIlIEEA3ZC7jlqk7JXpjvbbSI3Vh1bfGSh0mpiBt
Js67AZ8RgYoVMiTkxjOuvNrsgeZdIV86oKEBKhOfKpDKRHT4C31WKLQwIm9tLEWP
q7E3j2iTtkx6DrmK5GFV9hY35aX6wRha6KEGhYH0OsYHQ+rq1Ho7CcZhOxLoW2Bg
6GYuqYtAwDMtDZILm6qQsnuLE6fcJQjKqvNdrCVuLsSbgCrIC5h2eIYkDPHoPbGI
E9XhM5+W+acBael16IkMAVayLY+TLeVJuJ92JehiolSstnKM7hNEBxkuNF8xeeCk
afAKX9jN7Mb+4Lt1ocjrU3v64axJv4c/7NtcLqwysKal85wgqGlKc3nvBAmQLqex
RL3HrxQbRjhzYwqWtloEXawJ/MexkP3dF1GcwsJHThsC8prBlwmlJOxD2qG8gD8q
Ih3yaJKLp+aF5gV277z0lyPUI149IqHYHimemcQUI8TnuiLArTLv1g+ENplY7FxQ
GIBWsW5eo40oOLxSZfRGlU3x7DNivRpmoPS5XskWj/T0S9SEQbojIrH/hTaWXREV
AwgE+E/9RRZVHQRY1H2uc55Dco6ACyj7XGjMjh5bJAPoghpcTRy0fkjR4Xr+qm6D
rHW2xAwepavYHZq9ZaPm936XQMne/9JA75ALT7pm9ZrZP5GxR619H8d1tz5gRT/a
mQ+hRo4TKRiQHpETA+oZmTFfMqOKd9tg6Um0MZikRaOM8UnswZwTtBahZy0ZFjIm
LHd+81jkNt5yonuQTIXxgX92Gr5M7BIhDImGQgzJuFhcpaze2cAxwwqXuvT++NeS
v66t07cKyYqIrPsFCf07M7JEmkHCtSTsKKrkrG1cmbdKFMeZnXz1BlHI4NiQwAKf
kMJlwB4D6mtwmymDk711mGsDqEBkBy8fNL6I2bk4qgv0ev83H19wGfB+ADcG5X8o
0WrdqRtu/DSaKJeav/4XGO93y4upL0FTifnPifmz9Ac/luoLT+Tk8/5B6fPa1OnH
vZdq8VDVPwI1r/YiT3HQqomXwlS32C9YdmnF+LBqjtMhBiEoHqLvqDhox9npTB6O
XjE4iDIRf+NCsY8r/oTz4hSlkytkL8QKjXvCkh5DHPHsLq4+MXycpVNDX/xpauxO
+BYQBjkAjvPDFStWorV12o/H8/PplGFoUqAqVByTIk8vGNNEQuEQHRYw3+rIrL//
WCePcptajaofEeHChrLNkkl5JeBpF5b+C906JfdB52SjyywZ4mLNgogazaEftxqn
Jd37F75VfQIOm7fQlT27y3MirnxLNHXlqrdDHOHNY68pXd/mH53LbhP1zcdvjh4v
gBGFcimNrSFTfaf/zMji4jEcxH5JEQTJOTYyZh1PPWU+fToX2RGshH+Kca04Ja+c
gK8bfPXcfhXqWjocIU8w5LrLOeeBEg9AhoGoJAs9978fCSXaehxK5fut9GnXZM2K
yLyIyV7VF97stU6Jt1HHBEsnOeF6JTxveSKyp3GMeAEmDvWpzLx6H4H8JXFjFZgY
C1fj8J9XcScVjZSVnqHkt8frv1tm2Iw7O/mveznjQA8unwGNb1TroiR8AQAW4DIm
BNGwjfizdeYDTUD65Lc0OkGNkUuOvqMUrcDO5FC7P7/HBmPemTs6kOQaNrymKX9B
7px+WmkIqBn4g1GC/sz4UUpI6KDvext7E20XtcLdL483srdT5rdcAZcJnikXKpAn
1+Y4yGKbBGF8KeR0J2W2pUkDlszkqHTjdGITukYuz9frdnj/Tq+yL+rlnXXh0l6S
2n/ch9Y1WezLyb2vD9iri/ABv1+CLTpz2J5SZgJ444MYlP3a+oNjp95IKw64m/5e
veYYUnXTBS5Wya9hwKurwxU6ekUOLy7OVkiqkpnXbxiIkTGjUJW6si+NYKbl31CW
nAXmv44xW1e+biaZgLL8R9XS49IwtU3cCHOx5Ymyfi8Z5e7KFFQLdKGNc0BKB2we
UpGiF6m210borgjDXruJIEEFqCuLPdbwdUqeIWcvvGCTOWAmnwg2vjUpXfiP2S/4
fTFDEdsMuG3WZP8JTyVROOIEXPLxiOjQkKTBbvQnnebY0jWRwg1gCoQNAUb58ueE
UC/tlzlIQrpMll0Jh+gUSpyTcuUM9sS2ea5S1IrTIUcCHj13wRtRudaJ2MLfVeMU
8UM0OcgcIjjvJG3qDXHHaaOLQj3zAthMoVjmmA5aUdXapvijmbbBHOjrT+/nx2FR
/CL/77lmonyBVHmDGrRqB1nf5gR68fTI+eu1XeHMBSbRp4CGmctKCna+7j4MZ0cc
dlJMJ8zRzkjICPsCyFhU12wDnqX307I30cxj9w88BEC4/3zx/Zvf6UkhJhxPpG40
RuIJioXfjy8z8sCc4fTcQSVPx7yDXg9w5rgqn+jKlYdMrrOq4u5KrP17eyZcgfio
GJT8R+R/+fzqoRMauPhUjJR4TkRp+5+pHx1Y3UIoOPWEiegR4+8CMXyxB5BqD69Y
Uc/r8A7X9y8JiUkqCmw9bXkw0qPbism+/yfhLmqFRPrBPEAA5NKkCriA/XCjqqxw
GvKMsyK+I6ZHDYMjmHInw4cgI6VRjZjUu2AnZ4nkNyA5c9k80lP7hyku8IAapE2m
6MBmRXDHBVrP1KkojjNhEdtIjJw8ZxoggNLWWs1Hn3wAYzktq5SdRd1DbZSppwhI
BZoEaYc1uR8goR2lEuHtvAMaWlA2StXy7pUlCJ6FvwEaRk07PZJvvS3+Nr+LQXfC
VRTnkh+gtLSpQT7AOnyQgoYl1ZCHNysrRy2xXCl3Adu+CM/saFXv8BncXyDb1yS2
ijj1pzK/bmwSBxahabDDBPxJtXhvzz9zNEc0RyDJIOZy37jW/8JHx1Wcn68+Or4h
HWkW82qdgC7El80W2niXHpreqYk9VKI4u0Z4Q0gH7NSTEBBLaie+vwsS2PhHuU3R
EPFPgiYsrDCAS/Nf7LjhsJf5dYNb/Jaq3VNNbahIKNGYgFiktV29b8qMkLX7lSBa
VC6YuUGkinXALyXzZyu+KLninzMJCqbsWs/LvtA14G2w6A55sakMjgGgNLsXi9Hs
VeLPXAVGDeFQPOh414Mbakbtx6yMfnPUTlxVzTwXpJSNBOXGzc1D30R4+n0VNZq9
ZyIpicFkz0xfZOSxZvgN54zANuM8N1L+gGzW+P+EH/2G4+qc7JH9D1bMRHlZ82+D
6CMDqF2c61y+CIDLm6JqfmA2CIPAgUekS2CHe5D3gqiX8V1WUXFyw4bb9udnYez7
diRB+cBffMYmiIEpP0BixIF5Sr4xcT3nKERRDBStZi5YeO8V+vTrXOzG6rE/ru0T
itblTgzARsgACAM/SddqhiM+usmRuRWGpItb1GW43kIvS8p1Say1aoZ7eJ9iSs8a
N7/9oxU/RHpaQvMFLZWLlOd+cJrklYiVHqmr/A94KcZuBvh644K6BcDznjHF51ou
qFvcEvPXRPYYhAITE+scJbdAfJGoAU4ixQBBsXW7CiWOrpTfHUKyr5Docdq/koXY
lgQmIKeRFsoyLZBIDM41VIOp6B+OMmfyL/DlijisNzNa5wci89nI+oBUjUI8IsVp
NkpVcLNpqTDwBp+vui8/GyyllRiPynapyQVyTasQPFFzCC9EDE0I8zkrZYtWSGMD
2lqnLZJEDNOdh/ZrC4jn2HF/bXISV+4bI5UD2QRyDRM+OUm9H4i0LMK6/A7xmp8S
yZwxf9D4OsqZqe3Uf1O0FgVXz0EFUFnOTvsu/cFuyMIjVK9Iqo2Vu5jTjDK2uEKj
YW9XqcpE38hGQ3+pU8DJGwI/qP1fWWiInGTnk57P3uhEd77WCif8Ls2xFRAA4rpa
4sAIhcoR/Iao0nEiNTEtrt5F9jI1SIyrART14lc+OZXlPAKUqTDtnnv63IoefmDQ
KZ9iddZyyRomln/QGxcyaojGx5Fk2r5AKatBlITIjKXYiN7xMBeb311vyIG1JzZF
GDxajZbL6nG/Zb+4XOKxLXvrTCQFM+C2IUOs6nnxHUHQrUf5wvM8C8AVSYneCg32
s3dNc79RzDNQXIKgGqw8ICYfmph2KJFR7EwB3HVOCG0sgwgNFCEWKUwNE3VdFOIu
OOzwZvJlhK+cY2GpXePUeg5nLLBt0JVO9rwqQfhv70BAu2MD6e8zGnnnVTMhpCPg
DjXk7+AQQwAzsTC04lUfyCVWDWRDOeOHVaf53FGIbOUngbw79kZ/6EBAvJHxb9wK
ZUHOk3YRKqxZHGu50iXmIT0G/zxZmE5Qu1jhQfxte/FFQ1B7WCNnUtFAUHDQKZmk
Tb6nN4WRMPuEBO1x5ZUwCL3jqeDfZ9rWJ7dP6VOBPOkth+93xaoPfF602dqbu5cQ
r+JruJHFZjPENwhi2en0Xycd0Crb3fqdd/Q73+Mz63INTc1ykgUBOOO572TJxsC8
0lh4FY5NIwfmTQWLiyQIt8bm4TLzdGW5hY5u567h+2OxiPLhpSJrXCZiixD1inS9
C6ZCm8yYtm0eD6TbFCf/omg/ONg171/CkOu55VE7cXSx3Abwe8OctJQnj7v7pL66
MZlPfJcpt6qv5x2Gc1Mieg+DNUps5ye9voGHjXrUAs0TzjoGuQo0H4Gr4PN7XB/h
sG7hpeTTwjpHfQp8Fh7AX/IKvfGw1r0K5+YBMkToO8rS8e3FmL4rpGSK8rzPg6Lj
GKcvmURXQ8G6pKD723sfF0qZpb4rE6KuX0LJWS326qZp8tLQ/CUoOfsG2XxfRRx9
73KpMLU4xBCgU9gVtBmK6j2sAl6C+k4WKsVMrEKCxCA9MQvCTR96NI+uqCJnUz6H
XVm7FFb1MQcexECNSl7hwc4P6HpdlOXCr4AA4fKRbV/wSjkLSw+J/XO+pO3BfJKe
/BeuTeqKDQb3bzw+rSYc0YPtd3YKtTBAtwe74m4eQaanrbD3z3qCNa3YDZZN4Ztr
WYYQoLjWjqSnVtQXsRPRspcm92Rp1lTN7/Dx6TaZVd+TaQHF3BgVaGy7aF17oMvn
bcmo4U7gUa+n3jwlEhCiAgMR7p3AoVAGJbjR8PzOuDpklY7Ilw1gSlv1Mi+sDJr0
CrfOsaEkfa4G+26zVnBYe+6o/yI+YVuy2TgCfkkcqMDT8iQGGBJJ3nGjFH7XIXXK
XzMbXXBazuXJR/RcZeX8oLHx3IYvYapdLQbBCj4beO8Tel1Q0L3TMy2qQ6WkYbnx
Vcg375qfWPCcKIGt+Icvdeshs04hSkLeyeUWt955vYBQ3H9ILTr7OvHrdaX1kHy9
OagfJb8iOicE6wfHmwwmmtFnJ2o1t6dVwqrkJLA0HoaVzutnGcJOVKNiFCq1M2PU
kUkPmXRAbYppIxzpB0Av73om3VCxvKjgbbSlOzJFo1NhUPF7DBpIRu3wjmQwb55A
leoSoKKNPP7xbf8mn1H4g8zrVQBUhq9dZDuHrXyo/Q3XqZUfHi44I3pD7arzZkvO
EPB4uXGJLYqvLgUiWwPhLpZbm785e9F/a1RHjEYVLwll43hv5oBLWYD2F7T6T/PM
eXoxYcTbt663k9PYFNu5cMo9MTvpSAk+GxBfpDffCPS78PPP2qunhumD3dFy6jr0
4zgHJGFIy2heJwhk1T7FadVI0F0ghn4iQNJcu8z8BgMJI90iozwqx66zzkXjhgH0
lLzT5WcZwbFYKxKAt8bSRt68V4tsSNTWB8bdsCIBjFNXXZcJcdx7HTtMcbsT+8yH
dCe2iEtfjkSj/WagvnZoL+TpiTvJANqc9h5CfYsZ149fRIBqNUbHT+Z1aQwFg0o/
+Hl9Tr+AWK4xQGC8eDHWcbEfSp7NZcYg6JwloQN9zItTusCzYupslQxyeqiC8FMb
cC2y05wEZGOl/ta1+YPLT0cJisK87x2vvCq5rXEuXP0ntaklGIZ5K3lHvvxdgg+3
DHsQQu/j8+SKtnnwSIGb+8TEizq0vq3T3kHn9vQovqlz6rJE7Oi2qodancer4ofg
OQgpqCDdD7Q0zq+8dF77bCn5WZoflQ1yB33DtiZkDy4EDDO8LwIuxzXhWY1ZwADU
rBWp362ruvJKmslB/ajF6S2LSPBHTMk9SySjoK8QXa5s05++E2qse6+d3zkmnsz7
UxO3CYFvbhVaVEQcL3gOupCbB1/j7goTl7oNEzv9o8B0b+LCEXYT1DUtoEg7Tjzi
wK23d0ZJhVqKGSHKmHpPIOop2eSu4b+uL29cfyhFOkD4xXh5L73Q4fUdTkf7KthJ
Hh/ZZ1Dlx0jK7iSkcjJV+GvPwT7FhOSpPmI0oO5gXEoDVUrZ5nhlWCAkJ7zSfTzN
EbVNXi1uubBFnhSfiTbMXYOt31BRk/7zap/C3JxQObZ7iqL3NEkXAtIcuud53/+d
E0dbbazUf4L94mf1sUD9WGImpf1dN12B/9aNsUAoSxl1VTUHs9fUeCn6awd1rTEQ
BJmETVbDtscSDgyHRzSMt/WDYaTF5xwRkt5D4kdJzjOWNFH1/4FNCQ+dzk0Dz//r
MRsNTFcGzugpAl7lExBrUeeslV5Z8fKqu/A3evrzwnH1IQ/ePsqb+ZFWZjNFxnlq
RiSNJqw8OIzBqzd1/Du/zXCuHZgUUqqsuP46Nc++o2bIiHkEKbwAIVzM/s4UtxFG
bCp302l6DSsJw6uo3Iu6oPeOUl8DiQq58wstoMwilOgg4G5mVMgZw9yoPZOzPk9U
74Uf750OaaDxAK4bz9fB5O4ZuSWEZeUrzS0xh0QSGSW9hyt6UHTuRsu5LWnyIXjn
vOETmuej5XuqScXe7Fpw0e/KP+yrV3NdXtaFuzoyp9nZGFkQXGJJY0mq/e8LMnT3
9/G4TWTYqDSMlNS9y3jvZnc4faWRpbp6YCMk9czJIBUipMX43gP7cdXK1b87u42b
QE8eSh1AGtyv8AGg+Ui4hP099xXcjM/oZ2/IoFTrpawzDsSmt683ZQTGDDsKPhja
ly4lbSCrhgODpVgZTXy25kfajDs44e0BW2k8lu/49kSRppsMrPMmetW3pqOnhguN
DT6u/sDTqDtZP/G7DEuGmtz/ZaqkFhqkBpPOVrwhbg63dJmbnNIfyBzuWDSPvW8t
HpW7AxOWCj/5KGO/HNmPPw0GvoDw1mq3FDEaHCb1l7Yrh4J23+rcqqNt9hdwJni3
/PqIijdckNctrJ1QMdlUKRZqVzCRgeIDWDsgOHaGFRhNmPTXjAdcaJBweQa98kcc
UdoG1LCsYmedk/Y8yfW1dzhWpzDKu9p4wakVHl/a7pDn6XP+NJYmNWGeu2TWn/pQ
ktY3txDSiIVvdJXfY+DZIx9QbzdoEp9T+4G9czFx0om5tZo9ZF0l9f+YbPeZNVdy
PgOZcx7E2gf/bezfCycCGKz61iFYq2mpPFcvLo0QMvKFXAJW63w4TWZNJiK4Jj2y
4IUj39tLraeQfrZS9lnOC/KLFuVAl5oX8iEB638p6njuHwkczUizAYQGqvNSUFBG
NXI+rbndJiAUW/JwWvbo4wVVDfpMCn+i0nwIZphkewgqQ19Yzm/5O58SyzhIzyVx
IzpGVFA5We9C/Xfcqj+4VNni5wNAyOef1KZrlvi9sEOSPWw77sHlVbJFR9mkLKA2
EGZMhq0EQPN1Y2EwWXAgAJDyP0cimgVYyaSoutNQCu/fY5y/VorhuqHLJeU3M4V9
4u+RG21llWKpLvxvkQThbA8IEMczHJfg6BynDH54YjeT2Jc83ElhVXe4Il6puDPD
1MViNJhyoHWaOxCoV8/VclxrvoPZS8Y/5xEi6OU1mers0Mv2DqVJmpHegBrJwylm
+aB33/oPc3u4WTTGHsSHjSiUYQGYYJkO/lZuj7AX66F6ViAekxb+IR6kapSXqEtk
WiJvGGpUAkALNnoqfFCu0pM9piCM2fAjqa0X2gnPleqzOFQ7W1kPSyjSlkFbXAxH
cKLwH0+OwtDVMONv8Ij3Uvb4+ACNIyFYfd9C9zie/jyVfNELTu1bK0q5FD+AbFUu
ra2FvW12YBVVboSxwDzzpl/vOXelK0Ou7zJT4uvPGM/+uVdX9aavyX0qCkE0KyOb
Prvf6eJJ8mpKtBPGBvEN+h7WF8cwnPpphrfR8HFInsEgAmCKGF3lCRj+R3VwTiOU
iHXBsIIO/h56kfep7NkJ6B3UGNL2uU1dMP1mJ+mksbD3Nlxe07mKdZVR1npITXQo
/uwF1ll5ZbZvsF8GfnfnNc3DpjuA+O2Xcr7pGbGPDxM1tmicgypsd2n8AT5RAWth
lG9UYjJ29YZFdYT11WEt0IL1wVQI3djsaKbNUHv9lbw7pbOGBL8ziKZHQ+H3sX/i
RGIF/THsIPhePc2XPJw1YhybXVyigRRGHAJz3yeUliBPwGLKQtLNdGJ3L/HCFs+s
JgyAXxIJf7acQAZLr8xjVNFfVBLQ4FyDWh2ssaUVf3UTYrD5q0zBbza0ESDj6SoM
utntQDWyyYBRq+MAPM/vwPTfFnS75u65Km+UpZubZPU3DTbWTJu+KGSSL4hLS1ON
XIxjN4qiFwqAkvagiQEWbV7nAeKlE6vxe9ycXj1yRUcsNrgcJEsdJDGxaYVUjXEN
MiFaC4eJOEI85g/hIlkwOukuLy8KpyDQPyym/yf806gLFZSiSdGQEccUvWjNY+2q
0KnfIGD5UuDebm7Tf+X8h3uMAytA556mCHc7V/KSAiUXiXEI/oQFAYcnPhIALr76
Y+8Viny4CjYqnraRIgL+adc6VAj78Y9DyBMAcs0D+FcXC502HOocKMn5p24Xn66U
7wh3gmhEMEANzF3rI7T/+CmTJHi92EBAqLsQP2piLMRaffxGTsJoAKjDRz75pim/
SoR52npF1iLOgSu46Nrk827ZTTE0xaixS2QLkFEnc1QOGcAk2d+jNWFqWAwLjzEe
uyb0cfSL5EcwEGSdXW51rqxg3+v045pOhEx4LnAJhKtqFWL+Ieh2IfLTinwyBOTg
27CGMxKRaAe064dVD1rEBbLyTyz3w7u9VxYKRs0aH6seZXkVXayLt4DaV+981FFd
nVc22pMlZxIHS4IXQAM4CBGDwseypgTWPBwBg93v8C4R2FnQoi5DALjz+LwDXHdf
VtwswyFa1OQyfbyIrvE8LxmQkzqV035vVLphe0evkK9V39z4Uu6dpEMLrC4tFKeT
OdR+ff35zBtiYWrzqq8sXOjWu0z3Npewe83947P3K/7BYu7D/u2a8qmHszLh/cQF
HzcA4FFl6/NdQjBDrU2ceFDMgR0QOaVPJxVYszWaws76Efl/+sA9/4NulfkZGmCa
zIhvDgockrjtw+aHJ9turqJmX12KueHSfbqY4OVXL+hqflqL2lGq56SmNCwqR1/Q
bcc2gK4MAU1BOkkHiqz8PwTnk7kXtjC8vXB9aJNcubvslDETIFHDT62d3OhThUa7
Pp6DvgW0yB0RbX8zGgUPdqr3LAzAosUVSJAlqEXidMx+Opjzg7AcDA/XR6feeOUr
Zd4bMWtW7lpn1huFiLkyrRFsnSEJ3CX8QFEdDlvHOLkgLc7S8WU7XidDNJOpmxph
v+8IaT28VdWwHHNvCm8AMyF5Owe7kpMXkOvg+fFUTLdr+B/C05UaRdiY1ZPIy5pE
cATdFvHV0mYUT/sTNh36WRZDi5bdiT7B73YfhdSoap3O/gy5yR/FsqccBgsu2AEF
DQj1xYNsvUfcHVzG5gPWPIMN/BQjoMkiPzqVJaqlPqMd+W+pcRFlrpwAn/WVVVCn
d9d0peJRC0wwQKfordCf6ngOyrUlLgvorzF+dnA5EF5D0jz6sTr2KqKUjQuei4kE
chq+ukExCrynZdWLEoPnHchVEQT0+QuhuxJNghd4uof6Rkn0pdR9zN1FvP+FrIbj
E2g4RN7weUov+ExT+U8XIV0GSAymo1hQG74rove+jJR1cI48TnmhT+VTUdJppTPO
eyaqChV88lEGnVpe1fO5ivXk2Mz5V9wWdApZtOLp4pmK4kb3yDPmgc68k4LRXCgj
ymXeTYOp5RTeFuZwaDutqLEWBQzQELTgeUO+u6OxgK8NXyl7PS39jm/XGZmV0455
YWlqhG+sKCutIAF6eHxpXRA4b0QXuYEIInANXp6KcZpx4zqzSbAP6Yr1g0cvl2sp
7tlGcbeMjF9cPLrPfAVAnn4DRWjFQ5wO/oucxOs1E4FyKD/lSU14ToUYWXpf6AXA
7OytAbE+sBRRfeQyxjg9jNLgvsJWaXsTG3v+8UvatGghHG82CLE7TDuQ1tT3dd4q
n3neX2zBfAzLzY2jkKLgdbHofzXbVregGh9KWnlEc98M33uzrfKnN7m5gLkf8BNv
ePqaSVM1UrwxzcHE7kr0poEwwaryouZupitX0Z128oeXCW02BNn5bZp8KumoPREx
gGOBbi5/jkk1INLmWyhYNJgr2UmYGmGr6L4TGBiFLR4hmqoC4QcX+3zcTwnsFI1t
M6aOXGO2aCTgLrEZ9Bkc6bvr/sCUIK36Sfm3fZjyQrdHE/WCHEs8cEQVl1XSy/+g
zDDAR/vGE7ollEeulpC8XkPTfQSMNKcxl63fyJvFUgyMoEHmiILl9gVuX8czf4Zf
ADzKUaqdx38tPMFXC/SBb9ZOwnGeIn3zARb68Lrmb1p6xfgbTroFdKX+mUCkxZKd
yKfo0iDucABb0DuFBVrg/dlJitVLECy5dtpzHOOxtqOXA5sgbbYPqnPEpZuRBmSl
dsTV+ie7UFJTcH9+7qbRPAJC5Cz/2l7nafucQ6xpfI6l0gTaqbS8W3IVqTua5LRW
fwGejo0Bq3GgShndEUS4ZribuuS4jBW33smC+5MYD3CTFwRF9eP8kP1nrnh/BR27
RgrAQEBe8lAuPrAgQyp9Tfz1gWaFpUjQFa6+MzpGeDacOXuFRwnlkzz0V+y9+czi
Q76ATG7jGZVEI4+ilXOkvPLc5CgHSMccj/3AWICBnxCzS40nxniKqFlG9O6bAWD6
ao6nlehp1rUjl8v+bM4rHSE4OUq8Xs3KvUElYwen3gFm1t8YyeV91e+hKWRrB3LT
FcIRMHFel3abGQQFhTKQ2I8S2cuWEdsfVoCI3OdiOL61J1z3i1H9Yvhd62UvDxR2
98bX9qC2ets73cIcdLEKyf8KIui7Z8qCh7kLX+NxUaKVdcAlFtwGWUYZDxxmQzOv
dNWjDo/wwGPBR0SKcbOx/t/cjO+2dBrEhEe/HZuuxNqfW9ZbpoV1TthcLI/za1aU
oaE9gGzLrhzqXB/8X570602iQn5iILCq53jTFJmw8pWwPkOb2xaowwm6wvtXs9oi
gG4A1yzvGEv/EQ5HLgHr1axEzBgtxdkYW1O8lPMYQ40dJI8Tqk+MUOekQAYvn3vr
3/VZHJdOrVIv2vCu04qALm+tgXzSQgYSuGqhS8AX0YDssQllcmspl1IDJoV97YxA
cCCIuQx42CB2zg0BHXKLKDfgw1II89mvyvS9bMSmVQxf1QAZdn4ZGnQgialoF86g
QbTkcqqzx4G4f8WCBD7aPHeFume7XlFh1hQUcLZlA/GeN1fMFjmkD+IhFMYfDWvX
tiJb+kKW4aYws4Tp4Z8Ryr4l4o4olnLfG9pIgTygD4ZSatWwg5rzrFCz2O67qojM
3cTp50xtoNb4DG7OyWJ0UlrhYPcBrUi+rUGJT92H+4pn4Bs5YPIrOHwouphF3qRF
MBh8J1aIvoGcwL1R8ER5Cy4c4fjU30MXZ2Q3Dqxi7vlqhWC1U8GJxwGsbjPJwiqw
FIRYtBJ/DJCyOL4nbYHn43okTRKU7cmXmxaR4aKfFr2aSjHBYgGG4BB7RhaLXSO0
veEkA2TNn4HYX6FigFabIUcxEkrc26DWOLsBdNMu1FRhkQSMVFRStA0ClpEB20Lr
FygGq/ZL29Ym2bU9ffq028+tvOhfUjDwuJLedPy8Z2DXBhbbz1wfT49rzpgGg/9a
ANLn44/WolEZb2hnLSIumBhdatlftBpyqcgQzeBFmGmQCG2ikAosHX72ABAPfxsM
hqWkDd92lyRnDJfxO8/8cTPqbTt6/nQOmaa4XRot7QjODFa6GPeBywHngN5t8ejs
FGu2FSOCXaRCYtfo1AEVZ3kUlsOjBjuNVDZvzUA20ZGnpr4rx5pkglaRtpamWGcQ
sflRTf0IE1KnrgDHtXVz2dQapUNCrEkiWWDxGXOBQA5Xrn9UOchvr/8d4M8hNnvt
SGFx8DJMR+WFbBI4wI3rjJtq8UUe45Bp4cEgQZYGUGIxLnV99C70di8ArrpeKOrN
14aa1VxQ64h/mM7oLz35iO++X/KMXfwoZfFcaTUWe0SOceTmq2lk40+cP88LZ44B
mpR5olZft8GahA0w0LqvXyAPevfLYoiIkkgNuOoeft5IE+Isz3c5cyd3LlgVPS3b
uzouBm3I/naj0stuC5eJBmXAN8Z+QRsu9+AWbfXuOmKrVW6d7g3V/dZzhYImnMw/
w/1zC1OygsBJo0Z9NGsHkDe/fTEbIlFpJUJBV/g4u+GNTMRlq5EPVPiD3YMam0J5
+9WGupjIGuSkPhabxVBi8yKVUJppg+k28Jz9aS1fW4AMq0HwX7oaQVm8bMbt5pkk
4VlGzWO4uyy4lHQ1tgwAlJsBjgIidQVO0F9DTcMF1UoN7XFzKNPErKKRfPrRBfh1
qnHAIhcCh6y7hXtwCYYq3iuqR96tV24ariH1eGADosC44S8KTGccn4yPNe2CFxb4
cCssvGDMmVJreEIjdq6vZU8HpnvQCSJL3qMUEQ8M8vYmuJOtJS9srJM8iy3gJmte
lE0gFg4E/EbPtkcMivvTM1qZXED6ShOnRDeL+OrO2wApRz4kKCu2GN3HgawJ4b3s
lqfH4JpoWAOhFquxxAt17jwyd+wIpLJZfg/Rpx79z0h5+GMrXMkWX4xB+PVEYMTU
WW3cbCy1yZlYMZo5WE8rkGgyErtO4PwuZa2uaCLaTRsiDZIxGvs04zlXp9Nwcs8l
Cs1gaFSWb+sJlw5T2fNQQ+Lnk9US4dHAii1ZmuKP/+VcectL3vDAUIW0FB4RVRM6
eETebxBtGHqA8B7cnbaIycsvW1JHsFXEqakD7Zr6Xe3U70LeHnlD7nmN7MP5UMqu
473zQWXxl9jahvDpyDifCmaz89S6rMMfwWGQp08vw3pHKNSFfym5zr0FDngrQ5O0
uIDpczz5bookAT2avJB1YQLPl1SAY4Zo9FwmRjCh7+2f0RXJ/mLamWSc/LbV2zlP
6eeoH8gp5BejBs6moOEJzHiPzP7BiIjIMZXfsZkytW84kqGmc2Hb6I1fYvWpr807
SUuh95I+gBmwp0NgpcxyIgKFr+W2/mtBlDjPeeeaGeVNfcDyJlbiUVNjNLrTvBHJ
uE5to5XDnXjJvTU9Oh9dOVqHGnbnjkgEs896h4E7mCTSPfwVcQoZ3qnXm3sl69Fy
C7e5Y1+3uEuBdpgdWXHg8LD+GWTCeQVRzjbHHS/9y9rHn2JJRixLifQYeee00UQx
8JOQSafPvohqsVRQgxwjcxTvYiobBLr8IBu2ztfTwpUgcI4259Y/WivbKaoHHdem
TcA6xsU0TeOTHj43OlmdEhyt4CE9Aj56mPMDlez2XTg9amvlAwN45cuaJkcj3s0B
eoAOS3ZFPEYWjCxFnQpOddFX6L2FdwuUXrdcMKdYB0bDIWGXZxr84jdm4X1m2Ny2
QLTlj+Kjku9K6kxrqM6BqHlWZqllXamzLd5msbf3Ud4pWrzK7to9vhH5drrTlY1S
U0TTJqN1Xn4ibPXzZJIF25wUa/jqOj0PUAT8CukoDi+mv/uiBlCXkL0taKaB6C5R
JK+mRYAtLeOXlMnIkzj+sG2HZUQ2OmQUmj8jV0euMvghQUjaTVOkxMjAR84J0Lsq
qhUfh9yu6XNV3CdECmDUbqTZHHPEI3ypwvcmGdVLbHedxpAzVy0kUKgG32V3S7yE
Nm2Sghlw6F1/s0M48Xno7N9o1gQFP0SuJ+MeivGyzRIYbzu9qYoutT5HfX1GzRsS
j6HoYOI5YH/7CimGa2k/aTwiRsRYo88LB9+5vJPKJw87S7WuHBY+uSaGcGhCPAKy
O0E9GjUARLGskONfMzSlfe99bePh14hUmmszzTbxgRCfr7st0YAmY3Uc4Hp4jA/p
tNj8FYdYF62gt+xwqoSeNIo6PYEXeVIDKyE7Kn8cXzQWfZbfgAbnL62RkjmChqk1
TkY9T7mmex53S+FJwkPTNrcQ2Hfavmcp9qy4yp4kwI2hGp4RUqRsj9V7POSHiTQx
xoLs7yIp+MS0hu07osFiuLbZbGBUlsqY2xcQ+8kuMJyv97njtRYY0iSMiFh0xko6
McWRgaVN5T6LrznEFZKDjfes7jh7vxy42WhK2o0tAkua8d9tW+1suTex/tDMLZpz
gqSSaJV3hVi+dANi614Qua5ZHyjHNpTx+5xPoXYEWbwvORGRTtuLqX15DifZA6ra
5lYLyWt3V8w4esBOz80fst2EeZo+bGtkw+mB8y1rL0Oh2w58NR7XbLgU68SAmBrY
vkdYeqjuN6gdsizPNQyhinfodi4JpTXK5GZxjKdp1AxBhtK8er2emzYl9PD8I5dw
gSFENpZWCHrdsLHYIZBlvkbFabP0HmeaWzNZtEw0ESZppsufkDSul25RwMTLQYLA
ka9wimFhpCF1LJFSxo0gkY/RoJrTR//Ay4S9d09rop6Akzbf46yWzFqBHg0/q6pb
AkSF6mjMCpr/1bwRzM6wpXXmQLzfSfV53+oafWFjliU6wxwV6s9IhcJVXbBfFUCp
n07wMMcmzogQtMEZbuc/dzjFBMAGFoELDLahz+015zqP0pvmI0+DotmtkDEPRau7
35iPSM+qrfBjWMiSyj7LhtmzomOfUBFBtke6SuYJ2cLeGq/zKxxDfdeMtoQsimFu
T8igqmosOzKyC8ogdv5Ex845d+840JvKlDmCtFNk+rN3i1Ce0Gd9NfLMJKLAClba
zKspYBiNoqNNOdTkP6Ha+WKAzhw3H5Wh762OfeY1+bDElQfi/InEkpFBrVi1QnUf
hqgQRpZJKcuVo1gsZQiU5M+3jSG4+v2xrKLcsLUBDoZqcPphhaKlx/kXAwkcJS+0
svUgtc6pt42RL4j+c11hunilLWKuMF50bnw+0rJKRWMwSHauVnswo/f3E1ncrwJN
SeBgI7drSipaGfqlpwQ2iL3xV0spNGmH3AXWHaG38j1B1ozUEWQnT/RAkB/Yl9JA
P954iRoRK1nAryKI31JHNpaJT83IxtvOs6nZNSq/1I5NLF1DyZbH0/msgvTM71da
9Y2NegYKZe330OvAIHC11ImZi4S657aTRuB7d+pDhJJTkSUHTxma+E61FdOUVSu+
rucQ9BAz2HemV/Y020ZYeGfkKRLuIxpcn0w6ivWwpJX2QscLWfjwqe+F0xwY3M8F
TpHUtVfaZGAaDEpMXvRnVCGc04QDqm5ZK0QEd52iPUKjMEQtRjgnpkFYxmmmTpdv
sqVAZylfPFVowH+iDIc7FxwtRS800FGPbb+K9k796JDReN3NuS3fJ3oORmE8RdvC
l4ry+QxU35o/XIGy2oyJBWjKryvh0/HCw1ifXjA21cH+a8VNYzjHgMGONBruKK7A
BJ/7iz5XKMLXUkTGxh1PgV0o/s61PkTxI9bj9cQcjioZotesN62EybNeftZxYnYk
7UgRLYyGlwlI2/87uELDQ5iaw7fNtz/FpV4wIDvFV0IDN8E2KGoQq7HMzfJvsXk4
tvSnj6Y1nq5GyCijTXWXXMvYd4OuEaYueBfzhLu+e9uk9H0CRNEBpXN/TJKxmr0z
dhIdiSCT6EBa9gsAgjIjYbdHTqi5tuNQmfmIWwhB1fzPZoem9Ax48Eqn+3WyZZdB
VbVsyMp1wK7tlg+hQWMLAyIfwQ0JFXIhCXj1cvW/AgCoLIuI2/xFgS6fIeeS8uqO
6YLhRCJYKkczHAGWcigCbXK858h+VpMSzYCbPDuzc4JzMVyjxR3ICF+BtA6ltit5
/xv7wWpfCgeAjkF6yj3DW1I/A9kdkLEDehb95USAbjEdTaWEgU4pcYfC4pfV4X+s
LeNoQHI2d5AtktjP50OBxjgwhVQErQd3qWbR3FK/neTtfN0d9ZsgkIWbatZl07JP
7L17VbRa2shsXyl934Dqs53rAeFbByq+BjLRpkzWnpkzQskTho66EH8fr7nghlV8
kqM7IT9fbU9asuG34yiFElnJeR/XDLbcx0fV8fvgj8J9ymtdLKP8Je1gts1+THEg
3jKXv2Y8V1O8s51hZ70ZUdaddq3vGi8D+f+XgazAFY3BTvrhWJuMRpIPDCi155TM
4mJQ4CYkbpvY90y0KAvX7C0T0oB9j0uquzOpyPuzHFdS3jgNMUX83AQZfyXG8WWN
eGxB8Pav5JrWDd5n1lt/k8jEz/ShShg/Y08sn6v/OM5TtredWz6Sz6zKjhIJ9f7U
he/hid7wWwqVFU0lLPtCOwmbOH7EazMHPuCBk+LS90RSW17GFmtkEpQvZL5HM10R
cl5Wr464hR0m3n9VTqT8yuGec8FDtDDRfsGQGo50fjYvXJM/2yz+uO4DR4CKx4R1
vJ7bQWtY5mlLl+6XwTv9hpWSjaWIaCkWxJp01CygbzqWlaLAeS5hHF1rk+9B8koe
+N7JuGgRU7YzqR9XMl6lgL0CuG0XEJxRQyVOhlv62st+K03YAJhmnwe+K4juersn
qme2nlaUP/JgGeslhiBOGa3hzaFRwSOUQ8rk7xLNSgqrNmMxmAQGRLLPB9pPdDn/
k0L7i02jZvo5Snv7srT6AB6x+wUyXP1qq+ZGCcPQx+QHtOX2ccA8lob3HCYZBZVw
ii9erDRl3/JGQ/rVgT2DvCnlqTcm8v+itekxtICpezF5MYBuI5dajepriA9ZM25u
u2tre8YEuvagM1un79JM1rlB6f0W8MyCc22wDrt5xo+43vAVlgrCdVX7M1eQZqs0
NuSyY0My4xEHMfT0Nso6XcyAWBEeSMhGNuBXKGMdH+9PZxTJ6szMoyoUjRhce87Y
edR4PmU3k8tIhmvkXapVlcE2oNzuRvcpjVRDDTP8X+Za05xstEIazsA6B7CDJ0aL
/lM131mYNijN8S2bdD4kotLPc18WDwxXfXwb8eGmHmDnaEUzg92EEWC6uJpmmnBD
NnwpaQd97F9oxsjkJHjjgtORDxVJKs1j8oK6mrnOmaCRZIig6ueCl9iBxxB2tVlf
G2vl4gY+FvV4sNwzMBbzT6jOFp6shju3rrayQUprNjO277nE+WL7zAIFbh71BqmM
jJ0325L0MZa7PLbGy0ncuuM6y9cTBkRt8cHm/KhHb+ftcK0/HEgNkDZq/6QPNMP3
VWHJeRoKJYp0Pq4W3rrVWh4WRGKJkq7H/9d4coU5dudO/kE3tGPg3fEZ4gsYvQ94
DcKjLDDVIzaa9P0Nxq1FALwyqCtTlr0U+k1pQE2dAC55h4paLc28veKE3ByJO4Sf
1KY/67Gd0+M0Zn3dUu+ieuEJ2Sig2piD8HN24qxTxDDEykRTNOio1A8qU2Z/GfcT
k8cP96iA5HAIlmoI6hnjsomg4cdwwnq8vYqF06vrNO+Zr2Mfsbebsb30qCiDubvY
7ZLsDiSn8YZJXwWLRI568kZlsrIgApTKas5lgAmMWdSGBQb7Hkgrux7ziVbdPJq0
9QcdLBrLKPXgDmnE1A/ltj0Ph/1blST6TtX6QYyHxxCe+gUjQOl+qqPf7U/bSXZB
nxBWrTX9rji8UUiaKfUaH0LA8n5Xu1q0NZVXYBis0ZrD2yECpJdtrC7S/ZSIWkYp
hmBQ9F1H4r3VHvXmMmVF6+K0JFZg+q+esYactouvxGVG4miaFvdsutuxBIDX/Lsw
26u5V5F+DXBrqXRmfVQ8NnYhwOrbbmu+TlRy2u7C9hLo+yfM6fxugGARdXNnDQpb
bH/8Kd82Zr3WtJxoUZHmpUWyOOz7g5K0Y+qMMw+EbiBypx1N6krXTyCaajDUl3oq
M4UC9ys5aGa7uKWQ8nNV/2BUAfLiE/dIeooUWQeb5G5o5wMYGpJfrH3UPKKa3YJa
swiaHaGliHnjEFTiY5aluwBZ3UbM+Q3PNT16sibI9PSy3GfvGx8LoSAO+v/xC89r
7IP08cULs92L8ObsjrSuQ182fC3Wp20QZqkvKzUrHUjxw6l3nGR8D+fQxFcSwCGi
Ddf++07rqX2EuJ0ecvpX5SeiLZ3FeveV/C6ErIdZrU3EkPSTHB2U9W3Ys5SR7cpt
HlAlGTDs5ZJH8SuSnraq4xpEbG7TV0+B49CnBHwxTeDteW/s8gV9MMD/d86qSFsb
y5F6czBFOCvXYmzzhmZie6h3aR/v7UtrXoTfJXJvZQrbQI4TNiSDfjT0PLi4v/99
3JBjpfjfYG+4ENsS6NXiEyv0VIu6dVIhIMkFaSuJZiLDWWZaJXYp8g4Dsxbqtyg2
8nnMAjcG2CWCdbkIGqxs/FN+Feuhbtdv+bidvRQ/OT8BEfySMYdG4WN/BD9boRsc
TUCV99UCTrMEMtzGp6Oq23DNxdn/5eZSdHpXdf0CX+1nEgsbj7R4lOBT5bIxhKVL
Lrd0HrPFpk96TEKovks+BIqJBmAZeuxDJfHQ3lDMI1jPSWyYKWA5vv0mirQQj9Uo
RUY+Lf7kAzwtYjm2lXvZ7s3HUDSKyce0nNbLgbqHdm9SMiyXNP+xZVtDeYwL3kvd
dRe5l6AQosDW9BL7x6snXnHhr0KSo4xGPTYLEaygmP+o+PmBoFLqzwz4URmyYaVG
Ivv9Npq07+Gu7CVIqsRa5R8TWZW5Y6jB5ppKeGQM5hvUBsAifUzW8uiL+jLHW31i
dMapIp2LePEDTi/6SYddVEDZDYul09ooFRaKa29eGQJuvXO21a+xwl4lFmJUSXtx
57diauBvzPw7tbYM7kkTz/BWU+qZ3h5vt1wbGlS1O5bUCUz+9uwBuhvW1uV/dKjH
CboUl10By4T5qTX2WcHCgiHK8wF3piiPeCQvwp8DyK4/0y/PUadSrq68bBe2MlAm
ff1eyMI86T3ISi+W67s8ktD3d+pN9F0G+pi1Pb1yixWBGoX4gRdJl6O6TQKU7iJI
fwRuL3lf2kmdayq750Dxma41w8mN4WXwHq4AHKgS2HKSOrvOwJllyRNEdKGRH16b
tgSqM1G2OUTHAdtayJL3OLTPiJc0MYHd5EKe+StXxIdk+F5oEBh5i9E0jGniMh7q
dPbqP4k6yo0DeIk9mJpby6DMQvu26GNEjIApZS6TFLpOysgUSHD1FdEXsJiyFjXG
qFWhWZkjLagldT+o8c0wz/haqVL/njYoQ+lCtxiEOpRMT/hGCcGLuTQ0T06lBEO6
6lJq/VexaqHXW9u9+gecl2lFbov1aiVeqIpbnaFe+EloA3l0rWiJ8DtiigrtOzJ4
u4okwVcjv2Mmc3K6ixYBxrhddLF0vJpNfgTMyLm0R5mziGKrautgqe4Huef4Rfz+
dLCsG1ZIk3qMFpEsbqIsX/Iwbx7AK77KtCknaInOyHHAqivqwqjqw4MCbN+GPFYP
fo15L9iJt25BXVjtCmpFT7/iMEuUdjm2O446JToJvykm//6setw92h2SpgtAMp2I
7HvByL5y4Jo0qJkHgyeVNph7Sm++HbHkdbLnABgixxstf4ynkfPkE4q87AlNxcGP
iJH5QH3JZOx4lV0R9S33nQlGGNdeXWI6IjTyzRzVoWoA9yBinSzZoLb1wyikpZC1
1tbRPxkhqWIxz+xs2meoptqyaOI3k5CkDsW9WYkk0BOYhQmBwteNJa7arDZl5FnA
HS8oxBd1chSyjboh1ompZXRml175t4+ChU3P8aKYy/RHdc+Wo4/nfFCWUJ9gw01z
JvtdzTsUfaSqSrgWdQvpw4D42KfxpL3cvh9/Sabk0XdGp06aJ+Xu3CcXkti3itVA
SOVbehEbsb0Rkhu1bihKtIhXicPF/p45ALT2kjZkS5N7j1CGPVze+ZMvWxltCDlQ
KRC0zN4+jUhKZXxu8r58WlItYdbhlAFZHhuU6w8QK9wvR2RlxVF3DGR3WemJ/Kaw
LQAS8paASpDP1p+7iCzdDlJRCVEXD3BZgH+u4SZCAiSKipppwo9da4cxPHm3R7eE
z8mBqR+4rhbqrWpb4Ix3K+BiZ4r21/JgkwpqxQeDb842VcnbIUwtREOobCY4WIGK
lliDAoa2kVLrLxRuUvqr2DFiZWBtMvIGe0J4Nvt3MryVAnEVkiL4dCfFd2XwxYnR
kJ/Uqp5QcLWADYHCHemOSVKI7zot86N8AM/YxLERQGD1bXJ6sKoVpb7i7Bqq9Bfi
dO223mh58rLiwaGawYlAASB1+8DYDBurS1VXmOYIZQVniRwwV5vCEsHSj9FtTEqv
y8hh18ejBJFzNviDDwkSEqsTKGdHLutB1bIYi0OGdG0ANTnoMCVe+S/XAJUa6q2y
utLHM1qlLc8ggjGIAjf+xC/i7zu9+RQqGhhtOCfN/ZUuu7NhKPR4UMpSSAdYXIOs
8TigM1TmqQtu/VCjCDW4dSiiLCM+WBPRLavmMngK9bcqiOlawTA4MxxvAXm2hb2p
B8pNpRriCpHiCdzzeIfe2ybQKOEea85KW7fzZcsUXvXENFZ4LM9cBIAXoitQeqRs
X1SdMsNgTGcKPFZ4pHMuWTXWFMPLPJy5MEsZ+Qg1jZVsCTusTJ234NkbOO/3eIQb
LGuUX8g5mlPVLyJiANBGQilplyAHfc7SP6C7vztRaS+D+aM9VqqXYny7FLniRU4c
DxE8uE6/pSzmJF9zbJaSkyGfdPOVZSsxBDcKmhwFDCl3KB/vfd3Oj/PQgHvkqQww
vd5wazm/q4byO/jnHiJwBP/Dg4JpMASeSr39M9T4L7WZ14uVVH/JMhAyzKNQoipi
yUIgS/g5eSWDVjFNvMvYqZhdBZSFcaK8JQQbOZKZYb71zFNGBLjLBiogXIQGzhBf
v0njEUZ4qLmSxF9n9qRGGYfFkFo+rBqJdbrrjk36hxobTzeVij23D3CX/FnxL6qn
GGqMTwViHkzhGXtRGQqxrOWFauTMdFMU8w0yd1nP1BBXLAhUWpfIHc0sg4SBmuPw
VY7gTxJufSl5NqfJxXK7/TzJcxr3RSkL3mU2ECDDq5FGI0wraoMT9koFz8rWTMqf
brkLH6X7C4QNLTgKCSuU6jFVE488BRPkFl8h/xDSedvPKQi3j+Mbu2t+RGu94yqs
hOxNvrIxW9IzOoY9J83m8WnM3+cFWm/dMIIWQhl2aoDPEbxwUMMS16CpTqAngIXA
uHJ2+4fEXusy1afLG0f++DqoSLuxAbklP6CE3VcIP/rn599r3h7AknIHrQ4wuQO7
ey6k5Anv2gJiKd3MDbrtc9d9fw9G85wayLjbtsdxqVe5L1kjeU35aD6GQVePXunY
D+ejS1cTosATceiubieOrnuq49WkCyi+XTEIGpekW9yNY0LdP1Jo11Xg7PeHjZPm
vBhLzHMU4I8Y5wuFEAOGEMvYozkk1/s6hXlfLZOHDHEhh0Ke1Oh1zXNy2YQe7uJv
+o5s19gD7k4uZG0TxwGxjZ92bcQ+KQBjrrRv4H837/s+Sq1Y4C49y+wiL32qd3/I
X6zEYNh9zNKlzeUtm/P3Xvv0Wjs7Dr8WKAbhRoEZc2qi9HgKpSM4gEZrdmKck3S6
5b4A3HyftxE4OFS50R2nHzhoFmywRBVyZ5LTstaay8Z7eGF3BYiO6j6OlDyuyBNU
6xKY7dFxughBKhgbyr0BW9QB1yc0nq87JgclMV+8PqMHmjHLSza8zKWMqEvIadpU
vyswOAlkaXcCvNCUPmURfJbM+1gx2zjMywTGSavM15YbWbOo4xA669sz7RhVSiND
9TzE9qRRVkGOwGLSCFP/9KsYZgvP1JSattLGRuQPsNLp0THQ2yWoCP8ml5wtPQko
grLKXSY3wGn1hC1EndV7nIvXUC23NUpaJQ/e0KhfmkcKfVUQostL5HrWx4wO9mcI
8TkdJenbLTwzgjWOJ42ZBzAzYS72P5c8r3qVRabqjM1yb/QLGcub+xc9yxOLzS3Z
7PLg0uThK+KSXtC1FL2ScrLcJNMaE6yKnbaOJSX34CI40bg4LCyGDnmE3Zw11Z+g
ST6Eoq5pcN7mLBBB4mKz2f55xOM0viJceYxzNgeX5WBO12PjOedrfic7OLwqL7J/
UXwiEPb0DVk7z45+bNhwV2w/TMlllwheyB88lXjJogD2n+aG1wavUYBiyOlXhivW
CrYVP56s+gDqFfTGgmZc6uVutRZTBztM3sqifthZUBlNN9NIncIWCZ+aVYr9Wdq3
Nxs4407aFuXNG1EK8QHoeU1KQYat0W7t7lcoho1fKfe/C7x+2BG0Cb87t8Kyq0+Q
j3wpzSaiMj4vF9swCAO78ZzNBYXMDbkbsGpkgU+rRi5lBin2oz3rcflwGIFJ+uKp
O4cMmWJUPA5N8sBELFjsEv8ZuLg8RUCclDnrzSAmR00KB80/jBuwVDZ/r75FFRvI
XGIYO2JO/uRLZrC/o7Z511P0SVFBFxfUkdE7en+PVmCW6b+XzwS+yjPcnnwjSU2V
QWCN17/H+NCyFMhS9O4aZHX+20qL8ecS9NCeV9YZJax38JgVL1lG4vzrIRp23VPU
4gpYS04Az55kQ7lrQScNervvW5/UlUlbsdp59tJig+KOHgrRwa3/19FmruGfwqDO
78txYasA3jXOrWV8j15vj4m2r7s1xRQe0lnFXGwpLG8pHcXPOdiu9p39PXJwKs8o
6dna5SMLNC1q+V52Nfx5N+lB/KpPc4zuw4MnKH7sHjQjYBdZDa3r1ZXb7vdfiBtY
1ExlDsNxts1d5Wap4Yh5qwP9doRO84FacRwucVrGdbx309E5SS8LGssF4CBMVW61
Nef1IsaLAhO0DYQMfD9W/HUDmGQ1fTzjU4J4cjntD6zD6rDc3KyK8hLg6CFJeQXB
WDbjirXzbWDxADvsIfkxwiIlrTPwOiRTFKk9WOZP/MibegeGSHz+3kmQGQwJpLYn
t7VZ6qGj/RcRP1eT4Z0DCDPBjNJw1FMkRggCx9uZQhw2LsuelWqu8X5MpfYIGpWz
YL4M3Hew044h9CSqzxjBo0IE7XNcAaq8pwmIxo/liufGfxLMNEpOn0uG5JZUMQv6
LPpBLN55GZ/uOmtj7/pPJgfqFgOyTv00ez4vizyMEA8vlqISQNWFXCWsh2FwCFkL
8bUPIPe08qKkpJ9EddV9QNrIIlkXMzdQ9Rxfya3utqOkQ+X2lt3Y0TXYKae9oZH2
r1jBTCnuXkTnLGqOBoFFEeDD+XqRJQDt7JZaWT5zAHBfxGAjDE/QIZQ1BbJ0ixxM
1ToD8Vq+FHYbkMqXvRI9Q4wGBR/ckT7LqAmhnNBg9dWCDRqpsv/SEii+AB49oYEQ
GDBn7qfwwgQfroItR4oJGYMF0uFz1kolOShX3miwycE52lawxZvDSDuiuS+fGuu7
MjYIQII+Uie3shid4Cm8t9KMQOEtu5ouRLGh78yGd1Urgm1nufuPPsDlpEbZft5/
9iU7Xkdd6URlvpqczZnFeUz0CKBJ7ZHu0c7/NEqRkqWL3YKbjXAgI0kKAteLcQGG
5TgZF/H9Ru44JHslyhxMS8H1ORVK0UCu5XBTZMXygnfbUioBpYFLR1ZcCB3aiERY
wwWCTVgDquy6Zsqpi65NUibCUILQIL9hjaLg1h4ZKMtk8T1RtPSmOOYZeEeDp8od
a9GltM/mc91mbW0PpRxhb7SGwejKLUkER8lioyVkVcrZP+Rgt6EuBJ7rg/W45kK/
6JbuS8xoHPkvIVYvScaqFXaMKISlY8vBv2WCToR8GAFcFP+HQaNRaBc0iRy4zvIv
4qwQmb4a5x2fxjJzdSp2tS7Auf5W/g3Mt2x/h10vn2W8waTfp7dI/tEU8YTJInMh
Ymij0NhMtTANZbydfq26xKLjXM1dXJ3KuvB8b62am0bwIP5mKjzpyqqpiuhSkSwo
GQ0WZ/NhenJE6kwDciNavT9zSvgWBJnYaFXDWhfhixI2UBSIZh3Iyti0D+RxlN+8
gVCtHdnaWeA8cZpUXjO572j+L6hePlR3DkT88lo4gjO8anPrg0mlIQrnC7LehRCq
aktODyVl+zY/BEWiRWP6gV7IUFrKpnbrUb7P2G58avCu1wMTvjqRP8WIrhQ+L6qA
fOe63nEVc4VeXHrkD9zOUVQ2NmnKtOsMks4pN9m5OJglSeIKsXp3l5z0tl8ayl9g
yOD+az7BgZE61hSc75sQ0CnCsQ8GGtOAcQIkLvBewJNIsVk7Sb7LaamCKN/MqZ/m
I+LgnKa7YGshHkg3vywSqVOlm9KEHU7fiA5hsSx+G8hq5SoP/6fPVaOvJoGXETcR
0JD1aVdsWUDo87b+J3bCpcJ9S3R7MHDWjibq3m02MsrRCdmESTSiJws0jpIyM45d
V0Hw5R5t8B1e2GEYQa3n2S6wo8rYDRHClXD06npOAGNMfXYRtgBVOCDieCyQVQ8E
I/R38Nv4hqyMeyRd+Px8SQWjFRdoOlsEwcZTzaSJCSP0gIHSZglgnZNDU/QgQ2Yl
17xSh5waLiUsxV+m9Cxy6e9JtqjVme+QK9c5ImVNnfCrNw9BYfH4q5Xl+8UunzTK
DcG71bGiRVn2ZAeUKDyMXWHn1A/JUCC0l0E+YB/u3vNFgxkB3JqMDPpJpMfPzPrJ
A5htgEFBlXPZVfLEgCWiGXHp2kdmGvd3t+xiErxva7TFOK2i5jb5tmEkhTkQrpPF
d+h39cw0lCuJAzpAUlLYnZDU4GU0VE8EH0hgWlK/UMyxcyuOKf/jVLNoMPZKhRin
WdyWMollJCeY46pq5sDGsMDrJO1c720XegLIm7uVmxL0dN7ve65ovXJd6V9ZV+tM
/0ABsWxViCiiaou8a93QpqKj2nympd14DFEcvL8Cy3bjfnceUMNFxCygg4SqSPPL
5jgf1udhBDgJA0Kd3UVv62jbpr6PkzVgIm1/WKEF4fM9cCwJer/W/6l58d+S73gL
iWHXx47fze4EcSb6gnhEPDKP9S2N4k7GbrNkFWY00m1iRpF1Zi0bunXl3BA5InCI
IabAkJmCIwRX8+C4YmYpe7T6QVIkkLK978Vbl3/R1GSfGOsw27deGVU8CueeAjum
NAlTocv+aqV+jbgtXqsoIeY3/kCm5Y76M7BMpUC5zEbkpSuiM4WluKwb8Jt9Mhab
mEUkvuvb7at6+yMENpvhwDKzmGWAft5dUi7jTZ7tzKltHRmERKIZcsK87qfC5pq9
hz0beIXSiUR4cgJbGmveJDrCKHuvLzkJrW4g0olpGXBCDDh5mn8FlgfEAF1XMWew
es1F+U63dKRcr8ks6s/KXWzbqEsuifYZVqUoY5ZldGHz6QyTCmmZBOdU+hz2QteB
hP0o09BLWiIpOgarp5JiCN1eTgyzEVmY+En6dH5i8di108Ip6YwTV5vCy8qIn168
594B81mob0QQRA/ng0QETlMs/CWT/BqLekTGgHUoXgAHiVIMzjMY6zTKn369q1gs
XJ9iLHo+2kECH9k90Y7Qex0h6olfOfhYvOWr/DdtgA+gZCImTKCn/NPNY2uiTFiP
tGyRbGzxFx7pJRgsxNFHh4gv9SSc+bp1o2UBgjuU39SQYHE+6UQcyTvKEEFVKMHp
z9xXvmbDY1Y2gf2rd7K6yfRWe3/yFQa/ZA73PeO/wxbnHMfCtvc8I87jWCsn9Pev
iLqHXqz68FqWqZtZMx0u3/T3US9XJtFHzYJuT53PI/KMRCC+VRYZvCmT6Yv1Or8W
aA4ZaliQIyJ2d4yffGmHAjex7jVR9Nmq6OTa5Wox8nK8AqziVRL72Z1VLfr1u2lK
gCzv6Ijg1wofdD+p5j7zqvzbBZ48b8soJ/RynhJjTusGrljQtqLceUUw+6HJHiwT
FZCu8cQqJjekevmwUuEc57aH3fxjwVrB6NShWddPA2ZpiB7PezzeVL93U2dRo65L
2FCyeG2Rce4vAJjIYdvfMNZ4k8IQDJJ7rC1v5q7gTQYCobQ0H7/JlvKKTXPJ6tbe
3aAHzTX9XsvV0NGTOGpSRV7OGy6lqfc23e8LtZ53RFScs9V/C3QTxm5GmKzCyYCU
PHw3/HL5N7pcsJfbJ+5JVoB/aUhKwpbbi+hqB2aNaqSujLqkxvtSn058ql3fOUeu
LTcmvZ184cO54O1sWbsllZ5kwCInshcoKrn5fGmCas7pAlU2QmLX7D6Jn2sNJQxr
gb4qC82TCWJFGipth6AdDm3WPp1KEfc+dmS5ZDt3X15PLQ6NHW88kKs60COgYMlu
TUP179b7bLS+8v0RH+jsRKjl17MhDdvnHqoekch/NJDCLOacQzYoZLw/PDOUnRM6
NXCtp3houiQDjYHVYJR2eCUtZTdAYhR6cqg0TaEPovjo5HeVmCfPV3yQD9F7mZXu
yGDrBC4VyV64PnJR2G1SKT+PItLgwEK0Mqy5hTPQROVKBBxivgXMqVVV3tRmj1MS
1v+lIJj6HYYlIvB/EF3SSKKAAfDkf84/3GBo2tRf4UXGkmjvT+fjZaWPmixjMQpq
IzWIwGHh9CHzhTQ6fpLxTgkDfZ1UW8Vn0LNk5jXEHMjzE7QRBLE2u8gcTW5aU33y
HRZqXu9SbOlvYVxOSh9BSPi0KWGmSDEmguip+Pq5JpwAAan9AfvStUCFmfLZyeb8
9PXBUHRvQ1DgsTPg4CmIvuwZiEYJKpX8zp+jDZx0AZ5uNbL2K66zcdsSZqoo+Xr2
dVqlYwPgFxlRaDgKJpe8v8hF7VLnOf55bTkcw7slZgfnWH1CuSYNb36LzopmQzUI
czv6EukA67AKnXzu6vaXi2/RoSqi72W44CMUL9UYuXX4t71QIUChPX1Zs6vn+gK8
8u4pM+c/Oj/I69ES7wsH7pyDpkam/5Rgu/xwoXz4iyU6ZNDPRzVyyacyBsmjDiJN
+1LGQayKE4pm4TWijoahPf6kY86BJrkM401uVxMgzbyPaXFCbOn4ftWWtVCLHqFj
EU6/25zm3PoRSoQhsz8hvJs6YAnUBHSqVhEG+ImFV5sr6VC+uLTmTN89rgHAnuxd
CCOuRVogFnz38SAM2VOByEQnDsimypQr4M3336vSyBYODN295hdCHCVmHQdf9/sb
B7xd0XY7aDZ630E8VFXiPFbxfRmavjgZQuOBrhdZ8wh7MuIzQ6pliw5KBRg5qiJC
iL1ZBytcU2CbClkmuZ1K1FSldYLOYM5QZy3R5dj9MbDeAoeVR1lq8S0lBWua4j6e
hDioQOxK4GhWfWPOuX2d2039jXrJi6wGOCPRIGYwi6chpeMkmgr6rPL4wndnhA3P
OoMnSfL0+hpVXu05gvEYc0+kkJaQejwUddAz6ZKRNv9u2u446P2nA1nO5MVPDBDL
qvurIDqu98t9xwSuMN4BJrVB/wIpzi1AKYOf+nFFYPX+eFf+viIAMOfcKC7gUkHf
2GOB6CJJlKeAdFWdxjoa3umdGBt503wJS0/kp2jukL1GAsitPew5Sql/7wnBcxnm
ihS+ayvt+SicrOOR71el2qajhJqW5Au6VUPGbtya+EnOgr5nh91Q/AH9MiZUCRnV
nokpQbBRBH3k4LIfvB2HVORYcBxf+GyhUKuBtr0++NRb/+9QWkdEjH29Wg+ltQAx
yv2u6FBkkiuJytAe3nacPAHwZ4oFVIkg+EirHlP9c/KR3XM6+0MLS6F/vq6BExtD
RqisBYo1jc5Q9nEfMQ8j0Inh4Tm4/nibvGLwkOXgsyvWIclFgO/1A+/Ua2QiuPt4
JFwzXPoIOHdpEwUaSmo7TH42rwMTZp1lYGugwboUXyJTHD5Xvb/ABYFnb0uF5Jnr
tT3Qfl8kgdx0CWiGsDWumqLOeEj5GH1IOwQ4tSB6qwXVnNvJqkWotZYif/sjbT6N
8MZ+KC/bsGk1GDMEi+EQM87U1M3PzwtuObRof+6mbX2apHQWleamAkz91OGtiIdq
/Y5Bb87OYDIhqoK1AFLNOIC0OrC62KZUFviKe7Y7KsOXsk707MNojjM8jryLpgUs
o3dp3niyNqQaBXSenuT648YzR50Oc6gaXUrdNWy13udSlNbVjFIP0Z47VlJVCzub
YcWwmWMEMz/6vWWW7NW2UzKM2ex9HWHCOVYlUvY6enA7/WbpqPVLf9cF8RoIvHy/
llJObd2Lb3wCYTRsUp21dOf/MT/wEwxNi87ux319dsZ5D5O6MAqKv7plhUtsdBEY
UOadjVo/hXoLE9xg4RQkimZiBUnAeIO3B7yac9TjsaF0HwSX8HwCiRtRWjPgnltt
oG2f/mZEltGL9KpUjn/E0zKoFCs0rutCeLI4j9lNrtBkjUUrfwBZ3de2uzbACwOm
dQJvLCUnucRWN1+pr2Ht38MbvCSnubOktEpMdeTYMZToCcL49C9ZK+t/5YDEQasT
VQfrtekgLNBcELrvuC/rrr3uEU5afq/rVeHaBiF0avLHkHTLkdZ36HGjqvsLi81S
qaXOob+VxLif5trBskV8aYSb0Ga5+hUfAVJbcUJ2RL202mIrOhYzA/aftylVitKD
RfRIC1C/us/Sm1g2aIX9Cvhv2vef37hWFrql4tJLxIZ9HOuXCCTDAGPlQ1BXciPQ
SYYD08SpULHHA04RprZSPPZGOGt7TekCl8tj8Fx4HWafldjwwu7PHdWiZgcocYKS
aLmBtgMwe5TN0inNQInv5l0W0XdixU7hrvvSyNvWqB0UkcgfmPZXseD0xFwMwbxe
vgddYGwOriSutUlHHDiawaM5Md4puUGoR3p1m7BGDc4B3iwCE3JYnpZ0qzv62VP+
RBwKQjtYdVO1V9f3whinqw19oFvExuUEGjeYUuVPuu193o4w8DinCId2SkZpsn1d
ObQnbAQzAB9XTI2RpymWeIxIiubjhvrChd23pKXpgtZcROaLz3j3zI9WIXwt/pBk
2Zw5/P/9+P7YyshiMPgQ4NMAcr7Wc1qblFFtCJQ6TUD2S4F9jPT6VnZ/8uyDA48u
PVZzxALeaLC+C7eyyqLgSRV4Zw6+gNJYWdX9/rU3nmgeMkqZ5FiZ9EWByBQ5OgEW
2blFxIUXf5wACMuzZknz1kOp7tATdqo6aqnEbSj7psRCdmapYRf8WZ6RnW3+IctD
wo2NlFnlbk4EPhpKF501oUxpIuabPiCNNgZ7P6V2f57YwYEjcHcWPljUbzeHX4DD
boyRK3Lq+lMlgo3pgNtPfIqUaUlwJndtpbATAqM6TEEl49qNO8loC6ndeJHsuICu
ES/GB+/vOh85SgesYbBMB498VTT3pXVOVo6RBU+YoPqAegodkYFFwegnjz0l04FU
TtReMJ9X0oynja/ZMEtePWRPCq6YNnPcmmVmehU9DL9oO4LVOcoszEenyjpX3/HS
yuDf45e2Cqp0N2A7QOXBB4WV6pzqUxYKVA4GTVWco+7BwI8bwO+EAudyHuf7OWL0
RYWQlmYZC8YIEvfpFGdKZyOcCeVQFD/JpKTT8ja4ZVZJKReMfVQgcq3uEcFscmQa
owCYTJlKjZ0SPlQTuU73DEMKTv0/waUEp4cJcSeKe2e5vkPhVUnFDCl9X6DgS+eC
4p58+/RlCE8LdRt9sPkiccfc8LPMkoBdB0yR1vB+sEuL63UKi+wEObQjX587JX/b
dJYMCJMtOF+A2cZ6ewnq8W7omviDjaIFCvSEIAl5sxfZxA9s7zCwzdIHjgz8lm/B
7/7FzbdSIp/h3OiSjEf5mfane4u3O6j24J7pSkuyBBGMav3awOpicxwgylthVgeD
VyThTzlide3qrdmZg2Ormp5JaDmB9RAAsD/WThxFF3rjzgxr0W1Qta5UwevXDA8L
LAG8FVr+mVh0lIKfGXQXF7WFMRWYzdJRhWWL6ynxAVLyfvK3a8ybHMyyH7gDvvxh
xiuUWmjTb+8DR7w7gpx1cle6ppHeqBLGuO+a92o33gaWGfYbI9E7PwPEGfavxra5
QUe22I7RS9H+vx2lPOS7Y+OqXXbZxgvqccuEClIpQdQhycAiJNk+iv8NNRQSuirC
TqFsr/VANnTcZZ+Ft16gFGExn1mWVODPNVH8aLYaGR3F6+gmLiuqEm4m0lqXyDUP
D1oY6N3wS5SIwJQcoi8oJAU67pBQBHpxk7Vd80cdhRa+nQzIflbx4Xbv7IXMfcsq
dkSMsuj+toFeyzLcUSbiWYVWjxvaOLzk6dW8+cjHtwO+2+DdbCUR2pyUSXQNip7j
kLokBRZxMcwVntWV31nS1kdVSNybHiGaH5AO/QdV/Z4XfX0ko+30FkMv94Gpz8zy
KTldT2iYJJ2h84vvNQMjmUrltqun7RGe6wDAze5TrcMyqZcslHgUdPFFKQsVa4//
xlTVGzqsbF04gA2/UygAVBV0336JhLqfQkpPnBVz+SIgFG37z6B42Z1tSwADv6q1
QtjKVeZ8l6YR8g0sFbK6b1KNNZgwjoWfGPv2lt7Ipp0SMxuqwmc+fyIRL/z8XyA6
fwCIFQs9IWjXlCdVf4izOAGV2z0zgs0cEfAeBccxJjF2q4xvVjxYsTNT5JbEJFnf
Hy1+TlRd6U+oMpjWrKrnv9h4OzLfXi/ZK9p5/NN5pk9ycvyH2tAcobUL4URdglAY
tJ4vOBzc+LvR1lTRYFckf3+kJQw/YRpW1KO13uncmTvBu5gfm9Ua6Z24JZ5wbjDU
3K7HxzAQAdveizQ9ULGkH8/DOkzNXX6iiIoqu9avF0TZlIvBv1A5lO7BVuN29XV1
SgFkSRVyZFLO65DI9dtmzIGhP6u/+C+GXU0Hc0FbRire2l6dF2DRlBY/DlTbf8BK
LtqDCRf4sHqkdF6mkZ4s7TSeeAT2EEPCj5J+O7jGOY7qY8wRX2KsGxMQ8DbiKKy1
tqyuzVs8j0CEV/5c26ZYV7dJZRdmnz+/W3dRYrc5Lt9J9IjnUNlUtsAiQXc7c+h9
2jIzC6z+qOCoUlJ1LuP4/pzg8rdG+kDVbli427wuO/m6i2vDuFySEG35XOfgGYpM
SgCXq343xqbQQ8IaLjg+iUfyBH7aKkNMFLZ3LRaafaTR4kF6g9lYd09c1ZQsFdi8
IvlKlV0g86Z126vTwxqtz4whyAAtICETPOzfkLAMWFbBYlig3SsRSD4o9Dj12+DV
fxgN69DT7FdPKU5ODo6+36jgFykxWYu6B7qc5DZg3qUE0n1hCHC/J9jnbVDs1STV
dxS1PLu13a/Y0cj2fUGTOFRDJGHC3T/vd0anzxS8kjLQAPTlONYySvqj7qkeJA2F
YlHGFrWr1TWzLvqOw8DFxAPeqUX04OcVqDIaszWzmY3pniFDkltsvbckIGX99EvB
lDZvDvcUfc1CliIXlM8YYkjhXu8pbcuyImcH8C3vmha65bIQDT/xv2DIJ/RZ5wpo
onP9iQMw9+wJlTRWydSsCiVxTybXgHqBJc09EKBfJ1XUghxqfNVfzMudyfg9B1vX
2EgdJBnk7b+KQp7mbnYbgvjIrM45FajvlJ3crl03RC2kfdABf6DF5kdQ8bnAv6jL
qTjVrsx7tzAGwdqQyx9tlbueGbNxHqlq8XBaJOF4YvnU/9tLy4UkDMFLx2K4PkJQ
BIR7bMLQ/2bJHPdzSX7dPKMq7Blo23tp0BQF+cJiQhZKJSftqD2QIlw3MCQ3/Qsg
ejTcSdfWy9BIN8Dy9804ASWRqJUMuSkcKDZKRIV0gAfNGaW62GJaNpUhU1/5wV5L
B1uCN8dYNKHiLjRCGHCMVfsbWVRGdA/gvX5nBmRK6fF5tpdf8MloZy/JXnA0fhEw
CQ3DhFLMTnicjspQSpWWghA25T+FBPFeXQaHOQ4Yaa/tu3Y9sIHKrEmVkQ2iEFPl
3BFmiZuNfVOPNlDKU3mEebAcK3x4lBjdo/m/TwPx2I8S/dBpaVssm6JMqA7ejHuI
62KQYkD6ZR32/5iZytCiGt9rT3EcF0/0cgiJLs3kYhbiSKu4PigApMKXbJ8fzq0F
MStFNXyB9BHej0uDShgB0CwdnA7b3h5Ng4v0fo7s2TBszyCUGCb1Vs41VwrwPF4I
DJ2jPY1V8+r8yz8xoxS0MZ731abWnpTDMCoPGKR6aM9Lbo4vFXHPAJFztFIDK9ag
WrVaQw3J7rbwR7/D4Dw4aXep52S9gKVhwYwQRXEFvZqtVtphcGfSJBUToAAC2MZ9
Mt9ZROdCzZmpgvLlw0jh3VSxQL59xdGMOZAuwtFzHomaCP/JiPYSanAsJrRyMGHz
1CmW5QM51Xzcc8WI42webInpkNqi51ty53B2N5y+yhML1ICQ0MVWRwi+sjVAnF+R
nRRTVjv2AGkROJvyNoCNKymLznpfe1x9rDM8N9VWzeyKE9e/WQBYmYLJHt0w3DBv
Wh1qJ1f8kzTj434FHjlBOJf6l6VH7sXbsPSx+WN7e1953I/st65tyA3oeL6xf95c
6Bw3ydIpSUl2HbbnVJgw6W1kn61Qbs3A36VhjnyCIYqi9/O9r1fCh46FxdCmgp1s
wLeqb+yPMDdzqudBiu58Qe0eFiwGUEtMvN133F8iTVV5iNTXBa/3E3wIqv+Jjrcz
00C8XGk/vaXsCbEZn/F/71lHbLxkNH8QgglLZ791Kk8LJsosIPnmrbjee9AdNMbo
I4RG0R/tN57C0whtEda7C5GadjAJiZcIX9xEzeY+4uQWXusrccz2ExvBkq/4dIyM
5SG4mFgvTjCApBTLnT6edoUO0f0iEdJURagMwJ0rVe/gQtmJMV5f18vsFyorNFAX
e+QwbCejSR/vvhVwcZRat9BY/uS0z8bFkfNt9AoR0NWM+HTB+9P7GWVYCdQeYSs4
ynzvloN2IE9Zaevk+t4tB6C8wmlaQqGQpwE4y0OkHbIPtcRrXpjEfy7yEwPHbkz1
9b1pjtKOB1M3x46rZLYwIMKukrmLm8//8yH1eRQFTp2DrhuRdbcA0QJfbjEPsbtt
72gv9dIyZjDPHkojRhiX9nwEEk0t2cCWDLCA+5qy2ESBtWW7/AT20j/3ZAfzGmNS
JuOHbIh8BMR/8KHmoUMthV5Psu26ooaoVZM8Z5IhVOaZ58UdIV53f2S8/4T3+lR5
FVoxrvuNVdbjpOB1VdKOopf0igqku6PgeMK6kHqcz34YfbbWYIjWhcrOYPoThx80
XmpKqZAiR1A3kA0EJik0fBoTvwP5HD68J6ZMGCbpBUZoX29H7IH/PpP+NCpSUWGR
dhIPbNaBAkGlnZ205n9DT6cCEjnnPHKQCpbBbFFOmA9wMbyp7h1Gvb5BeQhumDHf
60x2oRIr/jB8/GmhMJhguFu/3Ul9HqAIiNWQyBTJ3fr4d6xJ3tH5ar8KbQ4jZ6yA
PGY+SksllR7Hcc8UyL4G92mDY7U72BGb2QU/Wo2EcBpKhvYEJt0zbICl+/qwPCgK
jzRR+gwssobFTraORhFmdYhnh1X8GR8qCLUcV4Jxsggum3pk8+PfD4vvGhgjEOLs
1lp542W9PSUcEzbHJRm6/hW8qe0h42TRPtoyVvyIpdrWfp0U4dVDLCDh5zpMlgA1
56b5AqD+cgLmdEZZFqgud6QqRgVCNkcXn2nehfwdS+WBlCf8GSVDWlpzi5jHynp+
Rm7/fqXCGIZ/t3wZ+97m08re+0VP154id7kUD9BlIJzl6UkZ6TVL6ahIUF62cKzR
iP4iUWDhclRUjx73njk6GyADNGOiI6wEzJDzOlaIsxg7g20M6/4qZREb5xtR7mUm
ZPEI7GWUif1mKDJDIZI2jMAYIqer3Yqoue+SLsGAz8AJadm0fI39W2MbepxIXqvM
bqwDJf2xO/JJiFLEBqBIovjxo2+foT6jJboHAqUIoz7m8J0dqQzTa5ARzZ+bODSA
YDTTQPRBXrXxL+ltDKUsEpeFirxv9+dri1Cl8Pbj8R2eRWbmeMohmxiVSkTPb060
7AvZo4b4dMdadfqidWixn3TAsFByL30UB6TTtAi8NoN+oyDh6LMieHtG1u15M3Lz
dXE4PENklDnpjEHWfrdV3jfi3+X3IE4U7H/O4+EIP9S3hxvyYVgOl7jPqfD6uEpe
rSX7EZfh1a4i130kF59L2spWEdgIV9ivj/IkBjHMnwqKPcn2FRBQFFFg29iyEEIm
hdDy6ui2se7pP1lVpgKzFnbgncZZzZMZ9n3PKU54EGuxViO1s5MqN0zwI+tZj2jK
EXMwYcNh17H1lf4Adbnql/et6Uc8xg4b0IJppkRf5gSucnwaBN03MrEsGgI3FQwR
Vv3YYf0r9e6kdw5xjE43jN6M1ZgPQc4rWHYjB59VPGbkP98g+tmmf6u/bKHZ25ZC
In9QELA1OeI270VkEmr8FoA/ZpqN8UwtpdIKDNrqdOIXFr948iPd41BR19nFMbRq
zSdwj2bq3S1MVDx+Lnw5TMMxHdoaauRzNrkBVP2ufstYAH2EAGg9h9K8rU3QhWsL
UTgHcikRL18uM3dnwtogkkmpAaev00ZaPHM7fNyzMERoFwSGWnXnZNZscB8hOKN0
MM3seG4unQNNeuVLZRzONFsFHvFo39ygULTdK2logsUF9TFMFvMxdgxb5F+wGoWR
pQmE2lzmehCV6bQs+bMHSTyqGjNehxqscJcFO5xKXkMVdhhV7oTfVZ5kAVP+nQhQ
60/gq50yJmKL9M3NAeZ1TBk6PkF29i0F36Rcsfjv06XSrO0qaLxvWrBKDTZKQpd9
rVUhMZO8hYx2xVehMXE75H+EBAFtyLo+kr+4tExr/b3b1UcZpTPMC3icHihf5j4D
3y6ZPWX9yRryz/p7VTdDvdiLnDFSy7/UVfwQov+0YvPXyErh7gpndMPX5QLYYtJH
DOQbPw3Sw2xqljX2iARI+8nIddS7XqIvgYuUFHdfaIZcTPPNYw/lcNqULxtMrC4R
TJfaXvx2RQ78tND2uTSs2jxjzMYxAHQ6dgryK1gnUeaHB58HoJAfc5TsoSXBFlhj
j836Na5ZibHM7jJT7DOnA8qsYAkXHkfUZvRMYvg40+24Nrq4XRT6AwB0LOC2vstW
h0jW2kX046cHYwgF9j6huQKRB+r6E616zsaDNXxSDsx+sRaQwsRVA3JbKd5XcwtF
6jPu6Izro6UEFt1phVJhxV3CbwuENYUzKOvJryibirFR6pCyHvVa4YmrXP3tS2+b
GS4OcNW+IREn0Z2PY/IsyHlQlOY8e58OZuP5dizojCgu1eFQ3K43tXrKHB47Vgr+
yY5CTSjRFXxb0JA0+/iU6tbQdeKOh7SQbxiX75GEwFXmie0XLgLDaRbZl40ho4vD
8sBjUnnJKBlJyFzbHMFRJTM8+chJqZ4M5syqMgEkXSWzdzodmH7PHMCN1t9FYVqm
omfKXhb/RhBwp2zCjV0w8eTEbElvlXHOwlDs0BeQS06zQjI3pj9EVz0xDrnUVGCA
UplCSnBOI1qm0oZKw1l1F6nEK3rKwNPXJ34OK3+QYNeX8SZmehoLRFkGxxs/ogJn
lxdlvd+JAaAdbJyQIhLO4ZScwMwLmQ6WuReg0XdelraIZqUxsE0aGDWWpE8Sawoh
yVG6aaOzX7nfBELLDlISKj2KjoevMvP9Rd+6FI0GTTL9Ho5/rFqOnk6mERDqmFRj
Sy+mj1u/J8dpPvh/B32YNXW6qoHcG1Pv3J3LU99M5cpuvPritbhvt+7W4uY6HQRb
1Cc96jJG4pNs8mDsHDtzAn3uEf6BdQ/CIoGDkHgeatG53CaEQwBNT+q+9VeYcoq5
/0fbB8Zi9kRhVQeHK3gos35BZnQ9oaxrjhW/fDGShxh4d3t+mvwYE1jpmQ6E0gzY
da3WIpafKvxMvrnc6wJmgWJLf+UkHHf6O7xINQbTldi0Aq5MWKIO18iLSZPqLB06
mhqV5MKkA+m1ZVaHzrbdDMBR1+d1Nw8aX2d3eFBLXIsEiKdjBV715fviHC9ZNSrb
UrQdtUbwm7n9iHb4i9gW9xUUgTY/E8w0QSErq+HNLgLMjTna4eLPKFahKfbfbgv0
D5yGwvE+eh2gm2Wvjz8cWnA0j4qV/bZ0VchBfsHaAs2+juGG0icZLkhuNDaVpzmv
Srvm6dsOwjnAJgLNd24BbLTVAFN78TTkkJLAf6WiGkUvWcvAEQ8BtCq9VjvZE00H
yUSKchmYM7RJoTa5ZiX3Cf9GOpOfpqsYwsu8uGDE0/1P71RW7quU/oQFi4spFNPI
bM9dKLKFgDIFaCII0yBnywj+hOKQgp48fm1SyYUVFQzKANTZGqmF77EVgYx3JJZ2
YYbJEkssDSBs76b9FvGC69W4BJkucbGfU+JphKUuBsk4j1oBS3uaa5QBygEI3a9H
klzTqohjZK1ZXtosEv+WgFo1Ju5zvnotxoVtyzPLLMk51NkTOGUtWXbtE5HvuioG
Psjijm1FzcsWo+VtjBV/jeF5DbIYD9uIhnKyY/u7OQFBbxoyl2FB7Frqa0epgjJf
sjo1uov00kZom1Iy2DBTDAyYqH4pRErimEkCOWk8/V9j+yafcDB7XsfpQnz0q3fF
Od4MSjaxFARMpng2iUPIT70HY8ua6HnvHXU3PqEzG61xviuvBMqIL1z0m9W5AUIo
9jG870Ynj9bZUSWQHl99Ph+emBg20s19K2l7NQBhFa3eOLw57uzkxzyegma9e5yk
XO7HLLWJMBdby5WKHA2LwUWKng5TN7hKhQGL2mEbVHpfKBSGhVPPW5HqsKJGTSVZ
dE6rj9xcIi8NI/EuHBurEoO5akDGJ70KvEE4w6KtHMOZk2GcPxtN017+w0bFflxI
LLxuDuAWH3wjlTho3gGoyRVzpTtZF5BrvtN5M8AenDIwTGPHz+GAxYcC1XIAQhdg
pSmPLZEheCB25YWvDbqxozmVhJk5odLb6DqsK66F/0IOoO/YTz0R5SOLQALfTUlq
CKgcGgAaRDHUZc1GM2rEYe8esFa5MbbqVHwF/RvbOC6crNMAzeY+0CtoopHGEcoA
mAzDSjixO/uHFdXaf1M8R2fSX1Sy1vuJoTQrMGFNVlvJb3tLuB0CUHvkGf5u1JfL
Lz+bLfl++hsNUgYUyqaXWABL8Mqp5oM/TTUJcwOM1kAgRQLDGXzZyfEB3hKVA4UK
NBlSmEjGSCtNS2e946CEModb6Rveb52fj7jN4lGOMDrwEQTRul8A+Dk5+g1Dv7GA
e8uZ5JfSvdlvSSpbDmyrA2yPPsWoWvPxubuLvXxxwWd1cASqVhGQeDo86Dzxbmhq
QJ95UAy+l5YQKKEx2+Vf26f2iDZVqwxRMO3ymDpvlHjZQPBsfnNFj1dwGQAuyeZI
6SgT4z7KzpmNHpv9QhPdtP5BrOUfxbVFWxnnFQZU7Cvc2coD0Juzy1wKQulyR9j5
MAoJwB8YkIGdZeMsDjEn2jzb0TBqn6oZ1R8af8grk/kBT5F5NjpNM/klF84wwrAf
zICNaK2FxEuN/9Td3qgpVosaIMeyB3hTDhEbM35ZzchUj+NUJ6fAtnH6XifKhIoK
OojTT/nMM0gGJWA2WWRnUWRy9+dGw4gopBPzkFFhHFk9FGHx/iskBdeyVrI+24bP
tqb+bTOWEsE7ISkdmhqfDCAUyuaLRnO3JqcJ84byL2QBtj0qNvjlWUHSy/sFGCMX
n/RGvMXYIb4WIPzlr94wc6GOi4dpTrDHw7WKaHRgxcT1QV2g4zTX3bIIwl507/k5
e2VDO6Q3beCtN6KZlwTPMo7gV2up/VwtrAGf0kQzZ0iXsYVyWYdqjqh6LRQrdhQn
/AkZ33NcXua3l6IzhLsJ5S8xR6G/baa/O/oeFtX7k8fdcdb4zz2nWOC2kLWymtok
crJbVnksIW8r/hsx5IBBAG+pN8XfjWW0eHdiYjLjqCmPobiel1AZEiDzuA1CWS19
06rULh/mHpEAjxFOhWOS/rzn/2gZVd90i0XKaLYnFfMyZH22aLumZSjjXY+L92RG
jU/1+iHNOk1B9jVXse82L4gPXR4I6ZhXkacWdY9FqHGpmneXgQHSwP70jAdsnqyL
noNH+74fsdr9nUBFsQJLnM5Vg/OkiVVzuIEw1ZlTsrLdJZkZTv28rSWFQWJHlYTw
OaOJT0hl+V9tEp1D9I8AIwmFTUJ5vL2limly1VkLY4xSFKyRZ9vA0yR52JzAGpNu
kztQ217rGW1lxqrSYeme+CpOCw/jjRAex65/VnzwmRD3YHo5Z/8gd+Qi31emr0l0
z5E/K8/fRjvt7Y31ZxddMxpY77aewR/T20lhKE/oPN1z/E99P49WQNxhHB+WP/Zi
yQuxCC0Csu0A4LbeAOqVFAOTfJk2Z5+Mj7PTs2IrjMd5IgcnaETfq9W5+G1KehPX
raBEbOmWoh5uJ4GAImtyfb/jaoIN4WN/0D+bk3BYzH1G5RotbAzjbM5yFpxwAE25
UZYsVsHHiqTzQ9vweubZqS91hit8BL/DoWMbGrhxm0pHBkPxi05y5BYzyXvEwJm9
INpRdTVgaougCr5xXaY5C3hKo46sPM+/2hbMrxn0MR+6Fha9kkJ4rjYmkQLnIITr
cPR7Z5A2Qz8eXwyIOYDrARecO2EurZRTcSdNdULOwjrnMgKCi9aZsKpN95kthmg7
yYi/vpFNMD1Wv6h/F77NT3OoQGTsYRWd8ZcxAXUVSUvSqNUyrKxiGRnxb0JvOx2x
JhF6Y3EanyL6Z/2zMvut0BUEJ7j6ZBan1Cjq0RBr0v6JIkFWes5DeKPpgoa7wQmi
phxcHQZF3oeJta+yDGChVHw6AsMLSPcFg1Y/BeGGRPaSjqwLsHQ/EZ91Dfu/NcPS
K7ZaJAn5mrIL7j2OU5URAUkiLA0u+dQ+BjliMD8zOIOnMx3G2GnaTZUZ2MQ2Sbj4
LZ0LJnK4/T9Gjx+c4VjdE8aW+Jl9r1kVugrGSsFMP5VmtsKZvtnnX0srBQ7nhDZn
oH1vowpmrXO4+yhAx3qXyrk/13QaIJj1HN49q7ZIzRg7jsSfgavDMeX+zvKEiYEp
SB5eaYLAEuefiNa9lb3nnZCx779J+9aFX+IiIm0Smmight3vhc2sBH9SGYAECNqQ
X9M0quK4WhsSOlcN65Aha6p8zdtiUBJEEP8RECH+Y95k7XF6iDgwNS88cB0YqPs6
1XRH/QYi1I1K41y1Fx+TCTT27EIePPp8ocCJPyxe3CuMLoEgNnw/h6SIehcoQFkv
tR9z1frVWw5X9FYNySM0Qv2DNTOVHZeCD8XdScud40LKYqyOSthTQY6X/D7HqzT8
7+eVJGex3bVGSxPvafBOa1E0LnN3zpRL8zEmJP5PlUDf3rXqru+SQwFLVhBCslnk
AfTa2mzZywIQhFhAZWEwFVw2gaF81g9RoYcJE+tCKIfOXX7Y4r7IHTFplKPmTLB/
Lca7FHRsnGmAPQ7Wb49KM4RhYgWNuLZm0f+G9NzdRqfJ5mVZKAQU4gIrAhinMbW+
3Lyk1nfm0VtyuzNTfgOojuV3pcqQ8fLiQENgl7bc+hlR2WAQd3m1K36Hrsuv/xWF
yC0vJUFX+gvib8ZObl8oywR/GAp3I8yr6QvUNP4e2ix++nhlwHPwfbNVVAOUie9Z
qe8xR7kb4lLlF+wyuVQMTborLq4W+Haplj77BKKIa3qC0rgMqFQHyM1kLwpCZ6tW
V/eqDkJybozZws0wNpwJOQHBTX6T3XSE+c7pg+nVFH4PIjNz1dupeUgpER5ajXBX
3QXMHrWwNj90TK9qI+PsFAmYuL4ep3Rs/JBZB9H1VEvmLiC1eki7/poz2FIGIiC+
QG5u8w3/SpU6yk1cNEOFZchIB/ub+sLLhUmJy4Zay5TOtVOslHorhT2IjOqQH085
9n9HUHaASPCjDcqGg7iASkFdlJK7JklIgKoL1yxpxoIxqRun7JT84iTZ/92Q6C3+
DdZbOa1blOhm33tWo1TXdIzTZruBmdHt+FVzJhXalD3GgpQoKGPzEAIVi5cpJckG
VaiCYy/su2cvrZKIvzvb5VkoR0NA1v8EjpPlRrEyMB8a+HzcBPyj8ZbE8T4cTb6B
LU3AudADzproGV835qTpRuX0yEK1RdYxBJ3z2UjfEnByn0wDrVb0LSOWpIIPrdsJ
iQJr/okay+dqJuydTSEkCKMpVxxdN/KV5xI1TxNdZ3SdUmq+mVOVpMzb0mWsNPVQ
Bb6rAupwpWOpb5BlLCTe9VtN/3wRl8rO+ZXG13tlh7EK52m3+zCGDHKKliHRVX3f
98/rdJ7TmdSnQZnG+L4e8+x05etyHs4I1m1p02Z1m0iwEH9I/FnQstNwT5PdtJfO
HhDj9wYUfZ5C4aoYX7gfVST8whbOR0+umLbKLEwd480cFRdhCQsyE17H67Yzus+R
uqjuoWG0rMiEpVHkhkTbQkuiljunl9crUz57oXn6c5vW+cdF/HZjIk2xuQXMqu8M
u1TFAOMw7aoS2m7vnbrVpHDHZQcg4B1c56bK62qU0RrHW5vGHbLDRMYFS+pESbRm
0Bnjsov2RZtU9RgselVSlTFJqr2Y+BthkwMN2F+srgpS20M2LQyH+K37iKcuShw4
kYul7kxfabs2eC8c0i8tUA==
`pragma protect end_protected
