// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vnsVXKCeYfFsMF1dBJ3UPMPVf5lUY8DRnMFBTR45JVfUYpu/Uj0uHgR/fM12UwZD4wk1SW1r26ng
kVFRO4K61myBrgVS+BPRNJD2h+KlBT5M0Dh52zZSYzS5Dgp8bx6AFsM0cu/c9kXG/1jLuBSOwOX3
tFR+z/ftQbIbYc04jibQMyQbObrNSx07A5s425wwhqz1AFftvXS3XMTt+BacgtY+iVZ6hsGmUdN/
lfYZpz+OINM7jwaL0wEpK8zXvVU2d5WhYoHNPg37jhNeoTCOu888eFYu4kRKejQyNJnxueJ2AI88
dhUpRXW9mjrGoVzlwuB9dZwUWi2Ku6VtmGrqXw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9616)
mlQc1rXX+gKV+WW3x7XooWchny8sFi1S9E5sQQXSP55ZH2/BKOyqScHn4cuhdVCg/iSAnETUewQ/
VcPJ2EK2A882rconYPG1cGBP7+HSg/5OwnN+/Smu2WJZFM5ITRXEwBCvuEh0okQjr0reejJt+l9b
oqrSFlQDa0ul9C8ULYTmjKwi6r6iZpryM8yvp4kQdy2PM/F7pnk1olHDi1SRjCPRYxSaR16RowrK
aW14R0inzrp5jDao8JuYaiz3IUzILmTQOW7YBEUPDFxaUSE6cqZdfzkPIv6dRhsBHn5FYnzKLuNk
ddGsSUfmhO8gobdgKlD9nLduVj0QVgoOUd93NwZHCZzuHdSGJwSZ4xkwsS5aoPAlCTVtUjB5slmB
MAzIVZbuiptgUdUOKXdgi9B9wvB8xnxq0nKlSMsb5CnhtRYgBbSuJ4qi2nb469VoUlz0GjLIcVyc
BKypLOaF7qc8nLVgMHT1tqshurYTv5mkDoKvLTeFLqUomIbJgW1sTIikqz/so7pvSr4XpXW49wtN
xtshtAgZ7yguRYT/l+EkAWK+AZ/zy3nbHpEKxnOJxP3cBTo/jQZPxT2kxaAguwGOqP/pK+1B8gnx
C6NwpTX/n9BXgv73vOSDoJuhArkwR6dax6DGpesKBjluelW3UpCc4BZzLv9MWTQ/Fl9qXGOqtfND
R93N8hn6iAJkj2g9lgEFzkBmRcLhypEm/QeBNtIv0JiaRS6PF7HMJ9gRGG2HonIVkR/HjrpAwS4C
sDuGL+1ZDUpTAsAWuZoDW4hE1k092WVKaXo927FzuWc8agAf5YWAJmMtVDbCCAAST8ie771iexzz
ii8zckBljkBaumGzBJ5MnkaScXW76E/1FsHaD20PLibkRpvlVGHrHCo5W96c+QxlxuoVxeujP+Z9
iTcp190VN6QXsE2+Rgi2XtAjqZziVBSlCHrCXMb0XvbtclfytyZywYUYKQWEXm5ipCZdBbZnEvU8
Dgk0vMUnX1yNK6hfl76htUwL6J7+RoOnvmcVr3kn6feV1Tc02nnDpYwyB1u9Hy/UM/EPQNWE6loW
gLGIvMYxHAlzoNByyRzBhx2CjPeKDVYOu4Y2cjWPY0K065BmyyM5Juzd1HGd/fFcnH09VAIXWXFM
cSgmYBrqm9DIJoCpPxeqzfGv1aTtMbp61+rxL86R/FS0RshUVHgnAIaPa33acF5epBU0xHdkafUH
z103Apx17mxsBhxJG7cOjWk5dEKCRnI3Ww7a6nKXMAHfD4KD1EMa3eb5uewTUoaXcYwrrPtthSyS
oZmFJEKAMekaQ5sgar/YnoLaStV0pJFCAbF0/KHVnzV5yHgnwZpgQ5qV9nP+VjNYKaCGuKRHBOUG
gulNh+8vjU4SX11CMPHRtb/PU1JdtXa7Ycrd675/fzUE1m3Dk3/0yTSkuaat5njytwiaKDF7k7qn
8fgX0lNUkGWcjlMApZBuAt5VFVg29VuJTJG3jfvvqDLn+ajIL885VZcPVG1p+Ucwie4uRoXcbHqI
xGGr71OVJMZ67UL09+1O9LzZWU2IAphz8txzzpnjVRYNA89KzlnL4aqdvtDyOBCROPvz2fpuCfmz
L63NNiTnter3r+wrb43AEYjsSv4NjdAYikL7HOJFOU1/hmnG71ne+5o/PtK88etnARQCq7OZAGiF
cIIW3X8xHK1TiG57BR3p/76zEXxt9aMKXVnS5W4WR5FN56pahylNA6vMnxIe998sHszuXoZmbdHJ
/b3K2yhmJG84MLbe6uwhiO9enf5ou3ORDWAlBf7FKPQcWmofsH4FQDI5Nmxd2QMgHWAk3FrSs98r
HDySHd9UNZbGUtriEldEEINfu03jia3kAJAW6sJ7u+szJRvieU9gv/14MYiAaUKZpxcMoiaICIk9
CtLR2pOgrkmsDlEJ81HpSlpom6U6Ec9lNYuOevnBPs3RXnCyy/5dMUT9LPOEwCoomvIx50KZEi0u
BX983m+9CUTD8XqCLyEkhD73/rBI5sNIQOUn8w9Vpww3oX/cGPVMyHT5yrBGTYSWowQdyAeIYFui
Ug+4Ktu0/IoYfrzQFs6y3YKk6IoudDhqbkDYpa6oNpbyTq/sQwXIaTKPCjXvMXgJ7PhvcN/crLG+
lgFKF/MclOGpNuXmedfY263EhNLuiARwCjW2uC54xUwChxAdBZStsqU17S3tWOa+1QyZfGuoDnqk
Pt7cxUDxjVKVnmeZtcJKbXyznaN9MwIffrplMmYhFPW3jf+Y69Kk8EXU/L0pMb7+LHgXDmD6WtKu
LVS7Xh7epyLspnGFlSMqcqmjkI39ZsKv6bqpyW5KL1wNIfGvyU9WM5HkAC3tpxExv4PsgYP2FgBT
Pzj1pIzmfoXhjigoFIBNz4Xlvlb13zsMy+D+9i2dE8nQ0z5f0eQwsX66SCoNXWYLwfqoHylULEC6
oMrtrtFb8y8WLv79k4x1b8vCtgVCAOuDVmlNfI2tdWMFbjxHwRklAiQavVznT9ja3oso2Gtx2Q8J
ozwsHOvCZPhDaZ2ygSN0gBHFLxbywj/ax0wU4+tzNAnpM0RqJgFbi04HB45+2vXSVi2quUod8y/c
TvCtubXcGHRz+jwVJu0ICHzYPLGSrdkek5IKJZ4Oc0Gm8uIxT1FRXeY80B60xjG+M0OfzJlCHDRR
fIsuhX+rlvJwbmnAQWcfHXcNeP3FU3T1tCYIyuRu0F7DCiDifDqKU9l4zQqbdN+sdaH1gTuqCFx7
fPsvktB12gUOSVaL37GZVMyFXdEUVcQXHG1A0eru9TI3fW3brz3CwDPp3k/+xK7dfwP2k1eGd16s
imYqJUc+0D78yoL5w4jj/dpewQuB8t3ZwIWBGtPhMLMBLI+/llUX48v5e4kn8+3tw2LuJSPA59wF
iCqdTHehyywDKPxw238l+2XRGLrPBQEWI+rOxUBKZgMyBiUu/iQVxjjUW8+6PMM35TPcG6wWcEtF
hB0QE5Kov8+X0xjRJHM0YOG6lkhAgPdAz0E9SuIxCjPe3eDM1WyHANBoVNr8ENTWaCj+wNlq34ok
2ObCXM+MLn2kYhhDlgzzo9bjnpzjc6dqq65PsFtHOnN8cjVqYPeyM/2zwRMvEtgAU+QhqvC5aS/O
ponu+BoXB94Rju4rVFrdIUIawJ57vL9iTwEqMf32NIz2gXXZqndDh2M8fv8lLHk10aUf0q/jwmGW
TK7ukHNPKZL5qsLy+JMw9oYZcYp5NosiTm0zTsvWQ5gH2kFgmTeaF2es9LMiZV/3+HEoa3nzhAkN
GeJuI3A/8OOoeFf/Z0XQAcEcTwFkVQGhPLlz86Dd+LrEOPxu2yagVrCI0kX1R3SnoWP3ej2lWWgy
qryX9h6sShFGNxyE3f4RwaxmpegIh46aopjp5TddC6+PSHCrTEplQivWr0Iboqyiq16QGU6eCddl
Sq+zqDyo1UlinGnOtLIBO1sD8wFGf/iI9XDi+1QhYlyhdjhaMNy0041aJlNtFgo1byCpI+DgQPN+
A2EJiKth2Jp4bHQu8F7nrAPhSUjoiLxmtC4zjoSqWlRgkM0H4qEw4ZrHIDQvayvwQQXIpYr+oTZ6
ne+IyvUz2LT4EGrq6MXOmlFM/O7Q+bHhhSOC3fu/+5Nakep98Xxgdx28Siw8hf7zdXgLeUgqWBOx
3rQtyCppMx2YR6C1R/ZY17c4/ihJWt/EEQmcdbj+tm7PjEu4xTfOPw1XBno1S+CojTp5rX297R/Z
DHAUaP2uA4iAL4+TRz2q6IbehvYxWpDR3MoXYIMzdP4+bhMVlTF6dgh9hY77rU49VBHdR0zFlnqY
0c9YT+9WlQMa8NyzLqZW3ykiPM3ATnRlYYhNdKuuEPvdynKNe+7GlWhqpHNcsB4NyKhDK/O1SMTe
88hR1e2ZD+RKA+mvF6ULegUoUsAZTzBO1rIHcioLeXkJ0tKDYg2B89NhcR3oXM0FGqVgA3TS0goq
5FcL0xZESrFIncfzgBL1eUk/pZE/LxMoKUuugwO6tHCRMJmjGuWrudKxl1NIxt3SPfHBqXGKfv8X
CXBS889+jHEBIG4kwPNO346oC1LlFGMWup8Z+pO78UdB2hrzzDL4tKA6mt4V2jaNQdYt3PROu2cm
VpjmPa0kyl6w1zJcqmC/HyCBZ0X3kS+vF1uDuj7Ku15kzYuDwjnbMMclHDfWha5I2Olv+65HOrSJ
bMkzRC0Ozcmf+526RhIS4Hpvf2sd/bAKdwAzDfcsBt2PVvqHacIHoJigX+Hdma+faFy9ojvwQCFM
yxh5ZnPMQZRXJM/ei+wFBUGtBFwisoDEiR9w4KSmc+1C1bUUZ0J3ziWMR64vaQc/MS5vBXpQzpyt
EMt2aBVqoL6/S/+ESOmrEeAq6am6vRPDQ+HMf8Q8cLIe0WmUWyniH80CINw4U2fC8QhmAhz/cfKw
fhy1HWZlvvuh4xj3ViNLTyr7xfCrBZ4KaHCtUS78U7a+FtgDXx4MrQHBJdQTkXmam7hUYOuRi9RQ
1PP0+XxGztf9vfU2Utc3Bre028rUIioOp6GYmYz42a1A0U+wqu14D63INucz0KFC9REQNaWwEgLc
VfECBHK2qsmpQxXxsSPu0j8DmRR01RKkhL8lqn8rEsctX/9STqmFRs3fUco7GMLvzu8gCDaJsxcM
aKJLocz4ibAlaFt8gCOpspCsA+i89tLEZNVlK8cbh9NxuBkn1AQtwthQ01EWi0f+AJI30fSY2JyF
h+pi+IRhu+7221gCJ5dmVGuZdJBU/+STpfhPcWWPsqbuwoUMSCWgU2yTllCBYzqd4qJK/xI2Nt/w
ZsTD0Im5A/MsbQHYrdgQVEYkY6CtYExe7SXjqug2gjizmCgXp3z8xGixCpzkUo0mlKZx77ZCDBCr
5i5IvEUGalA4aI2rCUMTf7GNypRFWF4jufLx1hnLi/MdkemrQIdc+0AzwMMmKyUJQvAYQSGqvhsw
+5rA38lkO4ACida0oZK9f+DxWx32suOWS1IfJF0N1erYPg5j4+KLd+Eh0ubwgtutjqk2Xmclhs6D
PYajXCub4lic3uZB+AZdOJa1YKICju4T7W1w56wg8G2xBd5hegLSGQ3xz2TjxK2LOWyHgxF3uqBD
q9NqPtN2+X1wHJQg185p6tq0jVESE1VNdNbIaHtulAvN8bPvcVCoqPV9PfLL+KhSrfk9ulBDRQ8p
p8Yt1nxDHTC6sp0bs1TS4ogd94T934Tn0dzCgjbPxF6CdRtyayVEh/GY11jLoO/7cGlbiWgWTWGH
4HieKCWqrtBvTcDFuttEv98LEOXJJYFTkQzewBeum2gY3YYeVG+ZZ8U3Hc3hbSW/Wr14XgkTYvr/
voKZ1BBcFDHB4pkL/V14/72VbIrVqBrFbeUxbu9KHWDU7173BNHsQ2u5qczav718hVSHjCf6ZFnA
a2y79cqN5Wbfw+gwP9LVmwa0663/lqoO0JeQdY/r8WmDRNBEMVFCNRR7z5LIJ9Gk7+4DHxIq4RX8
eHD7dDgYk9PGOb4Q8O9qu4ob2PrzQetv9Gv0lRXWpS8vuSW7UOElu+5Re6eWHX+cK4nxAfX/R0XQ
lHWfX68QPkdlf79i8dSVrOqE2MquotQdkNTfSMtPNiDhlz61xJTOzmlj9V9rzJbGKZoL4GaoZ6rZ
Y75yPJz9Y4J5Q1vtjqbykwxdhX0KIef4zA0RtzNuNhEAzKK9+VeLbnFwtNPWe1/K4qtuU6RXMFHJ
Rzi5Y8HMfUNHAfxkObHnTRxM3N/Sw8uxCgzS83wvimPxRiOVAYeCI0XKtx/r+PJyVAJ2kRdP9hWp
O861YIAIlEABp9RDuPWjGfmwL8k+vHhm+T+OZHTRsMtBdcMRA1C9vUJ+yeFe6/ftsyHgZiSXkH4+
WiQbVek+JQaljz8dEEwkU52+LFJGNcOL18y81j+z/cSzLzxgJQe8FrcaQZsfpVYTRXVEFzgNxRDk
uqWPAtgxBqDEh3r/a5jDW0izDZ5ryMiPJAHQVU4sTRug9tnT3cwGDCYncNz/v3s9Nfyh0jAiTdbH
Mzi7C4o9tIu0W0YIhqMcqv+8Q08wK0FJO8Aae4rJt8QE5EOvTCFM1LlA9vF9kZcKepwfvUPOhiLp
N/4KdQ/1Vh0saPa4ICM01zAcuRjdMh+6imnczAEAB5peXg7917CQnYDqH27dKbaJOFZKZUwqAlma
4p2laKT7GqrBFOUdmodJMyJWA0Ez4jZMrtbtX0PbeA+uxlyLRD0So+MFMZ6K3I2JdaiauFG+2aI3
q8oJai3X7ssjLOAG5wZH/vyizwfTM4KvWvj+PSLDVofOW0k2aSnUdefjbdVGS6MOBOyHQqK0o+th
PWR4q+NtA51SMolwBScuqkQmVEN9TlEkvmrXfXhtPdTKZUKndifIIac1ZqtBkRUy2vorO/Z24Nu4
+Su8Tt5urz5ypgFNQ+wuYNFU3nLnZs3vAxZw+4IuF6OFWb8/Fnw2VFskw1VWfSrCU69xc0rkyVwv
Mfo/bsDk60D758r7tC4py+Rp7LywVo+LNs3VIVNm+vBSkg0iV5dXR3fRRVQo1lm41QnpU0w0lBRk
aBHuK2JoB8LYfGoVoyXtV6qjcg+/LxdqqdYy06xOOQK4yoU2sF2V9njho4HHfbBMT3Uf4ge7xOuR
Dq6MQ17A1xm/fPdJWQfqHbWhvTG4K/nqBrZuff0za6ZHnYajaVFONWD5CBMPUNtExSXmgIyX8r4l
7UWO0kegJJLAqwDJzKDSL/ovUs3J5xCLUUF+nvs3KfUFQWNB0etvXLz3BOrMCW42yQwwxYl+TpYV
bDK5EAuKeTjrJqJq7yBw6Mu5aqAzHavwtW8twhU28blXooiI5gWN4MXMEdkuqcfyZjofCbQErKHQ
M1DhE84oXe3oKTnfCwMv/G4lmdrx5+VJZo3OUX7yo9mFyuUZ9SidS0RZ1d8Cp5m6Lc4WYmom++Gv
k7rGsDTNL4VuSfL4kp57kE0sOyWu5KienxbYvvvoFonqf0vpJexQGmYmpr9+GpLN1xuCqIb/Fsun
7lOu+TmoOOwtMcvWVsWqnub2rKkRreV/owpyhOUUhZHrj1sAHUhTGJ9fWxYPEgVkeH3M4nli3PLT
zuPKDzVH/tEggKOqXg+DshPn0WHQ6E75qVlN+cLLcYNN6SBFPc5yiUyUkQP4P1yS7pjqurC4mI+5
R7m3kSVznZJGSQ2Q+QPIMbQRhRM5AGfZ/xmMHCLYWElREBRgzp55VEvP0+jhyXVa5dJBTi0pFIqA
EtvQrN1s1FXlZX1AGO4smRerN1uCxSsTqml7WULgHOjXV7cZWZyM+VEPuztDx+abBhTyY8l2ESeH
8EJR3eVRYqfLqArBMc5FpxlMM/4zqIi+Rl43abMVV5mStTjWv0E5P8E9IhbdPneKLT9LPUNqbpKg
JI/QD6J5eLxgPmuOFwoQLTatNPHCQ9tz9dGIJ3wpS4r5VxuQ8e/uUiXuIEbfFyJE6aBU0meQx8Ay
X1//qN2CBAaQMQXXOyzPBAZCe8IBiz55Xpqmf/Kf2PoWY8Rdg6Thuvwp2S32TiKB8tDFM4CWUHx5
SJsStFkhhTD5veZiRSnJU5eE8FE50Bjvs5tJENobh/E6rVyLrE7DctsihcsF3iYtlNQwVPh7XjTx
mN/Z74F1dUoZ7qhU1yigRBZAI9FrBWLA5HMK4PG4CriWVrrDzMOT8aVINbvXlvXQKKUWQqlzarBv
jqLtf7VSD9L9M7XCHJQZR4pyhiPuH4Oe8bs7/PaT66K2f+Pm5b/HtDXShcLhMeOTZRWeX/EL7UkD
WCvsOqXMCrr1CwB7D2Bz32YpHhV9XjNZ31HVERl0tGMzfWmCl2AKVvI544bEuXb3yXesJ8gwG6pL
dE4O8y9wFMfZHR7NxVirpsVEHts+W45sJzhBfNUET6UTH7BF3JCQSm3GulucpAiqve1IsAQy4buR
RQdB9315TNLFSQ8QyqDBtkVRNj4f/AeqZ3GnEr2g8TOR0IRjEsFpUDtQY/vNkkjXanqQj++zCymC
c1sf5b/A/lcFH+qKdM+AhD/YtAAd5Ure0WWANJODxFfptSM8mS5Na+AM5IVVFJ3nxEISvHBQMK0V
m96hRwwQLNW+ahBU0pmVlXmmvqpc5ZYOqiNp14dp3M2jyfLgxTphJVU+R0QlrJS8JAHKrBS/0m6L
DWhJdu7W/ckNW3fYjC5RSKXikxvKlfBWjyRrQMTZajOGVilbb7JTNtmq+7rEN6Bs5tFwjQ4cxD1y
L5owhG0VNw+D/PlQy64pyC1Z23ByTxSpctkdCK2hT/jgJVg3YOZVbUAY1F+5Q5+0F3JXz6AfDpnk
MYPpx7ZrWt6uzUCLkHcgWkV8tX1+vYOx1w8sA9JgRODRh3rTR4KnkHraL2CwqYw7u126Pc3U7DT5
wD/2+W6y+4uLDplAeEL+s8jglYK7RUWzDQOuwPsjQhuslKHlRboLF0zLCg2+EFiGjhLhTW1A0R93
vfQCbTzE3s6GPizswUXcdQ9rZ7Lf11qcMovP81qbYfQlAWple4NUIwmW8vQY4nQuFrHifW71IDwb
4Jij5nS7Vt+WXCnZtIKHfaP9eNarLd4I+lS7tIBg/fQIrM4CzM/5Dw+MuY0/KzT+zd31Uf4OK0bt
enjGWHlo92zbgrJPsT0xy0BWxisX/MCMMWuAMwVF5i+IlpQ0H9DQ/z+Ewo6glnqjP2TQv8R/2s+g
GU+cgYnEOqHbausRehRA9waEMNzf6Phe63ljNUs8hXdIVZLPT859kHuPzVotfHOXFHuP0fLKWB3V
aEBLpU8tISqnpiz15sQy/mrVNpwyzE6ALR1GQY29dIktDu4h9NmiuzL1ND/lqiT6rMgqnvJ3Gk6J
54giNR8as04N+exqghxag4xAQDGviKQxiogGLBo+qvCOb7P2vCeaMU8rA1TLKCkBAXxXiHtFbtHr
Znb3XIOftj7UVOyIYaPwSMRriZwy5qP91Jd0sFGS7TvKsnIyL3VyEUtYZdND7BYY82yqPgzFS333
O5RfK3PuiG4EfaqtVTl3At9WZzpcVki7MEXqVzRqc+2sHxuvB4VHr2tYzMI1RAIuqO+q7uoBe0jF
Wre4JJHgAZcevbDPVXUaoPUBFvzBnBa0QlQKParTAee7RVaH0k5WcK6CDWGmZlhGW4xU0vAjFPhg
kEyVhqkMMBCI4xUZGWL0p2vnlZ1V3OclB0UHnNAk/ilAKDkm/we5iM9h8+3q2F7ahJ1tjpSdPjBH
lg8w9qOcELrWjMwGBndRVVPAcitbuYbBoJZe+qc1b8NOc4BOWm+TxvEnv+d3SV1q9rq9EwNedMFd
64tZYqxTt8VYvzygT54D0Bw5vLXvtBbm2nKZyo9epFPHD/1CwVjLIcHDpE7EFgTDKPN6nkYKOeN5
pkAeymOG/ZPKToNZT2y+ybREC650tkOO7t9LPW0nXXymEww4AKBG9HwrRE/9XRWrxUD6n3Qs25lj
FxQIP6cASyNOxwjctkYLmGWVOzzUr+I99vvWGtW+ToqFPKv/tSkEwNAU/BRjbnOrVcfwR+YG+LNG
ygE4TGsskp0tEpVYYU9QOzuA8AW6M+9fvxIHFVCl07jyKON/luOvP04fADsUMNxZjVk6Bclx888S
Zo2VGqxV2VKTqWaJ51+TIQGVcAYu7c0cpGeeHBpa5TJMIs31mLJFVbPjobLvZYSPiaA1nsQYBFmo
8aRh+3q+1p+t2ckPwnXDG9Zm3CGcMgb7EfLRbL+ZqMexgkbBxdra56JQs1fs07kHeUSxfLKqX4gE
mi09cjC5ZcYsQXtATSh7HR79hCO8NRSyHGDkvWoqY4LtLhBV4fI7DASFGQiYYTXmnysG1x5ZNHdX
DlQvMqagbDO1VGilV3OE3hlaQU8wlF6sCRBLkX8IO3plgGObrbBm6TCSbM0r1opcygd+LsRj38tV
bI+06hRgKIAvR1Bz77PgQS6fINpV8fcMkf8sb0Pr9XKiF+Eu1No0hwr45onic+jSOB4q6QDN3zAD
oJuWAsjp7zIdemJo/92AQbS/0mdwR9LExQJ6KTzwWdZD32Tm0UZkalNztQLweok20AZcgTAFC6Ya
cy1MQpJfupQ6M7SGRQhR7p++AwyENfvtRO6tAhIjNPSagCQIQlVOL2ad62mggMu/BHpFrl8r0Tre
yY212a5ALxUJuw4pBLES58j1jziPQ3DYOibdDnCgL6Df0Qby+njsxiZmdTnFN5UYPrUotqRYNmUd
Hwq4CRQB3EMfRoUHos11gXqgytVF+l8w3RJTdNb3Xwhcifustfb2pLGWzQSuT2Q/VU5kaPv80PAy
xG3HibcpGQpAa8/SiJCcaycGB8X9YIIKrDqwGrPqU82fNF+FK2wry/QUdcDWICrse4qWEWD0NxQE
iKoRJE5ce2t6lBtmZOmsigNQab2g7kN5UYTRiWQgIAqQv9a4WWoMGiZx+mm4MRqP6/OHgAmxt0J9
XoYAo29Apxj6em104jm9Amp9JEJGvvIGHr9W2Wa6hmPP5mfx0zP/wrQlVEPggqb+PjoUd8hPG5R2
zJbJXPdyZcpSBqIbEntS4PWOuHDbIuNfDbcZ5hhSIyvimB2CSRba+nngipab8gMTVZnzar17mQX+
r6Rcv/vIZGOWYRf2TwIJ/LStz858DKrRgU29xYEcR1u5O8eldVjz2S/jPlPDxbjt43FXx+EFOmJq
gYpRqGhaqVv1tEGFL+KEXJ2HJ5/j8ZXou+9+xN6mH/v8hFANzqQvYtOBvf5F3ZQZ3JL0VXEh7PSQ
BLOUpzqvPzw2N8W7cFtZcwxgaJIgxeDPg8lyAWxPwnCqU2gmkIxjVHEn/bnEq9zLU+KPHbwFMWLC
YCjTuDZaSs8mw0cl8UQyeJCq5BK+r6CCPacUeJ/UoWC9RpzUuIv/Dii4Rt4K/MU92M950/6XvtLc
Mb6E0HvDdxyxzXeHYrO7ozwBc0oyZ8s4pA6myQv+XbsGr1TW+1m0STjfEHkPOsJTBXvluXW89S62
5ohh5sQK6y0PK52QmCqZyRohUzzmgLYjlpY2DSz+1rUlo/Ug+sU4UHt7ktz8Alaj6BnOey6aEJNZ
GgCYl4rsa46G558hHsd1QEEmwfiFyLjQDsbep43GngeOjW9aVLiFv8kZTo1araOEMSKQvIHnH7At
jwvWbaAr1Ce2g8yQznbHh0axniKkYTc+9RQ7NXUW3Vh64ohAcvFBRW9PisVucN67KSr8lA5306FW
nPjriToLs5rR052eehbe3v1LXX9IP6SgPuU68wCr21DlLbV5qJPZTC7LxO/ThFupvZ7eVU5Zbg9s
p+y/ayaewrliGTrJadpe1k9JWyfuzxG+4C6uxNN/z0QC3MlBYk4evS2VBDnjeypgOrS0N4aSub00
Xy6FsThXyVikzR8YpNHlMgNsyYyU+zXeVP3nyrAmXVGLjl4P5wnDhuy1W170rejt6BCN/qF+wFrD
3LPUmIbKs0eE1IsVOUkyzCBFJ7oWZsrTFlh2avBm/OIhm+Wc/EGe6d0JPGgTGaCBODfgiDNGmJ83
Ua0GUxYyH6BlZWQ6NEFF3RFyH/25Bfr2bJudSZrR/evSvHkHpUa+o6L7GrP43ytIb8ANoW4dwO2F
LsgFFbvrNUUzAkRFsTrMMvIqLngyh+uuxFKShQDqQ8y9kpG42c+ofDETroAhE3K08+i+h1khLD5P
AmQWhLLV8mz5R5U3PquehvsVhn1yixRwCmXWXUC+HTlDZWzG78WN/8D+Eigfrttd+A5EYZZ6boc5
okf6tJkOFyWPxZF4oST+X4RE2OV5f9lmYhzq98WVo+a6Ksrhoc5xlioLZzIsuGH4mkNddsOYGJRT
Ca/mHDkA+h4YGMhzZlFCFmKAPhpliICZc0Pj9lE+MmzsgJZq3JbGPldgnER18fcON6+G40g/im36
g6yVw/XUGkhwaztOt8daaSatzmfM/BwN96P33kP4VMSn7/hn4rtl+xa/VwrPSb3lNc4ozubQ/Kd/
sTUrhlJNSALotUt/lIVPinfFP/uTCNM/o08tLvknhaMKegP7ZEsErCoxz3wldeg3e7GhR4GMe6eJ
3Sm4GX4XBQJX95vNnTOcAe53sTlHKkg8dZyQqDhoCGr+7UXdtsRfzZacjTtiHrGmjPVNcQGieYkX
b5xxD0aZl3b/eGj3znnDzLm9KVdYNO9t/UDuCXPdzOwOJcJ9siFwcaLMg6rAKJi+8h0nYAeNt1P+
zDtj8w5W7w30a3Z3j6Vm4yOj4kIl69QrRApQkWUSdGMB+BWn01RgaeGqqtwK+XikWmkkNGjQRDwm
g2o/9k84j/W8s1U9xtOoV6okVTsnUgvVUG2Q6KFoEQZACNdpNKp7O5n6jP0l1JE9WsdqoT5eUgnX
dcDtJJqBxyByPbWjmC5CYeoYmAgfe3zVX9sBgoT01mLFg01vFRrGMHu2QJ2ZytY6RrT/nuu3RCLH
8xJ+wK4qLCKUYNODF8rOFtzvVg0NTuz+W0UwUr+DJNBfpXBcIFWNESQD6+i3X5m1Imlc3svFrb1y
hjx748LdCRS78knxWs5SxXIVmDRiHUswGKQLQnxpEKVoa/77YwYBMf+OFRLD+gbpE+4ZdK+jwAQb
isVjk7QFd7NQGkJZ1pRckaQAnbBHjV/Dw6ft/k6lDXWclnLoevXsZs17wnAl8TzhhXNOKejIMrHS
ZAkOsPynmZ9yfLkbFkmJ14LXFjBNpgKm58Wbw5ylNtWVMv+q5iT7M4KVHvoQ7XbEJ2Xn4UKQa+BY
189BUyMjOBLaxz3nGsewaK2zGyXJhpO3w695v1rt6qzA7O9r1ADuwx3y26x71Bnvo0oolpUsoq7M
sjALK5E0L3WWuWfcG2A4h4zUkzkX53b3Brc11XRKRgEtbimkvMlRgg==
`pragma protect end_protected
