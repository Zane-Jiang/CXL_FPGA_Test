// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YEZ2Y6KBFOhjOH1OIjbr0K6Fh018GAiFRFAEOBji/A9NX7oNbsLXlI58airw
5/uOUaIihxSbWoSNnzswpnyrRAoG5GwAy9yVQ1B+8h06LxsnJeTorxoDnGUJ
drZ9ltsK1IPyL3wKR1JDL24vPO0hw9lJj/e83XiTOXb8tuc5wohNOTY3YKMp
O5Hgbl90qBFK8d5HrUr1HTJDz8t1R2kn8QhuNZN6+l2t8NVDbVztAIiFI95k
kPnd94oNFc4EcWmdHNGqwQkS/4Ygaxo84AtYeN7F4vykVgGSz6490GIh1uSZ
REVDwSgI15eWguzMKj7iR15GH/hNqIhbX17i0tqU7A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DoBG0Wv4j54nxLys11DZf1vABLI121Itkc0SEsFmhgqE5MKKwZhW0bc+PPmo
ADgRGQG1cJC5rXfeaaQCVfmu6cdVxNoyFFlgLRoPTf8dLxoik86GTk7SDcvY
3AxTeO/KD2Yik9YX0k3peGuaiFVrHwVTPZlZ1Y6jF1RCXnprd81M8GGEix2/
QfdtybgXVVW6mKO+SmU9Y3jV9sAgoRuph7GxYPpD2jjxf8dTopvX3JThBqGC
gKQghLOh2AeGjwRSIXoWpCA1XI2c9o85G2tMLPIVIuESj/7FPvTG8hd0uowD
bKofIrYYGJR6koqQxUqxIjC3kAZQxlIH2Ge0M4+Erg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qP6HSHlWQT39rVwPhzwu92UMuwvSzl/OGUdy14H3OHd25pWzkMOsHdqEkF2j
79FV11cRhJRaF07N23F+BIWNg+ghnkwGdlCA2iAxHBLlgELe/Cy4SvcNc916
awvRFdWj4CToBPp+ul/nrzqmwhV1jUmwH8z3fZZDEQO5k8WOjGQIs0Dvdb7y
EwNQAaUDBT5vWuwvOAietgtodAkFBQ7/7EWLxRZyUp6rKyza4k/Q+oaujtwH
O2qZjl8CtZZ1snIxKXwZ+TjCRucB5W3q/mQgGcd+vfklR8aG8ZYHPzCAgUwQ
9QMUyXu3RlUpDiivga7E/QxDK0jFnRy4RCcaUJIEmA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hEcSWwmg/Z6PnRoCdBQ2PK9SMfeUfUBCiJ7xRooVWDZvvi7EApFbTUqZO89O
j7kmmcgO+elx4w0EDdZHvQRmsiG6KpWF0fGcsHip9avvZoKGJtZiR13onkNa
VdYuvEpOypdMG0rv2zHr653vVHSgL1196EpEFVhQ9rzsRBjWrr8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dPknA+8Nq4VRIOKVkS393ZgTorsO83MOg8caHZTl+6I/04qX9FeHHcqJjJwU
WvKDFZL0cVVg7SZwHZsx46d2OyoT8uJ3Q0V1KuEk9Zxin5jAYsnmtJLIMIGO
o7VqDym9AUxCPbMW7yU7v9AioGz1QmP8XwZHfm9aKssOUQAFB9zdKFTPPtmg
Id1auOcyCV9Ca0JES4lMAZxjC+OVN4Yfr5Gt0JNBM7XCkSIomsXDBCBrE+xt
Qgko3NPLhPCx6IRRnX4dODeuGJ+aedcf7ztyQUjnNlht9POCXEPPG9RBm5Yu
tAEEWIUKM1AV+JNLEvpfmKADelc/BLz6D2s1CUJZSb975LkUyDer0DFS2kJm
DkX1/WeGD2gm7VP35lyj0u3M2pxMa5GwHJONsqF+IaqPDsQkpffcRkgxxrQG
qiUCP32cv64gIhJMrsJ/FO8r077g84KuAcBXWSaja9VZbg9fy43UtYszE52Z
SacpAaJ1GcTI1B7bpF4Z01LHzBGWcxEr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fDRD2jAwdKW2XOOnMnNuUAV4GeoLjmsUlODusI6/UIxmZW1sMVQkkaZTYoMX
ViLQir976D0WL7XSmEOXzPycbFl1G8ocXypUv+i3c77IcHcfztx+DuKJCr0k
AhyhUeYlx/rZLDdf6DVjn6Zg4cFkR241tV6sQ8EDTreQ8F5KS34=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VtcQXCanpfjoqr1BXce1BLCSWvj9m/yXJCjTPr5FNXLtoE3lLgIzMrjOg9Eu
ASO38biQ8qQ2LhrXksHk+mWFPByobetAgjfCtFHXDq7x1bDxjMWPUXfKcQ7r
tc4GNb5MxhT/0lWCIulFPWCJZMLc2Kq5JSPAz5te9iZxrKMp1qM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3184)
`pragma protect data_block
oz2mnMEADqdNC6kPSrmcKduQHEo8RCjNTGCXjCDq/ksbdHR9qQDxhA0Q6rjp
7XI2vD5y9Ib4fJRahLD3k+c8CHwHMpQYGYHern+2SL9NYOKJEBCasknZvq7e
6eoFQAr6HodTcY0TIppKIlOezS2x6fxmjzYP3bVW4G4hszMejA3nf0ZP/Meg
ddashQ/WbxG6qpK7bkdHIqDtCCIpWIcaYkdPu+J5GE5FMKCXsZhx5xQ0rdL8
CKbbGBL6fKK2WSRyqTXnpJZ/gRkJQ/HdD9liv0E+RNuHG/ivZBRSCHkVdMy7
jVkz2tqVhaGSIBbuxA8AS9aljWJAIsnnXLjJltSzqjQfDvwL2VDfa1suTltW
iMQrSwljdnd64fpOpzYcEpyPFrMiUAey3FMn4vpw7NtmJa/1FIqk9ARv/2Tv
Tnw/ndgrVfe1JkH5XmhxmMjSI6wB1AOxPf945tocIThxwiIwADz1FOkIO3QK
Vo7n+k4QvHFehd0pGXfAch2QIEOnukrIjpxBmtsEBkjdmyYI8LZ1tv9jVQEq
d1X36W8p056/l9yjBMtrwSivhue9PZun8ksZkbtgz/JIauOFafK+NPzeqnBS
glQiaHXCiI3RgX5QE7vzTQDHMfW0ME09Q6topaGhclagjzcXyD/pmrF9VyST
OpcaWLrwXpJDzee3Lx1wmFDfku1EuSBEF8CNkC98mCG20rH8O8xf7TyOatem
ihcUAcTcZ+8l7hJm6On0TZyem9p8HCIXF/tWxEGOoebmnvOk86kCcMTTVvpL
rtTNyZypES2ih9Y+CNZEtvWZzSYufrg/VF0wsopl+hAD5FoO1P58pdduEtzk
JNwOE6oqT/NUneygQFC2pLXXWRFHuaQ2HTAsWdg4bI3/UwzQQ4mjXt72w9+8
Y52v4AQZfPEf3vqbjN1DfFO0H/hy1oTLLxi4d9WjlsZ3HB9HNoIdF4ayxupC
9W+ge+mq1s0SDZzyufanqHo1Zk/A5bbz0PSPEBoIAnvRJ7vnf6teQcBRcuSx
kQUwUqXL1ww46FDSISR3VnMxiDl//N2s/ULsTMqjuIqcY6XyQjXgkdOrzPwl
4bOC5qNOZ9e+g2JGInjR6b8Y1nCJlZfHknPu1NLig7BcUFvDxUQRGfC4eopB
kstBgwM0KblkZTRSjRB5dX+nvjgp/o3oQUczMVvOO9AVstiGa/M7X/oyoV/r
4rxAb6tHMxU7UGY8t2A9FpQcO1X9oUtG39jvVzxKaWt5dKKUJLpyE0YGTj03
07Yk8WHiut3jQGgA4clhdE4tPT61X5pLOC92+GtOfr+arWb7oskixbVtExy/
Bf6aJP8m4RApQg9OwqoO45wa7xDjSUpIlHybAjFy4M6Lmbp5DKPmcLVm/ZjB
6jZJhCxuG6jIdaov/f+aniUNbcJ5w7fvOxKhf3BzEaJYpqygPInzJbqhiOU6
T5e3/s634qGVEty/wkVEDktGbj2Ngn57SZ62sgd9cAeQc/nLpKXOZnjJjmCi
xKp5/OWcXNvMwjutYWelgLsrFgx7h9gtgE3Wn/1Fg6IGLvHWI8QReJXVimWJ
b61xUaqqahRcHsSoVEzt9cVdpeK0Rx61YCyVZLLE6G3LtdcGvY4zHAXJDAtI
EPLHZHmVku8wuWUqJbXavdU6ejeVMGHuHj2sMWBpOWbLMAMzHqv8E2VRHHn+
cKcrAGCkH8zJnxoQkyQ3CPJxP0dABIil4GBsqLnsBg2HjFccpyTq9CVA3O3+
y7r4UfctqCLwW5O9x+9OzEAnxKMVd7sju6yda50toS0SEAyMNwVXjiPOw6KV
bTFCMbxwwW3x7g2zZRmPW0HUETLLUYSq538Ne1nkUW3PgfdzQyo6Mdpmv4j5
cbXng8Ugg4h72rd3vJmqkY8M2Ef4SXQUowX8PMDb+jotQRE5uoR3mB1D/S+f
pI10KM6FqUFKit7rclAVLhh/xOSYVM2rIB30IpjbhMwBBIFy2lTACKnGqFXB
6OLmB6BlWxvGiUVbUf6sQQKrX2nZlgaQNomhtbwukjX7/2pJAaVmUiOD2j3G
/0YyTUBdoTld7VmzTAlNfNH81Wtj9MmYe8v8FCotHR/I9I7h1jCAz0+kJ4Tl
xPB3kCs1nVTx3z308uu3To0/X8lktS3RIn9jEsZYFpI+HtfV1mjdtd/2wqUN
od0BPO5j68YengiiB/fU6RUZtWch/hChdX3qmtr8ib50VlRz+u0D7Z6KRdm2
5tW8YiDUUhQ8f19aGXAUyLzlf9bfBn+ToKNRLcKvdGLexrJJOnIOI28AuU7B
PsCDBbHPNazTHxgcoy8o8J/0QLSPem1ob2VUfWppnkAfGP27Ttp+yLVGwAes
g7eyXvRR3ZxyxiEIS3MkG1CfXrKun1Kexq0vu2GF3+KLtCX+Pgv3WchuOmti
E3T9+wXUpjEZvhf9CANdbvVZ2+UpzaHL1isN1bIrj2dxHGQVdycl99f9AB+E
uWznpqJm5uBIRk1/6lmO0ECmInEH6MJq3nTKQ6xNJEIaeoYq2b3t3QeyZvbA
AxAqH6VrpBDkpMXeW6GzCBt6c9ZbtWDR+whISRO/8i6h6uwNKzaimvI2xAyy
zDpn0/20uQ2VRFiKqViqRKfEbxgcos2e43XKeHGGCXDSMNTOqGe8aISGf20b
lFLUago/mssb9/u1NhYhHrynDghXLn/3hAgpnfiomWxBRRHsiPysQwsy7WLz
ZSOeXprkuMlaWZUddiE3sNw/BPwxOn+MjfOQ867QoqXG6lE27iHCVUQQiuR6
rib3aE75hkUe+/c90WVJq1+SvuStAHQwF49xBm5d/oxW1Ot3+TR4v6M4i1Dj
IHutdNzOyEtqKaD/V2T0Ma3jaBed4bnu3fcDkB0rt4Zmv4AnJvUgWs+aBFnj
RAoc6y0nq+/+8y7tA924w6QLhWTRwB7Ylie6jPE0lMtmYsKcopdEd0fi9K4w
8CJ6XWKGYYTxrsRl7QjDBv/vCt/dFw5eBHjBOib1q1gSU2cfzuswxsk9Zlou
NdadsJx3f5575vEnCHGBQD+1mV8OO1WclvwGCJil+CYIoxWenXvWksbyv4i2
eNMOW+LUOkzDKNpeBIxSMJyjGnt875jo6W5Ovg/BgUGBk3Rch4uPrKC6MkCd
MMGjZlMBhLDS+l2oqfRve6Job5AA7Xw4fyaVsUghVOjchPomG/0z57kpCPgF
h6V8kX/zFufNeSQZNUgq4gkOjLbVAxsG46829IxHJKe85PmClbD+yB9kItUe
GOKftHFKEq95otwPRlFswGUbV7779ZxSj+J2DIAJY8CT9T53v19CckJJUcQE
4ZFcOIGcM+29sHfzUlJrUjjkL4PeBeo5UxgM/rapBN9TNP47zgSjpQvbF5MP
F58V6KkoEZPugV8V3NWHGhKsZZI6xiGw3hMOQ+7hAoqa/DJpYPtq8vFPaSLq
38ybD/lzt/dpjF91tTh4DSJmxC8WH+HynTmYU5laR5PM2Kbfx4VizBQkyRx5
UmgfQJ25uk+o3IZM/KvhyEzFiQoasPD7qQGDAYJVXfsFXcT4P3Wt5s3EEY0N
Hhf7J7qPG/18g95aQh+sey72ng272m5xUb7XckCP+KIgIGCNiwl/1rFlmsmJ
Q1ia6AdgOT0X4sQzzEcOJMvCDEjOR5WpklU+dGEU+bnp3O9f3QgcGYVJFwX8
RgM2ave2Xv4zqaRAbPjny8rE2Wu8pN2nK89bAFe3aDMj/uiXlEicXAk37jFu
qIEaLk48H3SblokdKWIJf8VSHRX8gbBJt2LhBuwF99GW2uQd2A0meB7XWpRx
KbzdY3yHHUCSrAsL8LMHbQczFSUwxyP+wfDuJF1HfAYMEYDBxxA1ewYUn1zS
7VOgqam3n10gFX2DZiErZPNeHkL2ScjrNuKZWL+3S1WAf04QtryReh2ogS9a
WbyrlGgcl51gwjljXEzcbmiWBEd9zmZcAuljHCPvKztlbtkqaT9ex3rWgYZX
nvhqvNFX2FU9uJxgWKaspljiPQ8xefvFDKyQhZQD1d9mNjTPhIji1d1/aBRV
yqdeooPVJ+nuKjHbaIOlcT62epJHZt+QCJ/0oFeUT4Hb+fLYs0ISKBwZNulz
KjSCkaz1a8JaWm2OV0XCUjn+coyAacrGCgVkKntHZf//STvXS3rxr/b9B9w8
48x2Fqr7B13ADEFO364PCItrMt5GPtkET+6Jzhb4YwOXe7Wp3jwkTG3v9ny8
LUmlRt9hbDDVrhsxZHqgUU4/f/O6UicMeWUSCq1mldHIag==

`pragma protect end_protected
