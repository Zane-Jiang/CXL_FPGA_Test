// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
RYwShzAQ3kjK2ewPpqYQ6j87KKNXOfpFRsUXsDU8rT72n75//mswjlybuTPFOoh3Ug3/WiWXOXSj
MMTOejG5WGs3Af951vOBoKp4z9FW1hwyc+g7qe2HnmlLPOs9tOI9FJXVPh1SoFvnBKQup6M7GMS6
MojGkw29T6UrOKnbYTfwwEoGFlZh7najnStSD6UvyPtyogmlfSHp2sd2IM3HxVtpliK895eZcomI
BTkWb0wAJqOI7CkhiTYBFM71FGjqsrlejfssq5fsh3geMEPx7QLktxAyupyKFENIE/YdsrRUuMgN
A7Qr/6CSdz7FtH1bb2g3LIVQQ2fBhqOGKjaXTg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
7gnpONAnSh2DPjonUo72InXvv6zd+BHNbd+KxW4cE1zNVxde/hGDsn24CbI4XxVh7C0nnpi4oTa1
gabdGsh4yJsCWIy6GW0PcFrc3KCtNwsiBz4L0nzkNhEvJXsW+XiKGsTT1GwY4cUtrQoey9e6DXYp
jZJY6nChogeiA2kUpGmtrKyksGXj3LomQw9iiQiL99dbNn6z7chioQkkiQHYfgQKceIYFwg7udlW
Zo53LCVGSqlurio6BOPdM0/5+N2Zb3yZkTTOF5qplBqwcQMeGDgDRu3XY35EoZdrl8qqdG/SWJEA
n3KnwD57g4HOZiI9oXuiWe1aFJi1SY74kNxzvnEH161LmYJcvCUw+h1ioTZnpnq4+l+pqk6BWsYu
WP/f+C81dBLGVxAJPOnC3ZITyy+UbwRqFccZ5Ux5H4a78deZwvxDIMkkjD1gUB0z+r+Zz0JVwp0P
SDCdR4wLL9AN/kVA0b3fmxYHWtmcpfk15yHJacqriCFU9Qqaq9qyEVSdXDbgsxCp1p6kkvTTfqII
ZLNGQTDHZ0g3B/4Kt5x2FBQiv/8czAFZbqnK8VlTqmEr8aZfzY9slfwFuotUhXlqU11I82KhAn/3
g6FmzbJQNN7fQXngfnVqFtc3EHhM1yKg4stF2GkSB8wuuFOKmOqPENHNcCzUUvqPeIxp7ds+c9z8
TRo5eJPU9ojNwk+XzwJt34nyAkQuIqyk1iQaBYgRD02mkpFnJ8Jxtis/1H/EYY0CBkUF00ugEwrr
rHY4qhuEJIJMvn2TetSq8Xsj8xYqa1W8ZK3xCkHcWin/vODjGm+Z/kZN8ajJ0V/LqzTH29dQB9+z
vvQYTXcn3gyVuAf0C4U8xfENRT5aIu034rIJwq2YyJ6s2r5RouIGV0Z/NdP7HnC4utsUgEJ+n6vQ
VbFQIkEeSmt2CX9yTPN+3WEs56u9VHQyepeG0EJ/hAB4TWaw6ctKBWLmBtx1IPoSwRDIPFaY4BWS
gfM6aLgfVq5a1uffcT4f4Vfh5gnn1D/HOlkrx0JD+jCM2+TnCZyuNukciscbmHZmNjpd3t0VimZf
7Unsz0YtkBlVhEC06xMbqt0Gwzy52pI9y+eI/60Y75y4Y3tI4xTB3INSX5We4V4WzsV+ssxi/ZTo
hny+BFWBXevMrbqbx+IPOA3AHoQaPggDi7m9tp+voT8TCTK8e0SLqS83jPlG8jV/UvC1AvBJcqEN
849YpDOO/mimUaBuTZvZFZJ+6gBiaZGn06/KxLpasQcVxAq9kDZMNVhgrtx4nPr4OWxbGqmf0Lug
j0MHxMAL/RI9bt5SLiiJ/vk53zV0I02zGQlgNf9ZwwCVC8zwlMUutCTpscW5jdNeKki/RowJy7mc
Uq0LE/wuYkU4X3sB8Rc3uEDz3m6AnmGYiZy+rZEO0Xz7kPiRFykZ0o4YtuLbnRAOdo20NAG9oPO/
s+jjuSupjDIVOSoinG8677W0WuNXaLUn/CvHsY3qdBVisybYhznjpCBMwjiJRdDfNY0LhFbpRaJ+
FqbRS/OjvBPs5B19RXxyHuJRvKrTaP3FV1yziIoIWFT9lKJ0jh+VCtwPuOViywfUF9IeWiFxzbP4
eAFhrftVau9VD5iLEGZ4GtskAdz41FxZcpLV0vVfmSCobyP3IcNY9+lYZTWTGARRAqKkuE+TC5DY
JcxU1UPPsIv3o257kLXbSCyTPMe1JGpd/3PJYOAXyWklxYuZryfxsw46cDuQcmpcgiJCmtusU4M3
+uNE0hkfQQ0nNPn6/kW/gdbtovalp2icllEAcezJtmW54Gr8OvNLAGHDNE6jA0WcG3WuqT7v/l4b
HsJKRTV23FfEnH8UQEpaidVHOuahnkosdbZcF7i/VqD/DHJMKLf4T4aBCC55QtfMWEjE5KZKcVr8
M7135pwXmIH0EEI1J9HAOQP6zJynh2Pmt0bSsgtIAUtMvAWIJOiZNH0rghha8hdscGGxi2Rw7Jgf
xVGYI5LZJckAZd5lnm16qPZ77VH2E3ztEak8n/tyWxxNOkfN44VBDGO0VfoYG6eURVpSEAR9k1uQ
wbVJA39mF7uaStJqVDUYTH8J9+GGevTZ908D8T3x5zn+tZjJGroU9L2IO3BwiYhoWSPcNfNQdjlz
oGHruSHoAAdIVI/BLHhNi5TMscA+X8SwZ3YbfFMGDA/iiEfPbBEGlor30QPVHRJ8CTfUGKnQXWoy
71SKPKElT6Wu2QVDz5Hcj5775IZxUYO8nqPT/wONbU/pgHMrjqb1cidEj6GxMl/JF304Dh2btgH+
9D3ZqLgZiWiCofEDu0DANsUCSTkVR1fkV1ckzXqTAE76FBkUfPg/nijjvA2m1GQa065bewLdduLU
8FThrHue6hNVtGwSXJMxndM8rPD28KrKnTfHniOqYSXd+9AfFA8bH5sf/fCvw4iV5MJ405KhxBZu
1CtNM+8nLhODmjfCj7Z8Jzw5j9uHW8pC/juF5s3vN9mRn3DpDbZh/jjoNBuGaiCT052uitMVFA+2
ikQv2wUPlzhDrpsvz0C/sfH9N91BlSEfqB7heg+jburx1+gFOfMBT9CQn78++UasMEkM7YgAUbkl
LM/fsb9tmnZ2Wisd0n6IyZmvJVIglWJI/2U54WFv+/3fjOZernHNWJTgtq6fPMIEv/Z38RPOdfj1
8n+eup+U1DLq573dr7ks0/K+CZ56q5PK6T0kIkQ6n5nhlu9BCYZ76sEEFhreWu6EfQ5YVPWhniyj
PCkKuHJek19P2kf4haOnRIWmgiG/J6PEvc+AY3xLY/F+7uM2FTWdzIgJ00lF+2VNO8m9pTCbsiAp
9fzihosUe7cN0fVkFg9wuyDe0btrmCT5CRNSmuqygOl+b/g0B/+Tf/lT+pbQBMulz5RtmL0yHT3D
4UFpwd4XEEJtDT67mNi2f+Tj7G8LoXcXylGbbIGjuYElGfan3Eou5bDTtYVPCDuCXYqVgBwQ5DVc
abKZF/5PUA5qYm8Cbgukl4fojJywR7+Sg6T3vuauUSCASSFBZBCryZenIRtGliFyrhIRrOUcpHep
pKCbNs570OpwNfV5ZpmeQ8Nw11O639noNM5IviK+y4vdRUezv8gvGnb7Rj0csQpCY4xJOhWjlm2n
4Y0HBA9qzjr0kz2uM4qDm/DODX5wUJVD9Ka6NGBclBI5kuYfUHHrSWduU9g7PV7pMHVkw2o9sfXl
cR8JjGuk1//3yWSuxV2Gi7fPOUld4yZ4sRl1ou9i82CyzFTVJ5Cdi0JocDlJ9xZd/ha/N+GgCpAw
RT77QjBGgXbSFXSIDNZTqonwbw9gBFiA/2dq4ZQB2o3hS9/FYsc8WMt22CAviUfGnCD81lPxFvHs
Fy+Jspo5+BgmhQ7ON+PR3bHceRDYTr70Yba4xY7hTqrwtTEED9xaukW+hSl9B3YZtPuLE5HVk/ui
jeWsal7Spt7pi3TW59QG/FRsYsk98KHzF3IHAu7PRf2oZM393fLnBX2f5OFjbesaVfVjUHSwltHf
5q7DxMRB+xy7MYmdM25APbQHm2pugoPl1df8E+LhWAF5Pmy+QPI1YuIG7jk1WTnlcRiP71/szISW
iBQHUTBomboSF10VmlRr0KfInDeYP0BF6hbpuiuQODBdV22kPWTabLuipLUCTsr7xWop3QxcETvZ
RXS3UGghevmLAQh4FGdaMEr42IosWz95ufNVtKYz65QsIA1UIjmF+KrLWkEla7vCPwonF6N8Rxll
Bz5x5Cu1lrub8F4wTcrU851MNqXgl0O8T9+rZfu0HRGcx7TjNjDYpo9/AsTNL7TKheDL7oyfHtAV
inhk/igSy1U7LjfVvxiPiqbO6e0qiBDSQm0f7+PJpCmkf99IxoCikduEgYacE5oEQ8gdnE4wgBoG
vEc7yG112iqb0kcKxwFuxe4ceA5EFFzX1oZ9cSMNf98100R/ytOzIQGQwxNdU2t8FbQBYvEf+aOb
QSPTYsu6hAq12Hp2Xp3lzqdoo8hC3NUkaWUwkd/JGxN+QcKqQ7izgtUniewJONO/G8cFd9GcFJLk
5DBMzHv19mQb/sfH5uXSKwH2YlI9BU3+hr98YAFBnwwWGnpMqeUUogclw7hi0JKljcRlkOywtszK
p7jTi7iPgLQvw8qIPda01X5kghvYzQhTxFrw7vThrL21CoVeQBZ2FhLHfD86ahTgYLQjXbOTytYT
kwlMnHXFahcH5qT7ZAMhN+OmKEzJzE3rxoZimdc4j+Ng2+1JN6ejGLUtZS/SvrO1IC9usp8UhpAk
xRkM7fPweJHBOgy8xjnxtjgDIC4lNsqyOblakrIP5XF5EZScZWAmc2LYRPLNz38E482BXX2sS3Lo
Uhe20KK6xEFrxzGePMD+UONFRDdW/PmZMOMLFNnby5YyRCFyqT0jPokSwE3REteCLyWVuOCtsNVd
VyMms26aX4/RF/vSpG6ykUFH6xvPGTXJHrYTBBnmeNz1N1LUSdRYdj9dU7zBApustcWjAaYs6Idj
KZinAWcgO6xAlCLiBY9J1eHKK6DHlxYIDgIkbunR/SaNkJ81p/CswRYWkQDFNOto2V5U4UFSiBXk
R7EFvrbB8FyccYf3vKPGblx/y3GL/uQ5XYSBPuGtO8yA0VHeiWU4W8u39Z+lckk2MjLYGkiwQVE8
hD7Os/iclvuj+fA2o22W3VcOuIJQT97jgpaqQ2ecXCpREfwM87OUHIsmR49wxUju61Xp6kkLQ2KE
yp6SqIP0iIEtVPA/T/sqETtjeI86uO19/F8B2miSOx8Qf14Bq2d1bYBP3lcYR9KGH89R8zB8BltF
O3QLpe+WkL6mlMqyP9IrGf++rS9rwUuX9OOGRK8aIYWy4OtC9BbKj5w45e4rxcnZ3oQqg/34LXvN
+YzhJUvy7K0+YyrBKQceZs2tdzT3ps1rqV2LnF2zynWYXxmd4AP0fqry+dq5vKtFWSB9a2F502Rg
VS5fK+aByYzcT5iq7Dn45ILeM0ypGT+QySv54SFcSY99bE8ENX1B/59kR4Cd3sFvBN6RMvqZjU12
Y8K4y/uqQjafkoibwTu2JbZm4OakHJhdW+wuU7k+0O0qXOdqRLaUrX9XwtfomJR3kKRqXSZj6jNt
eLP0hkktYviD6iTaJcSeIKiuSuuKjtlMzFLI8cSDwMvb8+wBFyrgX5XlLr8AHt4IpHjbk8ntzCUW
pYJglYMakn1tOTDUeSoBIJm6Yg/tZFc9A7JgqF/A2r3ReVZo4p7O2Wzwk4ccwewvkCCvF0ZPh7HK
sODQQOfd+tm2dExhc7mUzM8B6j/K2n4l8xY/umVaQbEXnCUD/JoA3nIy4bOwdLxVpTlb9u57MFJy
7Y1AWroYVxshtje8uvxwUZXrkpvXSt+AxikcihfW87uPWiGi+2WPjkma8XjqVTyu+b3wXHmtFg+Y
4AHkqJh7dFQowdnnnplqxl1/NCGoXx/+mX/xvpaZY0P0btMFu4GHRJcSxUUTJ4nNTysI9i2WI0H8
iJayn+6FLyy++RZRqxbnIHRIxXppZ23v5jcqmtzy2oFLnqpP+yzp2tcqc4/abXJrgh6kOs9ZNAxO
OF+8T9ilSW70cflr4e5JyJuSbLdnGl3nKrdeDQCuuQnqv6AkJfMLTUPAtdv4pi3psBNiKJJMrViI
EBSsd1MLH/NhyGGo82dR2rqy8eHtNfTf0NbJD8ZZ+VT8xfdnOBI12T7toN0WYVyLJDtJyxnQXj9t
K10zWJsDNgQ7/QxWsPasGNT98nThkgFz9Lj2YW4VwlH7GWRLgaMPPVJSYGrJdagdQLGg4fbIdKMB
qHzeBoX+PQPsWzCma+ZyXsatwoLVMm3TlkLCemhPtuEK4WDQNqj4l/h66Mn/WCt5yLyvsyMno9dd
0lM5oFCv8lEg0hRLhTQSTU+qywkmpBaFu+jHBIckmWuclZ/dCIKCaPnGDvpzWCYeoxQ+xIpYYcry
uvUWuEAR9QnS3gy66z7Uz4LBdEoE2hXuWqtPIBnNBVWWE6X7S4QYqMI7aiDeuaPicbL3zjx9+SNs
aP3ZR1/b5iyY/3TUVMXseBkYjyQ4exhFq8R6EbP7r2HeGP2nPPb4wXB7cotl5Wo86KaxC0+4sE4o
w3k37yn9n7PqpwyKGjlBKvS/VBCF6+bEchd/Xk80JAiRRZagLdV9SMYTa/XtLNFGPkaK/18HMDNA
vSAHUa7T28Pg3jGIRxq4zZGkL9bll1D/oQgEtD+0QZzxR6qju2x9spKwmTdesihwLOhf5LTd/g8s
9omfxOjk6zZDpBJcv8SWbVjA+xTG5f2pCGwFrDh82JD24YGqTR4DYhca2Zok05TmurDHFfpLQz3c
/9h9T51ijrPHITyxymqYW/QcszpSEUfaC6XIbGxpofhEySZb4ngHr8ZoMey+hN7PiJRn/9iBPWKC
HSrYeFraN0WAm/wOK/ifR6twHdkPC1w7exDNGCBEZOtys8rWXhdGNS8sU1GKSv72F8qB1dMDCd2q
C4svQIrI5mbIaNSEBd0nyGpuc/UJxJeBTVuoPB63sPsgCfuXBM+1nZEWk2GwCbGpRL0ZvVl+TsFT
gwvU0OAXCpra2j+AZzA5i0knvXpQKfWqJpdjLcjQnZUAe2pd6bqTws9+naydjAn87zZe1QqGNqlP
+dZZYJzhsd0gCZHVjc6vk5zKqbjkafHWCp2bWpxnszTPD1gLfkwz1B1sxBep0N8gIu5gqjHTfa/G
pwk7tjIsBGTVJUFgq/Nt9o6XJ21VdcWUM/QRc8Iq/fnyoy4E9u/2z1xErqaHYBsFBG449tMooc1r
qGeFv7h6vLwwMxSFNY0onw3NQz5SmdG1HYBqYYKzNHDxLvKrqb7IS+jrDl+nSJ0qtPEgXrpAUJ9t
2QsbDrJd1WGzFSycvOHboEixkQoB7I7Q55r9b2E2IXpej8WlpgvZjXDWWRef/smvWEslSefFPQs0
xn6SjVbRfJcc6Qzke57CZuYXcHbR43BkoB+nd0VTsbBVUzrQ+jKjE3d/ld0lAQa50xkjhj5f4uyu
DvsImdoC7aQRXxVv9hdU2XgZz11r65F1F0E0Pqu3Eobmnj8AwdbLVf741JrwdDRHmBBSN2FeS4ut
WuZKkFPOK/9ziZUU/of9Q9J39OTVIu5rSybcDlEtuIvKZnfPdTNfLT/5o12oSDFNX6cG4deOe3aL
hFxDqkU+4pEIoUSG6dD6pfw8y+1N0rmD+laI953E+ZKGI2ci/+ZrJLm3zzxWsSHHD+OrtQikEGQL
YGB0po0D2XziSc7xl0AtSr/tsoKjSYYoPmD5dX7qBZ8OXRhwld9NCTE5f75oqdzPd7FbvTdet+6G
Egkn4prVopHiL/zgUnnReloVZAdtHbCQbwh/5Ik1eBwgyVOjySDNgV/duwF7eskUEkUI2jec5Dmi
tmbbbnCloL1SVBPNfEr+OvExVGLK8csnRw99E7UoWzaJwrZHNxNTugATdz62YwquiCY93d0diD5C
JfSYn+4pZhZFSGJxlzeXh+jlEzlmm9r9UmrhRLIykq20a8HrF7nMfhq93SoASj33mf+z2Ssmgzt6
h+FL2U+xdUrwxrGzMMYAp8hIjaKKg5fv0B9Yr4xXvu0aYKpMdFkXi6l/raAMpv0PnA9HSiHHGQzM
s9+WTYPLYN0AbCHgc8nhyCPQPKTiVzcyy1eZxHA7zswjps+6U/ffwTde+mFhieu5Jq6qnfTfGjue
YT2KaXXgCr3eznP3zD6gAbHDYTXo8obB+PTL1E85NUlD5ikRLxzCKUmjKwSpjhKvLmWT3uad82Fi
8vz9ucfP0m/4H0g4L9ay3VtzGYNFr4dOfmK962AxAiVZ0yD4dFfRcCXvjePCIcyKgUalOUNdTxDC
rZk+WqW9DcNpznZSVuRu+YVx16JFqysw8aLU+ezOPL9jMR3FZDfB9fJXQ+FXnkNxKgp+tqSoSpCg
uOetFhn8uDuJwWXT4/7tyuZ1n1+U6CQxqCGoeOX+Au9pnLI+p0Iou+dnIvfkjKNZYKGz8r7B/U0U
0qN5pZqHqcVz3FDahNCZOtjaVSkTJ6KvX/zVZqf95kaP6WsNyDFJtX8dG+TwNQHYOUf3OErK9uaX
cHaryKCok71QAgrAiM53kXTBK41n3kh6yhurdrVFAgmwOWKCYVWD5t6yYbIyhbU26CMQSI7vGM15
+pWeHAa+QfXgbTiwdMv+lLkg2NtBUWNm88VP0iZqA2PM8wFlsplRUx69G99VBLI+4dZZGcXhJtoT
KrsoJptDEwHa40Nrp6KHXRFp/Kg40VajY4+4SapJ4bBt1nULqFj+9Fyzf+iqNilt3EyszxqLLxdR
U7Rr8WiLF346A/Ox92tCdwehebX18aMPoZcX/INe07OWDi4keKyKO9F08FfKlpmrkURQWLm7j+j7
IFTiPaMIaOJH54VzI2pzIh8bhkwoPK2+WSEdGFlaxdxiez5Bk0kqk2B+ixokUK88R8vcgY3eTOCf
aLbdfsG84urE2KExUS3tAph2QIuAfrqglWwe4MW9Lcoa28L1KsELd09un/L7SLXSYras6/5MoiNK
4yBcmBjZW7CT4MG0K9S6a+YffFDlxKh/KPm5roXr/I40A9cSXD+YJAarI5xaqSu9Fhd6DUiFBm5X
BcjbUb5ef/kHzQvFneQbOg5+vAziJFf463/ma6ScIp7w1OksfryWq3gfOcJNZQlpdkneDTnijVC6
siorCk7k6DWPRlTCmaTycJ5DcvxWpRK7w2iQXFD3BLz6f/Gofvf62Bv7daioaiVw+UNecz7sOCdx
acSyqjVjwLh0Ut33Iq3ONalX9C7CgxULYjkG07McUZ/l5mvb4vHQOo77TIPqpNK4zKh8Ol6ngld1
EU2b9/U4WEx6Trszg+hgydA856IONr49wfDWNpeaaL11Lm9THU8by6MAZVsYyL728MuUYWWAsO14
asnBMLn53QqxOP4eqKE77bn5H/YV4LVLOr4cC6j011gFk8ldu9yfmtrBa/aBx/s+If1m41akyK6o
d6w3moe6qdQjnWgQSMMaaNE2tMchm5cvuG9hOGiVXhYj+fi+WEKsD6K56RamiMinyKFY+j1n7GnR
nTxIiS+IRk4iQZu3+nepkQazoZt/xck+IxVpNDZVR99IHoBMQAUSam7wcFpP5NlKFKVaDY89zRfC
EoK8oFA3pV7QazKBYsypfvVwPmUUiYMAUZO+Fapblbn3mD0WfTlWwT7lDg8OhamLIqvXfvnXdfhQ
K2DDFKDifCa1s+C5KYdcYJZa/9i6aVK3mYTfkG+E30nPQldlD73NutPXWj/OiGhLuRjXUzNf2icP
rxtkAM1Lpil+ya/dhjjhc5tEKe7KXtxKdTGMVp3Wpcr87cimvifFiIfhU0F5JZQVt30UmE1ZpkSp
X8G2s7pu37UGG8ZPpG7QrwowBJ2qYVIWapRSkJpHGAck15a4Vwsf54mgRBgpYx17ikJTDO68cMpW
lStRg8evs/PAnh/jBdIEtUoivtkvRRTG0EPTsM+68IMfm2is117p+23nFogevCy6Hn1EX4J4I80X
1n78BcCsxAYkAxUFzWa9xwUXxpN3OFZKw8FFOLHMs0AGnlAgy5wHi2gSmn+6QUezzImqwjkm7Vqz
Vcw0kUrgQ9o5+1G6bpWoZkvCAbp7BhJkRpm9Gfihwrv9IJKglSlKeF9Uiw7I2vpYm0bdSBzMEa47
u+WwNRQy+oYNlpsA69tNcWX20VZntkCpzCY6FzhElOfH4SqLvPMafVLkpA+HUXd6oUz0DqQe9Z6y
Xn/ylGe5QHHXcDrNVDBS2omdEhjo7lANO6zBVKNg6ssnKdIj9SlGifE/t6q55XSTmlxh9F/wlYIz
akYFFMQJCcKpJKTfI5MqayULH4bMMNeIohcKIOgbh9E3s+RfG4tDI/iW/sZLc0NPzJMy2hJutDQm
qGQJ37+Iu5QnboB4jI/VJHQu+18BhPFKK05iy4k727nDba0caROVYN3v8ifs3S+VtHbg1c5ZEMlh
aSI+L7TmZlMb1w7mE4SxaOlShKZHm5VJ9zAAvdnGZPKO1gjfBsEkL5uIq7A5mLq5mTDQgW/mYtpQ
Je7Nmijjjr6DdVe6QeOTh5qkh4J31C1uMeqyhTnuo7ZJ9+EPD7cZoToHbo+0j0/vegJGfEAhaWV8
pbtG81KrhZjgCDxWYvBAgiuNkXgEJSpbGynlLJqyHEiqPT8o8AnbhcrYAkK566PXJZ9Mcia2bFX8
xw+m/MC8a6BJCzN3XHdRn8yAz3mg94bWSJ77BIDIJ2G254bfgN1710X8KD0FznaNIvqAn1WFD0Ev
nu2YhfbYpR1idYWDX8E5VezJgC1a4IvQLKxF0wjaNEMMwi5xNVos5N5CO3f2KM5c9tgeVevCPkBr
6MyzhIsCFZUkBr3z7RsirKBLJ79hXN0rROfYmFcBatbKcvIQt4AmMkNVVo+7XHqsQSSn/DlTpqSN
qOflj1QZ4Ms0cFkAdeOeIeVhGnFEC2XbqxoK6ESfakcFpq8QJNkZPbO11fyRuLYYr2GPIvmIB5GQ
rfxs1UJqmmTSUEGKC3teJL+/qdnFunBb/D4KfUbl371wJbf+G29mffH1/Krag4JivcMcr8/2Y/i/
4BGKlIuGQBphIWXC0NRjnSUUZypeU++0BwWkf8myLDnp/1VHOujZbgAj/S48oUpU/Jq8qMMcum09
oOgiA4Wu+7xiGD106NUJeBG06CZhMcMt7/E+OOgTWGrMtMdWlItADtBRN/+Kp4BWU4WD/jQ54N9e
N3329VHB+8oYr6H/NF7dXAi0u8c6GjzbxrYbpXpHJgem6A5zgSG312kInNgFWnEZQBUxHyugaD8d
thba/iwDI6jrsqYvVtnYPWJyF7K/oPCzwzHt34XWWczLUKg1n74JcMA09bGbD9IEO7VtKRtCJMwz
/nmu9JaVlFqq4Pv/SBernsH/7GDiw4yfbG8yDbmD/1I01kSGGR3k1hS4bxEDlyosh64COqncYp1O
EA7ZLtXCZ6rj27BrPQ0h1zDF93sbBKMR9t1bqkDec4CzJlyn579Z5jKWDpxRwYLH7P9gTnIbZr98
+HgfQrbPhLr06ulZUdINqWSamzB51XvamNt57tzE13cZ1+geuzL7wBGeeIUW5DbVf92cL3rxjEll
qOQOoZezYwBc+eDJFCAPDjMmp0Gn2xsu+63BO9SKEvtHBYF5ojITbUtu/uocRh66zejWTRDpns1g
5OP2u5ohd+GAxA8RjrD706BTdgpw7lfJIUaRPjgT9fI0hyZwGpbjHXeDhvjpU6EokW4UIb18NUAN
1A+Q+UxBOhuISLmEUEXsB0630I7785IrdVR0NIxLzISGD6LejIucgN26HH+4pIJGHH4K7l1uq5WV
CWu0
`pragma protect end_protected
