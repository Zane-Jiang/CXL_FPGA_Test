// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Ayys50UUVZzZIYxDTfmIlFyKl0xzqcnpTNbYWVevh9xOwESAk5hre2vCaKYV/pVPGsECNzuIvt1v
uPa6eog2AnqKd695w/7XnEisIwtyBW0hp8aZsqOdMVuIqQTKi5mZtqiHjf6NiTxd6mDDcABd02M9
uNu4V4PMIPf8iJXpF8G9PqhcEEK56y8mmTorba18V02ucWvCU+ZP6FznH7eFvcjKQ4x+NW8/z0LL
zb5BQgd/DRl0cF6Y1abmMhk1NUWPlLoSnZBX99+FtPsaDjqy+pmEqQRWNdWEXU2xEQUbiJCv2tJ9
vEo9zumAIlx7gRMJB+fSxaA9XLxOsxHfUHXHQQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 31408)
9uGS6D9+DaRUW8C8I4FuCuXjU0GvqY7q0XnjNRaZI5Ab6oUtR9DfCOT1gsSW30E7lD9DD5TIkBuL
N6M6LuxeVaUtbkxS7Fk88j+7FomIGnMg+u7txWkG0UAsZv/Uc0qMwo4aOZUN6OxZTh9IDcY/ey+y
6skoOgdIyrAiDgQ5avPrBnfbLzywz06wyRov3cbJrdrI4y0eEJaEYGFPyz2vhBMxJXGYlSCf4SaY
Ry0XRS9E39LAyWY6h1A2axD6lG70l8RDM5LlvsTRzVrQspTsoDKkAMgPBQhr/21JvgxZ2B9dliqS
7/vAYRUm9c+c0B+lDv3TPzMKVdqDz+bD+Q+Wda53qGf4bzCKAb6gi1lilrkN46aaIKz3yfoJYWlY
gECFLtETt2a6nsEBD6gG0zqYEUMOBLtRWzMuKPixmMGqM4U6WpDBtfac32vu1wyMvuGVMSwA6tNE
wGUiCGLVJwqftr1v7sOqdRrOxoBDckXnXMWa10TC2rtNbMtEOj4RVPBhWNK3+XBLjmBFuSg3EGuX
VgTN7jphqGGGBK7VF6qzi9OC5w6PmVtnTuRyK+ouK86KBGTsqSW9SOEiDGxc4Ile+ZccuBzGvjhE
9kcYWwKpE9uzr4D4UI6lE9/j29dW1kmrvsH6NNX/KXmZcjG/6Jqu0nS08K/BHyzizz3shX6502wc
+R22D/g57czbnPi4kkC1wuABnAiclli7Pq5xDmchL9qSFBclse3Ut+OmMOH5NhX0A1Hd6SoUdEQZ
PUSBy7uDcAXlw2EJm1aWkXdN2czvFQG3DhANfE+3HtX9pdjPQk1Cx6CDtCk7csGksDCknGCRY4Hq
z6RuLgDc7148MSip2w7ah+cGpFeBQWjgmr00dIzUi8w5pbRD7r4dtB4MKV0M2dfz/xjzZEiMdhT6
GmQxxXLplp61WBiapqnlVMpgP5/zGqr35rNnNCJmDMGAaK8bKisQJjxKxHLxTqlqJuzZkN84MyhL
Y03PWjMZWjvvHz+sSdnCOtM8f+WmtNZH/ZpvbEAU8nhZ0NvXdgu/sAzTIoExBijUQzLuHBHMsr/S
f/3iARQr6ny6UJpS+WDni2/Xr0IXFdZq44Mqqv9NZ/KkOyy8jr5uxykgy4tzgPrTE/9Xdnon8/kh
GnjXir6hUTFpjNHO9t7hCi3+XjLg/vcgDwvAp5Ku/4TNc3GJYdPgpwEzTNqLeciSDmo6rMOzTxWm
rIqHI4pCJj3AhuDkXsmr5wOjOSSG5obNSPIYmmHvJCGuX/X+SyH0a4pANShSmjjegUEA8Pi2Oqj0
+r+mlaJOQkjnhD5zUkxeOP3WP7l7zPYJ9/A5nz7y125me6F64gVofrluLuOSzssNRAvYe5HVcg0I
xBJw+UrQuylS/rKE/aj4pmqbixJYNJmyH+SMlYIkg8XKbFbIVTWPVO9t+ZGA7bEchIVPff8BWvZ0
/NazOBFb9jlCNw07WKVaUpR+9MJEMGk0YgFEtijox3P9IXE4XXkVIZqLM1qyihfUshBrjCuIPFJV
GSgHCNGIWpmPK8kMjqd+pUAq0JZdZtyXDsw4LN8O6vjMCC+OUoThkHyNRM1tEE4nyOXJ1UITuZUB
LBOyOMOXw3RP21dN2L/1JcDP8QV13lTh9/9khcoVVgQkumDjK+sEiH4ie+98VuLRO92fkBuWKyFo
/hMN8zC36oIqLhxS2m0g2QDVmguiy1lbJmNd+CxWL/414PfK27+p6sKk1NM5noiIll83jjlc+xFI
unyOeTBGDyAEnzyuFw99riL8xGpRDxJBomMUizd4uJo8WfNcfxLJnOfz8F8Xh0B8PRP03C5qGv78
WvAu/6QsjhHjQzATcWPIYogcSgIvNzbC8HcYDTdoL5K8+MSeHubyL/pqnow1aaJ7ud9jRh5QAWHN
kbJElYgiTFxn/xdCffizJJhG8NE3wrbaY0O1YyhGrCPChiCozP0bc2YE9QpZ0lxkbNfRJsVOq84P
Il6s6Mol39iVgR1CqmxruqPQTlkIfvnRAMvcOX6cr8hmIuV/c3UMeuSl2bp31EgnyNMYaLsM4Dy0
7FBTHyllVlG4R3CxD1Xl0J4sciWMt5fnIu78s+n78Dw2IUgcn69tYDpBqZz/536xFLetz4ob3Txl
/Fy4SqN+DCV7XdINPHT4piTedQdSKyXysM3mkzSwRF2n03206BdDcO1CXre0vFVnUXslsDKNX01f
8VDwFQJ/dm/wvqEqZakm3CZzu11DvYb/YpKf+JIxGYvi/ulzm9k9w1JPD3Kq/5fqxUADY2QhlEC5
/AXd43UZfTzcU8iO5PMEIfRXE1dRboMY8AViThGLGfmJRhYKl/BZArAi6TPRVQuZH7PSdOpoPSdo
OCQV5dhq7MC1gw6vgz1k2mWDIY1tNjkZX8RJ266d+V9O+jSMdZGXoHxua7OgonlgnngcHW17nnXF
FVdayp2+O3BJ/rfqcxvt7hMglT7t/fKQ+8Z92uCfw73tMiCdQXCYFP4K+8xix8HTrp9BMvA5HnMg
isbCMYGfUfn9okCpnRfNfEq1SugkwVHh/QPV/yEOYnVnWePRpxdfVYJf0q8CINvVhSv+YCjESJiO
f+O0jeBmTG8OsKNndKQhTbb5kLh0FXNArZkarDdwvV+AslpoU9knlZaoGF1ruByLS2fN7zIXc1Er
9ex2TQEa0pHc26G09CTn6eNWwndJZ7chZESSjvXIN8RYJETK95TH6SysW0WsZUb77P36rl1QHOzb
1qcM32AB33OAcCgZNjiExWpUJGTfmWz67QElW1lFjddg+LUmQyRCim+ewtzF74fatEL8vF4BJ8ks
a5K3k/QRtAgqv84DpYBlIOZxPgPwv/V071l4JZq/JxjM51NtPEEksrE4J0iIxQnC6wZQZSm+i72B
/AGO9oloDTNnmyK2QfVch8skN9maHbkv9k9jTjgKxfo/si9aOVGJ3cxgl3tWHOKQ4+YYeOOMGant
clenX7XKMy59UCFJ9k6PpuGZ2njBQRidkn6Nj29lS5PpJXvwSN7HXydDvY/vdrcqD+bRdkSCPg4R
p5+/MaPyAIrwxh9XM13lU5NR3pmzCSBD9a36ixVGDMGunr9dsGTH8Ug0TRcg+6JRobjQs0olioTJ
PexHo/ZJexneU3s3qVgdK9IaBWjtQ0XiNJxhrNQLaj39EmiCTqddoJJnvCk12t8O7C6BihDjAss/
6Qon/KkZ8yLOnj9VM849nKx5wAoqe85j5I+mGECIiWzt0tRdtuO54AfIJdSYr+nt4QHGfmfe2uOS
pMd+CNBNMBZE48YAfCTxi7EjcDVfUZjBgNjJpZh1T2I5cKJbvEdeNoJm9pjrc+mmXrnoyXQdtOES
98kHhj8q1QsapobZaCNisjvo0nSEUrSvr4l8cMbSgfbL0HyD1lkVfDqk6oKRgr8B2qdcB03aVkE1
GwYS0qVvUUjkwVuAc1QH/zHyOGd/M64al5wKcAYmh0zI0qoy/DSquak+DnM+rMlO5juTNJMF65G7
UvNJoWsOGkLZFLNjCHZxnIbEua3An5d4ZGzfj1pYL6lZdA0z6eirR1HZRd4knnE9Prr/ZxHtwvt/
rL5xR4sr5pusgkoRbaAsX28noQ5cYM5EXAUjgOO9gqi/ia6Whc/9viWjbF6oFtFxkX8CV4Hufof5
/LFkpck8GgfaqUTX0bY1uawf36gzkv2KKf67NFrzI56QvSi90GZBiMK19S0POK6ItALXc7FwOp4w
tM5sb4e1p7UxfNoUfKYfVfIVD3a3pJyeFvJNPobZ31wIwaYsm9jZOJve5wATBQKAURpgUE042UbO
H3JZH6ea/U6FzIsDD4UKjyFUWvWCcw9daRZvadVn81qffhLxZV44UOXjNFH8L/2swSYbNrc37Sk5
DMNI3F1yUnTGlsTR/ZbkCVLP9dSh6H43NUUBVBGCUA/P+AjOjIeFj+O+fOL1fUv8rzMTjXsvFVvf
iZwKHMOF/YtAi1sPT7tGFm+tTCBKG5nSql08ALHHjnisIjiCqwMcv6wpAP2lnPUcJ0VutGlZC1AI
lsQZ5cOIdHkq1U9VxZdQbQMJlJ5pgJiBrVxP8hNZzhBSXPgIn3x83LLBwoiQaJ6BuS4L7rvLmifR
CQDnnzKzb5bR/E0HllKC5T6PeRLAw1E5qqRmfvV9y7Q1kLibcPuObX1bYp3ZhUCDfrFckKiUrX/2
sm+UEnYNBH4X/rn7ZxAkcslr1DYn9fJCJWOatx609oTgO5ccmQCYXgq8RQB0gCz4dh6lk1/3whkB
KJrVJ/NrVI+e3jp5VxQrh+SFz9evtsxd0PocTpOxZ0i/w9H3SEM/8wAyoYwEKgJpzOhHl9IxO1Ej
8Q1PCVLhdSGmXBpyNTFkZQ9R+TreYYJVa9IB6wpIxISoAe2wPGYXgB0p4d8+QEXHu42/Hblga+8o
WoKfZGqhx+NY1Kc+2AUPv8EmrTQL5bauGQ03LgTpZuSyr3VPO5aQKZr2/DiAVgU7ahQ51psIPi8T
Mo2qTLBFjEk7+avVyg+WFe6AZxYSKgaO0YJRzNwQVDuV+UMNqi8fWw7/V8EDFZADT0FO8JFLqviN
7IzlL9FbdBBR0AcCvor/AQ01QjBpTY4Dq/5iv0b9cSmhd4sLf8BfuR21k+NUfeJJv5+2u2+1E2Lj
0W/Qaemu/5MLKgafBztWuXiMYvYxVAGYID7PZLYAIfP/X7Y6T3JsOLeHYWb7YIl5MHN3+8yMix8O
SwbTkGTGA9jklydt587toOAObSyEM0mLxTMjk/0Laz7kF/sYN1OGZGkWpYdousI6/iBQVOwJjVlb
WAnDbzuGCcAvkHWRaC6PNuu6U687jk+yMUNU+tLn5lipU3wev4qLa2JYum8CNdkBvlTZZCGBBAXU
WiFC3JA2LiCS7tlcJ9cjpqWXd9XsEoi0cFKGO4nlA+nGQ3jSVemucnbmyVejq8BlnHSX+GZr7t1L
+H/XwhBXKhUhLNNAtyqMGPNCZOyyDFS6RFaNa0UV+RhKbK/fRPX8IHAR1BzVZyw+jFYZZpuSDASI
rSqcAZnNHR0UngP7fPW0YkKMnGRTOJIWjBTGlYVXBynQE2gSdKvpD6kw3EGYWRHc+Hs7f3OTAnpI
qBbtZfzpLtr1mhS2w/IFF0PUKAOhwvrAlk1KjB9ewneldWz1jNHzRJoxfXM9CeSgNJsBwM7nMmVP
0YoxrsGu764OC35SnMvq2cl64iXvFuEqb7ig9lEWD/cwJSQUzYVOgGPziD/CLqCacAfXkfj4lmEe
Yc1wsqTzVstY0ryJnfD1U4GjTU/24X9kVnt+ZtL01GVXcInRG9ys9LSGMWkhlJi8jo1muhDjIoKA
mvrm8jORk72UttknahSByzXQF/z5Sq53eJ3/j/B6HgSH2EtH35X8D7IlFGee9726Nj4g7DaAAmgj
uG7EiQOjIhD/FdSTOZ50wF1Y0Ay1kVO31QbEvkRbBDdFLIfMIAe0K/n6MvSo+hJb/ySJaUAKJG/d
kjs42qudlXkW9LHnu5brcdNbz+4buHGqMNZMa6G82yvExJ6LhN8hUDMEX842An2QTQbfM+zhQUvx
tWJbRuvAE7VVUNm2udI5ggxHc61C8PnautMXe7I8sU73HIkdjCDdkqKES3GmufihYEHA73kGybNz
Qfu3r7/UxJMSB27q4llhbkLEiYOfZsZ30OQRKsVveDrx6XchewiT+Va4W72hiqGFbfItJBSG8Pri
OFUD08Ejqrh27gfZOMcHa7cCMDSXkMgxyj/XGfgBGFXt5TF5zT130yWvoWbXr3zZB3FEAlNSf9zC
ypukufy9wfgJPI000kxSWzbOGFpVn3UNyNeP3w9EmuvZr6Q5eEO0zS6xezNAZ2DiBmSUEqfe1Yy6
cGKd57Vn3wTXbc/bQ04GY+zXsyJNKYPMGcsDdsL8gIEEdAZdEE7Lvkf0HtbaqZ7A9H37IjaKVeB3
sbJsPjM9Dbr3U3LUTm8c2H2MyryBIo9Sdl8hM1E1TKOXf9Qe7dLV/qegSHm53VSQeUu4UUnV18JA
Lbf0tzJ9LDZisAsBl7tT1NXP4HMQPx2W2k5/8E5Vg9yoT1BmiROotbMiTzYjlYfk113HzksVuApu
IB+jan7ElO3TYvtxT6PMgZ1Bk+QJUhQLEg7ZkyKCkd8Rv5hyTUCDm0pC2VlkhFpVEMsQ6hev2wbm
cKBe6ishrndD9t8nKs8q2vqNK8w9OHIvv/7YW4TFWVmWnASOnO2phVIZJth23I5b8llAD5CG6zhD
nf3jL+YAOF8VAu3C4QTk/61q9SCuLVfm5VrZ7nC0zhSsFhsztxoe/NV1si2Yc6eHJVOtXVwm+cP0
IIQK43d5llxoQZTl93uM1mnYHbHVzrZN+ZthQNjGXwDV6rnmH4tI2zKyWOkgn5vpL2yBW10ZTYvs
t/ZXKkjbxpZeRLXtlDO8EPo/VTN4XbNmIu2QTEr/A/Mpfom0MNqzMJNFVuMoyXdZNYKsNK4iWkOe
1TIXwFxaGDVUN17hoRilVW2JZcaLEEuRE/hKvff4rU/3r7A6yFWCKTGG/1J1GoFlZVN7MEcc8FWD
r+oMOQpTo6JV0oNHQk+PMtXsnJz3yVF4EOCkPFD1/COyDNDY7okPQJVQu3eRJz6Sr/hx87pqwVlf
9J/ol5eytgYPJVXLgWZe7VkTnrmkTBh41/qRr5AUmXz6qUCkyNWrWsI4ARU2wiuO9Q0PZwyczsfi
j4qN5lzTKLm3cuexRXEwhAhui+CdOKeG4s+1ooDFhHhLqGfLYGBzU+S0Kyu1wkMu03k3HV6S2ABO
QyeOuj8CRrzOcnyUyguPZF83HkOq4xCa32dwoEbW+orlGLeupxwZmupfZZ6BcYFSFsYvvdQNf1xk
NuGEquQymiI2U+ZzHqWyMDguIuh1oB6/hOKWO5giA3pq7LTZHveowNxaliDDY3YLn8N1Av5fGg+T
Iy9YzIRmhrzZyYKJUceJD5CSAj2LprZnAZt3UWh0Rcx4vMpI8iTAAWb0DBrS6rf/HHuGBWewsk0S
LFh/hjuXOzoh2macIpVgWfeGQVP5ZKiNAkTBUtnUHaeI8h2jdCEIoNeqhpzFHXOf5cE9zI8wALiB
ldUAoth2fKVOANLBnuMGeATqprM37rX0eW6FQ1dlOtJhA0kDMMJXbndk1DQb3fl2a8tghtohWqz6
XZslBRDTPG1cXeijeVM62LE3mDB+Xbgk9Wqc+RCnzMeU6F0fI1PtQmkP5AnEvijRmrSRv90ggbR9
7jatp+ojS+FXw7nO3EY8+HgdXEOoMrxO83VOj/s7Xv9qlpX5KugKPcIArwYgN94HCefZVbO9N1SO
Ka4BlXOPilV1PsmBWIvo7A4lP0HrTmlRzRVV2ngC3XgoxNU+64IhcvzR4/oNOkdJX7TIb6BlRRX6
tJAZrtf2rKYNc1rVXDUWl0tosEjr4VP2Qr2r+Uu1tDjEG7syN+uR2hQdLX/c7cbgiC4xEK4BKyDD
5o0FAos8S4XzGB25GmLmtEBtwICxJChpHrvTh5GGWhtAkPIDyfrC4Yxm0bd1sLAzPFjMuif6prbe
6l9Ba87rmnoLF0gYOoPbqjP1FO2GOC1xZ1uyl4yeI+TjOGCG1Ae8hq2LOO5qNWlYvVk8sV229wyJ
40xUBveCqO0xQBwWMKwicULfe2KxCXpPN/cQC8F9eTkbzP/358xUnQYvAZNOgNUEKd5Z4iIcZoKp
/zJ0qvJllYZIzch0lvgesLg3gTosvM93E42M/J8X1/I4OJFVGysO9Vc2eUban8laOO8NakRZBSYA
E9wOqLbw3njs3Y44FI3gCuFwYQVT2wiD/jQMfWWL6V2pQEe1dhoen+rfx6mKmHBv377/x3ltBcQV
pAGNXIGXuytXjQNIYaDtlsUCB7w2H3J/cxBJvYTb4ORSjk5aLNzrLxj6kdwOvQGLnEXAIG098ZZ4
7G3YkBpx1vPeB5zprpR9Dp1awUaxXI72Dd9vwx178n/7QZAPk3PahGKj1C2NeHbzX1B+0M94waim
oB1UyVaw5w/zyi7LVNdp1NsZ/yyd1eTDlnkaIwy+0JhL1bYLHQlfVK+mEJSpzWg+4D3/SEVtOFPI
yF1HtUECwXJtLssbrdjRpgpYM/0cGnlMnfpOPc+XeKNm3coqIuPskLD6a5VDB2Wnz1NLNOY0pHiU
PdegVYPO4KZpoAhL9XG7Jrz3w6jY8SWmH4BhZiCZP0qErDQSwqExgySY/2BOZqW4rJqRQku7u2K6
OxpDtgbgqgFJKzALsQSXm0OQr+cGye+T0GtOlxr54fsfyZcgbwUjsX0GuRhJIDoxMc3AxBmw6t99
mzisBgL6BWrmzT6AkugZG3WH8rWT81t9Aha0fjNFUSE6pKrxKTvr3tr2iCEqClyfZt6R4mj68jj8
TZvqM3scUxFkfXNAa5/XDpfS1zZnZDuz9TIBpHY/5SdabKV4WP+/T2nLScIkKGDHRvkV2LaKx/8k
josW4zKo1dOt0PKmESG47V0On3CA8lniTMfnzPCFyMiAb+Kf0bn3Kw2vycrPhhYCwyyXWZuEVMOm
fxm+kwBZSXmu7Nrd+mcyybkdKQSmJHGdb1TaQlrSPbOcOc+UiTM+PVE1BN5eZSxsVsHULtmhccQX
BlfgTXgWLA+tBmpP24bee6aw2c9kIeRIFmFcdwd11aD7mCfbasXnQWamoXoBG5AwxmiiYJ1/JgqE
Yxk2MVwUZQmIjLTdM6TeP21DGdzLLF8h4EtDVpn07DDArUgf2A6rkdKl5AqwpaFqVD32H18i6tey
xiPI2nPZUOQgFgFLgPIWa4xCpTwflPeliYendlr9ZNeRM/0YzBzBDNFMCm53Mik8kwx0H3qsadUj
EncVNtu/hMcKFlEbinK95STz8dGabxJsWnI4euXlfqI9mQ6sGBZwKAoNjh2TMl+E96NZZOAaebZ5
/p93u/tr4RTFs0EhWLRZ5nATBerJeRbO+5mXRqOLqTdrDXlAba+LR4aSMqaQpEwRmzDadok6lq1B
L64vE5Lg2+mWLTM3rkLwWsXKRbAYaA2m+MG5YKGQf4F6Nb6V+tntw+TnhClZuzBbotGYumdygc5H
RbTjrSAQpU143Ow2VBAOOYIomkF1nBLM1JlttPC7Z2JriLqgSu9LcySTGSOKdrNMZI/fFt9exyJn
PuL4EiuBJq0qx43O9Ry27rA2fcTu54YAZKPcws3f74oisDRJOwzbvVOy16c/ULIGfQDgrmV1im40
vak0MZLteQLG0wgqPFtrseozfy7KdU96BmXjUJJQSVBp4yxuiV3FtIpaPxudQxgc43E8YcfuUmHa
KgxzTWeV4IPVyQTXXq5fhZL5K8vhxR+W96NY5intLS6aSCtcE7g8KmEaAqJv2rXDa49JjNlKvP7l
8Vp1gkXuXe4BhOX/pWO+Q7QughdD5vK53nWfOtiguAmaNOiIUOaXPWdio4OjfiLpNDwkX3VDoIjT
5P0ADiKjWWcjIKWClWw3QS8WUzx2eFn8/8zRwr1UTikknrRAiJTu2D4uU1HYuzHU9QrmxRglJu5l
utAGHJUwA2qw2iz7xsaM87AMtPosUIAwcmJS4uTMZoYYRxrHf+BXC6NpHGdmNnCUUiO4TM277+yp
vJQF/p2avIMklKW/fo+u3zBdjwpvLH62yZgfVvmZFTnPaiXg5IjGt3078dATgPKJDevOdJKVavz/
jyFpG6/9w6byolnRPMGnki7mPojYHPomEkO1nY0LUaKjJfrQW8Nnq6mZp2KjbRII2SLyd5TH5bgT
OHYrXf+Om8452FyAMkFZ9tvuDA0cMDtC6VxtS1lKE+SPGODZSmUUS36WvYBNdArWI4UKQ+CwtdNp
lUMrKzT6cPXz3bul2miQNonluOsh62Wf9uZvwR7YqjOduJ6+OPOaHg/luCBvaOdIMtsOJm+QL4gO
zNrcYejO3oEgaVmGiyK3IAKAPkqYBGzml/yY0eLgmhOhi9fpkXQz5CRHtjKYpuovFic9/kBePL+4
oSyLiQuR93OZ6vC1JiMaJOYQWAoL/R3Y6Cj7D1C1HsU0eRNS6D9mTtqjO6c5XVCbATlCbXJmiH4y
PPcktI1X1pSgHPp9tXlfnpoty2gWUso/yvVO9Fqf4rfBUyjv1Le1pDQnPElp5AFQPDE0HyYlX/ON
fmQ9OHrD5WmaF150oc6U4SnZ2DgpdeyoBmOHQoR46/UVEtWrY9dofVA6LM2Jj6YodQ2bHJIMJ8HU
23U/rpDPdu6tSojsptdGZIyKSPYbxnpFwe0ejq0Frx5zJZKrGetrNA0siWB2e8E28lN1gPVQHwUb
O1ydhyeZ2r79dmznAhgZQbJ/IiMbd5cPxcyYA2T/oDLcMPKyXZCoQqGvgLZaYeI2YWYsM+Y10caG
IwKZ00KkMNj4TWdVsglDsPq1wczeU3kWE2mC3gVCla1/T45TrmEJzxc/DAERTJopO9jHhU4DfTS7
X3rj3JgCCuSJEt0kuzkqgLdLc2PY8Uy950HT9yqFyePbt0+E+fZ+c4Vn82Ayxr8tQMWjwnuSA6Yr
rvHFWJMes6IudXY/LNQF16XADJTHEz65wso6EiUapITN3to2YPHnipPz31Fvkk+vlNUHCxe6SY2M
irXRwPVrR+c+k+LWhtGTtdYfmzzYwGdXVsDXUoTsueVTDItd5uYZjhoPx2r+mmSdi1NnPyzm/ryv
2nFcU0W/HRh2ZkgMBdWhewVYRRY4e5Inl7+DpMozYVFr4ZLU6ZMnkNQSpRsWoggj9l3SSQvQLBLH
g7pRCmM9NX9DfTEnpdj/Xd6JKlvhaEY2XwiRV6cgLa7jZzM5LFUwnLeZCXA5YipC0/jex//72hph
1CDXweS1cWZacON8gJoOTXLoQUTUDZ5xf+6ud0YqlpexOKtgp0GWjHT0qRsXQGkYdXGT/GqDZKSt
dJhY9QiroREE4L9GO37pq1bBVvoiVUrKsMiSR8YyQABs+VqGpYtnyipSC9SsVvVTu5j4ihSEqnW7
iwXY4tUXngygb/PHNb3JP2XyWxvyBCBtUVrPNqgVrnQgU9RLtD2fTL9IuqgaP2H54yzr57nj89y1
oQ1wFUDkvBhZseyCKisR0S9tzWt1S0kPF9x4/5NY0mBnoM5RgLFFkkWUFRo+ndv4+LsQOF+K7aW/
iTEDLvUYINCiBt1p0sHD3SxljcLRjW5CPjW3RMshbbcHjlZWWkeItb2SOW7HzppHiImW5cakPLOY
ctTdrhnEHJna1o6Uet3czVgrC/uZRuWIkGCZ+cwI+ZPlWjIUHrNK8P+3NtuvFugSBSw3Tp5XPFC9
5kPq8a511npTov54cWjiwd477BOY94g3xgoMoHRnan36yoeita9zRjSkQLdDMx5xuBjT7fCs1Zpk
xkVw4KGLxz0A1hCj6MtYvx0vws1Lq2FwLIBmrSGkM37NhFsghWeSrFKXO0PWPiKSxnTfq0HkZlYl
GIDD43RCfr49X7IFtOCjJuyVelu5tyGe+aQA8vWdaG4IHyEV4S/WwjJ9YYO2rMvKL/yRvA0FFLy3
5hsRRbC0VboiiafCbvvy8n1k257nMzMpjE57JDxNDoOY/yKVyhHDb2DcW3yxevvfP0cGwvf+sy9v
yY04htr99+JMKI7/aBTn4JbUlRKcGzK/onaCUSn3B3ZcvYIj7+z41jvzuMtaN1z9PyLYfzpt9/RK
CQxmWuAY/aLRIVWt825cU9KzBKkrf5PfDmzJCE9oyKEh508P9aYgTk6cmM9AWv1ADq8PWCOGY+Js
Gy37DIs3en9lErCo8I4oMIFpgdEw4HzqyG92KwDQzRbVnjaqvAf+UCfiquPgbGXHkk7rB91DvGmU
EY5N3X2QgvpVmOWm5N/wrF5Uj40qY5anzUtyhSC3QGvaEv4wbkZU6oEMzzAkHAM9M3F1FO8Ilvq/
BCnpmoJozlZ7OYZWORKESYWZExxlJ2SrnAB3NsD0hRkKseUSE1Gii6ykmXdaoWU123IillhAq+xv
+xhfRAr4xwgLiovFFKp6PuV2GV3SKivDvLOHuBfvtxP3SUFl/RX+R/bUFfwcqB3uj6eiBR4S1pwL
i/UymQ/4Vz2znnI9V1rGNdRzfetLIB3YjPU36pRPXtzJS1dGl8qz2kDDqpGOfJQd4BBldemKL0tc
bn/ikXkTJx6DYJFa4uNgvCGKIq7szzVW6iBegCqqV6QWWAt0p54OlAuLAh8jF9ziFT2Z8SgeSJn6
NCtjtEiQfRtKzTV8bfDJ08K0qhMf1Vq8WyOuVq0KelIVVViMl2lEk5jIst8mtsLnK0kyxlGfAJWl
Pt5PYPGzo3vEhSZ2FjR//c1UySk3fjWmAd7gIadCAQKDwhugyHi0gwhJfILCNNM/eVHjogfeKHfR
pkVm38cGYOMYZQeKqI6YOde+7hq/c81wTEBosq8/LRGevnkKsyLsOwqmCpneYKJHyA7M5mYeK0Kr
tqQ8nD3xwdnxX1DRZIkpiqDGf6h/5z3ALU9YlOFmpBWu72GdFz/PWEOXLZxfFjfhOkz3ISFDe/Gq
A8T2B5ZXQJN2MJI2jm2TZRv9JLTQaUC4h3jN4eWkOuAS6BES41XoCQn1nutxnTnwUI1RzxFcDafK
1GUnvgKXMsUzrL3sW5Pp0J4Xod/KBDbn9Nxmc5N4DnIe31J1QuMq2RYGG6iovJ3llMYLOCv5Cvtw
msIxOiFSMjHXV4j3FoY5rAW0wKmAZe5dSx0oewJl67ALdTV4XRR3ev9zwyigSYlHtKP6Loq/PcLn
mv5Oa87h4+WinzYj/UoXyv/G1K3Udelpu4ysKB/Jyo2tT6T2TjtE9WO3yOP9ePN4jJZSo1YhHLsQ
xZpY9khrMk36B8I1s+xq0xoeIvKUIKh9ZFMhxX+ZzQDIDDNaGzGl3vGZnZ2WAfB3CQkfZFSkqrgs
hs5CALaPAULRefGN2rvtukzx3fSbCdzm8srT1AvrMj4zq1lD+uzozCwlUaEyS1UkIGEheR+M3EET
5YZAMHhgD+0NxNuYrP3ar6td6CPFzXaIaI7JVsd2ZiokKhse7Po5hUWGwwtPSEv6vK4Tnlo1Sfi4
O4N0V198N4n/QYMfep3x8RMH2XDZy3hEU1Sl5NN3dbi8OYuphpP+CYn+By0BtbF0KBjM2gI/DALB
98DUFda99QzMvRw47D6KNErTnC2f9+efDpgUU/0wYWG06r+BK7RpW+4V38DrW97+YHkA9/4Apacb
7Q2sU1lYa6NGk259nFomHE5nX3uGKZH+pH0aV2/iB/JOWyDOFoZbqeOlzrwwizjql3uFmntI+ErA
ts66A/yeGkAw1bUT/fNadCKVLhQNnMRI3vNxCzXLHTwQdy4Ko8OwyV3bb/WXiUeYszt9WMRa9M18
8kZAlRhHA9Rhh8R38v3lYAFRuTkWaXXEmAe7hU92esI3iw6GdeUupozRkSkNeLKDgNVUA+FRqdKw
TsYri1oDQ7FTtGf9ipRcpq8TnzL2pZWi0FYPYR57JP7ew0cv+BvQDIX0FneYbctwjenoHAEUMy32
rSlTAFq0DeAQoMukjcvLnjHKQDSrRLsEnWYfQNC9OGBzqY7Wvg7rzRcWi1PnxpAFnIodOIQoGBiU
rzJN63WJtqY+bCorEXnZSEb+jHtOlUE62Mz+BIBo3FIsp8PuhVxPU/fULJk4bVTIMNFyjeuytlLz
awFLZUH2DFlMob9WQXydYeMMu5/kBQxZEKVSWfHh7bOar5pjQKnsaE7wjolT8IjmO9hs278X502D
VVvBE/pXa3YNhSFCVfptYeonromQtuusRNTvBXGJ2B6Z0Q6Jv+ik9ikr/6/i+MJmeS+HIRDHEGf9
VA7Sj/36DuJzLIgfwayWqZrx3Nyze2fV2BaFkAmNiL1ysiH4hNin8beeTS04PND8dIGz+Tfc6nTN
d24/C16k3ZR36PoOsg7VzN1iYw9+HcINyGqg4cAWWITw1Cki1OLSx2SXADzPJvKFhw2m1x4Z0usn
6FMe3YdEFqTOONnqwgHgSC2MNrpKtwE8fp6i2sfyiUVnuPjGolBKmDSc18YzTUVowV2ifkaLfl9O
WnfbBtSYJhZ6LmETCTxLu0lEy8EmgRO0kOldDpQluXOX5Zl4oC50+HFNpM31jZZkB10HH/fEBj+q
bgvdmldlNWs+xJOYmUDSBZiwF1JTkNVbdjw+au6ttfT2Zyck9EB2QEZr5mNbmEZnS3asqhykVZMx
XITHSwhRs5C2v5wm0hMBudDfHP6kOfi9+ZKAi9+jwo8MZjFELZRGeMt5OP0VSOB3Vd9InYU8SvPw
SfDn/SgRiolREylbJTMRhBaRu1FBkFDKBArtFjEygkYc2J0ZX+5ME8++N3S7e2vke8Rz0kmFBKW9
ELn/o9CCgurX3hzesLBlYwnl7t/019LWsq4mvyZ/md/ilLUX2OwoKdiDGV+p7b2ClJpbC4aCKw7+
oZeLPFFkmkYqAZ5U/bftx0sUkZI2f06OLb+FIFIsUIge6SWFd5EOegSZt2llGDSOuUbnCiI80iWo
VzmKZYR8oC6FcxNESJYEdFL8a6CwDnAoM/xCN1gb3QExS0h/+QtMXuumuXonIs/Gdc3A7kx87dA1
yh4W2YDkTqeYfzag8+dRW/eK/Eh8Z3qLKjc5t2y/TdZHCYkdiCK0ikNHLkzKCQD+v542v4yEV9TF
Ndrn8sjJyFyO7SqgHxroKBhj966zp9nHxPgLRsuYeX+aocGJtDletZj8psA8zqYLDQVQZnlPcM6r
hxGOjD2X2fmtwey1DkgBbyzegWk9R7QpcFNYIBu8YtdIpg9efw5jGCZ+2XP2rHOBW6UxHyakyY8h
obm5aSiVwUcgaqT6kJXDPD74Ytzdr0AvCAOMxfghWDInEb4SlDE0Rlwr/quuXQ0rVp/AbAp6+KtO
it0LWrxdza+wpZCEgjnK6/OFF3T3PcnaatL5OR1cWA2Zbay3zjxoBt2iUoGAaufVEZoQ1/WQkv5Z
QLUyZp20Ud1oIhMIWToIP1uZrS1Z9oaXCPJf4E4q1VUY9ODkIyiZNpAFTVGRRLOPAsZDiG78XsCa
Zvr/EUFyb1dESqXeu1tuRZzO8xudLXDnIBCxnQVjHH+TCOTqtpBaNov1kD3tjpa57Y6yl4ccMGbz
oyuAa/ln3X1JFyV2DcoVL9DFgfRbIoO3ogHGueNXHwFtv47Try1PjgI/MJ2QGfRWYzixhPYw4upe
cVMDyN6fnurnPSa/7E5pLNmExf+nTLOxUUuE55dXLCT0YrhEyU8Q+jA0tmdvcaSzz5JKpzwX+lsC
r3H3D/LyyPS3rIUwuSpun1XCHKCcmHgq62bLunqT/d1WixsgGUPBpFC50LU6hQdytkTOxoSQmMCj
aePuEZf0tK24NIz+3C4Rr4IkECCRfEPSxHMPRDKlKzHQUvmRutIjtIq39nJbE3QlWru2gNtDlY1j
ANs9yn/a2GNtLTC8uGDen89WEzK8qqcC2ljw7fuPDAFgLZt8PDWEcxuj41dW+YfIZ5LZIFwAmeK3
vpiXzzg9A+zPLATuUDbKtaXgLHDJEzHwhwzCd5mHXw+fJNnJwjcZ6DGzvl+DZILaCI1Fcd1+Eq3L
7n9s1nWgWUWZqqBDJ/wO+SvgkhSQ0m++bnl/CLILym34W8y10yChv/Qelu5qoYkCIC5n/HYiE/uq
IVSOeCmyS82ZVt79XnkQQBloZgqViamIInjejGFcL8cf8SB56mUgn33PiwfWjzHwjZ4XhqF1a1+O
E+veZUSXL2hJCNWp2qso0bjHQRtocjX39eHOFQVEuRKl+pKj+Ft+7iRjp8IaMf6QnEBJ6j3I5LrH
PBwSFFnXD1BA3croKIjoFHxa1iyrvTAGTacNJIdqBbOoVQA1pNEkWGXhNTBRJqlumaSDiN06fk1Y
Ntzz3RRfeXarVsdWvwgwqEhu2ZP2GpLv4Pdm/02Mcn7LL0tlZ4iDu8U9U61u93/2cLsNZBaD+9ME
26iTDxISRCpkmA5OBM2scxf4ZyOxKd3LJ8MleyavzsjWXfZ1LZkj+YuiabXCmUsR/M0ZG90GA5/f
cKEU6+wH83+qvmzRme+VqLrAYAu2e+WZEAM54MOeCC6JUP7uuQ8l/a+t7YnwEkt2Vs3DDZPhxWIl
wdQ5dV3vVYPymdj4DKMLFY/OMlIvh5tkcXS5R0cW+UXKcZIvFSMA/WnbdFHmNnWDIUGZ1t4Ky9jj
9bkOXrTKunJNY5C9kj8vhZvg9s0RYfKaGDG8sh9CriKk6SizA7vxflbTfboMGNHw8IOee74TfwAR
maEcD+bHzBToEfWFU6conAlQ/Is7InrTVvwegSTthoffaA1zcZYASpYVh9hKH2i7NlDq7vpLjVGV
iObVLAEiAQK2cw/3qFcIYX+NmN5ijOKwJtLSTZkIDMPHcH46NmNvEZNzm72jYBSPg3z+C9B2TqL2
/4rRsBsTFRrwteu7U2kQ+GBubbF78KUC0SzV6pFdfnwafm/6uwh61zZuWGQfFT3emPShG+Nf7t4C
lJHwNJsFIg2VLAtYx7ZTmEHQebPN35RSxs58P1JDmurpe1s16xGJFg6ybjbOGEWHqyYRdbtk2dpj
z2J/q8z38VF00tB1pY9FxEi1RWoMLWO/9lM/JX8Ku0QrvMoSAkdWY/8Ypu8qVedftFgPkO7XfkzJ
gSG0M+t/vXkNoai/sZclQE6xUPRKjjdKPLcBssQ3KZ82bOABHpbbgT1YImGS4oQoeCxp6Y/uEtYc
1ZIv2/KA0INtXrTOXZna8I1N50lW3h6To7bbBtUhwaDg6R0enSt4Q/HkcsxsQisuYDzzO01VfM+z
nCk2LtRCx5XjqZHXoa3XRf2nc05uNkbKg2Wj4t3piMw9kbr1teADqMHQ5fukJFS5bz0rKKklnT7r
BRuvrUHbqLedpyILBw/A9tel0njr1moUs5QFs1ybFVOa0qgAiYfq47Jp9hRgfNp9dzBZKgn+hNQx
V71Vju2oTEbOzupQJHfTXL1+xzL+5soWYjH59EbZPY+lG3LR+u7LOyoZHxDPPOpif2o4Rp04dmKg
Lf0WjcNizY0GMpQPlqOzRPR9a1/3tArXmcEUs6zlrXW8ai4bshxs3JxcShRSJ/4y7Ys3F915SIpK
bZXGi+yT0UmlPkOkPm53TSB0M6BiHkqHLebpFkxLaBLHDn4kOQ2juw4npfOccX73oXPR65TXC4sf
rsZEdx//0VTvYH851pGdxFxkbco4IXXP/0VZ78dv8rUFBCszu/goiCPs9snbr4HEydmB9Ye+F17f
aI0b3z5uGk3/K65FOT/IuExlianxFjKYCFt+mdcuRRZv0gf9Dd0fq9oxiWI6zj7HdLm2/QYvISRr
TUafArB4Av0dceyk4hT18ci84SSvHIvJWGxMqjNshib1VWRfqtjjR5AlK50P60QdMhM0DiMBeIku
lZ6nDJPT+TkW+CUQw6+KODUr2f0iIzWIFDgQmpAfTBYHw0c8IRkR9ha1T2tPqckWmxJyiVFLifx8
J5shpeLNJGdCQ0QtH6Ui5CAn1apXC5CCpSvgqNzyPpcnIHoVSWgVpdQ/Pnw0f7pz/ZDBJkVxpHZp
1NkW8OPITQpS7BREu/JpC0VWuO8yyBUlUZYWxNJWMkgKA3V7fnRQ0aoSnenKZftdW7A/HMN6S5sH
DuCSlSvLHpwJqGuUXY9QVSshgGtF3Mh8k7sXxIOA3vCVneReb0ZX+pvRfifezYfi3+OiMBw/Ag7c
CZLUdZSGyaiqpvq8hDdzLPac2rTLwmQRjVqNtL4nMjeScsOXtVDh0H3UQU36qiw1lUYP7p5ro0u/
W2jjQ5ALFJz/vMWnhl8qqzilTdM28FQ/a2oQppPbAhjBXLD2yonrZZi0NV1W9i8X5VvLRr4goGil
71eaWBSc56l+QAvQUElP0AE5CBOIzqz146416YA1Lze3WvIe/YxxlYvMHfL9vTF1I8GtTHAZ/zsp
oCaw9J96gE3Keyv0yMr+NwIEXrXbglzcecpgozrkX/5uojzXr5MMbikQ5TU9o+SYpGKQrSJxfwyY
n0q44XqOSe9GUD5cwklOTxe3R7e8Q6wTCfT5jmwVT9w06Z58mTnh27cOu6RZJjlkJbTZRyOoDV5J
gdY83RwGp8qEXaOXIRC2G29VDFN5i4A/YPZf4UB+4KUXuJY0Mo9qFozMek9ve/qfFO7OWzzDd6Jk
GdA9SEnlt1yyrvMFcj/ePqoby1Co4avKLh6NfSH3j/Pq+CxQSKvPrVEemL0aDnhy1PZRqSyjygPI
/CysizGDEIpnoE1jdSAXBFlFqnjC79qc7Fo6YricIO8U/eaLlZvwXe80s/gObT2dstGPU6lh01qa
pLDImr1B47DUwfVQSF1qbhEvnBZmchUd7gc8AMNoMUjL2uFr4O9hQfvbBk9GCPwulvDBgcqpJ3Cq
WZq5uSYXPT8Tm2k250Fvlf09v20yXjBdN7CQHwTPYkUekobmqDUpUwryqedsVmBGnFWQXMofdAHH
g0rPHQAwWtdeUJt5tf1e/MVLipcTjjo3pRLFaHSDc4caNenN6d7/5RZPhxo2s3/Yneqi04wvCF5t
JcowOm2Qjn0fqY2vw4TY8uW/VSjrphp4cR/zkDoGzluNu/GSUMejtaYQfaHVKy0BTog51jiK3GvV
bOY1VwN1YIFktgzV4w+/qZDbU0EpSJTONn7buaw7Gm4gmiYsq15AbnBJkVEkRsbjrnMM0k098Zu9
HUmnUHUZaCVz8rzopMD5yDRLPtBYpCJ7A3IOzXUvDErpiTF3lOnBwd6QoSGAO7n3BU2EZ+RIlXEq
vJfz5PRH9mPW2cJTmXkbs0f4ssg+qbM6lLBRrynHzTZHNq3jlUL1VtvuxszRAwxeLbUyZZb7JNHw
BYucnEU3d9owAC+uoGrsA0D0XaVoJag0MHrR3aGUTppA8sxw/QA4vVtIDV9jWjgtHiVYwKSInhc1
hucdx6QCThXI3VQC2KGZKtawL1G9sLeMmd1g5h8tZxsASiAkVRc+3qWEFTQCO4UQ2ogHfdhLk5jz
6gnMnufCXW6isxdIN2olEo3oa/7YGbouw0Aor9uhCms1VUeQblKFrg44MCv1pRVSMzuRLmUke9wp
Daj7oe1+IhnosPJatdYjvvy9BFNscyBChnZAXCQOSvcPJrmaFGqW4tZzvOppU5XUCuDkL+mCfKmQ
QBUNgJ2FVvdJdPLqca866MCLyqOeTmekv4T37n0FSvZitsHIvhjKARRVEDa+QLehqmb1nt/HqQ0m
YzbMCZ3hBZLZ40ejd8jebV5XtHcG1lAyQK5WmGOFaQDXxNxV8UT+I2eaY4BAbGu2yuAMZY8DPX1c
YxeGmGXLQWP1ohvroM5TJ/mbzWUIBKnUoKUvfrasyQcrcw3B55YoPclVVDpjCv4GxT91D4n63BpO
nd9eDEmsmGEOWf7FzgovEZh9DK2T3B1KBjt+qG6cAkF5qmcmZoldpq7f0ODeURyxWYcRJjzslobD
je+lpcZEZJRA9j1mc+Dep/GH6i6kaZOqL3PkY1VyooBHiidCXZkivkiiRhVmFMNs0NH9aC2TN7IT
94GYsBaQquKE5GAWBJJk7rss9SBxad+R4mCVGFkXK8pWcNQlfGKtqjXbFcjHqWd7pY+wtgxZ+GVo
1mlHHRqs2FMvBcorPEKggqAtelgeDxnMwUfP4BWzRStZC4qh2szt8CPNxMrGs2iGi7m486WSUFue
hmvoJn7lW6y401EwzHsE0AChLUpg11loSI/VusOUTff2f8SRUiPmSZAv8ONUooIWEJqxoLFqFALE
4Lv2JIepo/zZrZKnJ/ajmUXoosmTBEN89dJB9l3wFK4hNU5ZQb+t7LulBUmdnsOoj7LDNfQLQdMG
fo/ozQALP+3HSBMnRytOrzi3aIGnuaSc0RX3l4p6c8UEEpDpc3IykTK4nlPV9JoNeCek97hfhUBh
ua/IIO1IgBn6/yBzCUi3do1j3GafEqfLhZVNtaBrIZBIT8zDlbR2/ZzBOhtOMnnqdiG6pMTJ9TOl
FbE8b2Hu7R8z3KwUcR9zjjYjDFNkBFr6LEcxthvPBZTaiUPWMwpph1MTq5rEx0K6geQvRbkpmCtv
R1VAzCvg+0BpSjlTBRCGnNcAVsjTxl2nyvG/2mdaFJdarIMB6kd/+K2ezv11uMOcyFvV78BvaPFm
7DMTBUf/wxuhgA2JB5tkw0HMfzLYfDNfwEY0h81JjGeWRIfznxiJNHCwLROwoyLk2Zy885Oy7uGe
ParPAnuOYH05rSycUxLtBrVQqXs19/OaSw3zsY9rEuF5MDp2SeabtvfNmK7YnEqGxgbt+blQdUR4
AgaVH+IgTjxeWgWs8jz+2R80giTFtm0enloWz2n7eQlRql0HqdJPgNc4y/zO7b+QaA6JyG37ltUs
M+2c6Q4LtYJm8E9CZSlNjjFA5F3lySk8F3FFJv96gQWAvVQCWHccGh+QW1OqNYGStbgEueC2efnP
vZJCV1SYnMlPimTSflVEjk4DAj9QkDojJqr/icViOYIUjHjuSTuN75Q8XrPWE6exJE4n8zYvtweB
8WbEb9R2LVVBrYUGGDWChDDquV45tipeXIDlpXGZa2CTgFhrUT0Oo0Ou0Kei5fXQXAUWsK852/fx
8IJh+M6Lv/pWo/L+9KIx3qjhYP/tPrHZ67AJsFWipcevZcjeKz2lf7KPqV9hRuqL5Df0hO2cC0XP
pzzoo2drN70ZZjbTC4Qpv89xfYSPs27m50yd0LUJf+kIvncWM+UUML2yULelL95sSK3gqzvYzQCu
MJ3CQudDsetdAcwQISElqct+/G9adpq9wuheiwfea5l54Sc9/uePfR/ZNIVJMdYEmtLj9kXkxsLG
sa1U5IfK5NrZEn6omnDM9cvqEqjMzzyAq5NOP9eQdrEQyjqbI6DUOQ7Pt+Vi3lryk6GTZOQW6l+O
RQsX9XSe/VVyXW9valSTBv7/PYn+zhC1il7x7v6FKJkYVhCbYJ4TTZiLGPpDPIzG7AqN3WAaDBU6
6/potwRcLojxmZ+UKbCYENdmdGwfbsKJ9mDb8jGV6FyAkRtBaqw2JLrwjOff9JzIH1aB28I/ijF4
5QI/U0ocgVf/YIdEz9X+Y3n20P7pfTgKyuL9T5dRLMZzK/ti1jXrhP67g4YxBKzbg/oJsZFkZilq
u0DTJ6kL9wHPsLae/ugDcbbWnFYYh0/TGfCCbhRLJl1EvOhwlf/Y2K10TGqBEoZTVV+pDZV/feFe
zzYdKd9HMfuhVrsCOzDeXRczWLpiCnLd6ErupED2++jiutDh5lVKRWYPNHZt423fS2AyYLGs+jfV
7d8lZsd4T+UI7FiojBRo7LC/WzklIXQLxs8GDbseKDETgbYSu0VWaAhrcO5ca/C6GDFipnMSWNfD
5mgXPTcqEykLRWKl1RnYyF2HlVe5r35EqnN2BBiQcXy7BIZgulwZc48+Jjgk82+picYio4EvQsDb
qcUFSrCf/IX6/wt8JIfcRZG7qDBbrqJQGT9rmkrJKOJcuAzpZfKWRR5xUUGVohj1Q7r2kvxEKIan
pfgJAS1Fm+GK0unA22IzSrhk10qLOLKNgladiViAHHhFc4sBrmZulGYsMOblUavGu69AYp3bIB0J
y97X1P6N6csWxwbz17oxbBMQpEsCA8EWC/zyIP51kbHtBG2Rg+b4PBKyTgVuLOWqlU5EhZiYCQOE
5oi05Qdt3ePID/NFSC/XFJ3X+fvZQuFvCwLctTNoZ5uMNpQ+W7q3ptUOzLlEemyCbV/UJfSsU8DI
prUKsNkTfirc8VPDpOEuKEO///SkNL5GCO7wCR/0En7OAUzPYPRoOfNBsMIPbnV2QeQkWC/pyhqN
Wa4ZrB0mcPyiUaep1Jr8Yl5p18WCLWoVi3QRZRNUmpRbCo0YKMsCkfFiNtD3HSq6ObHURLOgMHaz
pN+0uAp26F/dDuN3mHubRm8z7WvMrUFRPHASnH8ihZLHB+Ilz2gsGc6DqgBGO2GRnNQpW6nuo1hy
dLL29YadKjfH38NXvXv80Lwt3LG0rXXPsah0BRrH8yHLevCzEjEx8F9ATT6iNufiBHxTEVL4vhPh
AlkuKyX1MF3XbLrgZ1KylhzwLe7Y9+x8K7T62xw6ktiFl3Rf0kaZn80o1zXo9Pr+qtqCme7DExkg
9dgXfo4BKYf069PZ3+3GHa9m2qzjloI4WfIURxJiTF9E0GY6f67xVwTczwr4wWuOGecMP/2lYMtH
ueVMhAr9BVhnstUqK7hCbIzQDPWYpFnQpZ7kAQZwBHBKMcRaJz63+bNHBrwD8T7xdCME+2N4gOoQ
FuRHKANbAijccSIEN+rKNvDBYkcoxjW28s8Mme6GsmkNOL17/KxTCKcsIldqM6topof0YcNOAhhV
RTEihoPSXp/cQ/oJ+ODlfcXYlOYEY7ajnP6Anc8sf+UUXwC5el6Xer4ucI3RBEp3c6GFn3DNFCGR
40YSuJUNO1owoz+IcI3OEtNRTj8LQkjDnjohwOMvC25MxzXv+fCdeIX3XOj62VAwTMqWN4TqfnSP
vobT7Ax3dm3R81ZuPYMNZgDzv7n8DAeNQ6r5FRIUQ0Qdmr9KPJptWxuZvQaeQpROIhWXGbJnLy4k
OpWRpJP0Sbb45AjW5gehS8iJRe8nwHrsdnePLp+IhFl8838T05leeOUe92Y+gA9uJc0yfKuIUxIz
fCtLCvq7jx0n0drLIFEnT0A/dZbNoSmiKE8EyU23z1C4+isfEylao8v9sLulw/eD/tphkPPKcAsN
btvKz2McJebWTswQ/XZVg9YahbdWpgn6GT3B7zHwzlXAhMmNhg/HNGopY4me2Pp8Q6Rgqy9x3dZb
NJtva2uRej0fz1skRkHPw4BgZQ9a6+X9KcwNWCV5/RSo3+b8fS+S6I3zF7FrymwPKODi039/xPAN
2geA6Ka0yjOvdSL3FkI/hnIx95sszTNsKVEDFQy9Zzve1X1h+LEyNm86SxJxs6sedadYSVHCFW4k
ql2iOvrlIWQO0ybEavsqHt3DyBdkGBrtunDeZPA6F/utA1gn9831/mI53HczlSywcZ2Upkj4yY4I
Fg4cbeZM0LUO4geuTfzQctRW5xkZ3nc04zSuAEk1z6l/AueWnkSKE46zV9nbyqzpxP+HX8KbAGIr
ZJQMJg7b3zsqZnjZlmfdzAsMhtvayp3lHJgvKAW7TXqKlSvtXxQHhjfNw1js9YmQoh/xPdgiTgXf
Llhwlk6Eyaz+cKn7jy3W/Z0WK+7Yd5E1YGlTzDiQOswsz1SvRTUiURfF4zxPVVHAPHvlO+CQkcj8
76u/hA0tdWbZ1koHumOzH8i+e4Hel2gDRdqd2gteJIxQvNoI0sgPHOMFARFl3ROHCnbuDrepSNFe
FTqFpeet1EPEgKVBXks367WibiJXpTvczAwzvtgksd0gxQTCKX5P7s8ae0Xci5oLjr0NZhu0LW9I
kw6XQVf7f2WUQ8IPh4Z0DXe9IwAdWI4sr91BPfD62MlT/xRiFk22uCUTKlWqn5CLv3A6OVeJ8kOU
dno9BXClUko+O585mrqJvLZ4bmYxvpSh8Mjinq+bMp9PeWryykmD/ev5oVrB/1z8ewLDcM9zpIPL
9n+d+93aR1IuWNB1C6EGXG3rt6UCBJqjS6l2rctOG3bAeHrA9xRjAf4vMWYOMCfleGcjU2TkKSVT
Rk4uwbYLCQvQD+6ASOwHX8g5wYqWIcsNCa7ngWMtHmT7VPUYcT2LLF0coc64WHCS6WrLZS2cM9Ae
By7a0uSZRUBBRt7v7OETQ14mtd8i5CQFKtILDCszLzafgl17JSPuZnb6ahLCW9rcLcZr+lme+cgI
Lf0FT+j8Vg9eQC++R/RaQPUH6MIXANEqmOpM28WjwfAskp9XW9Ujf0nLlGryqLStiSA8Ft7909nC
FUlcKlLvmCsPbsLTYltUgoedPJ8YSeLCY4ejpPAeQ7zU6HXmljalbbxIYjpZC3FoAqZLLRNf+899
fKSZbPjm77472/S+Jk180PlYuZN9BCZSBkzk1VA7uUeu5p6b6zIPFmM/pMNxRDvx8gK73LKABQ/8
WfkZKvH0fJtBPq0xnkyE4LAGp1Fdx90+c/m38ddIBTHWSSNf0V0xAN0dqJBAKKoD5qUV+sytmf9b
iFo475827tROsow4yCGv+W+DLrRlw4DoMx4zwnvhmwcw0rZ0ZBp6wYsNv5gN5+RWCWgefHMBBVuX
9ArAfbD8Z1sIgUzrdQgjH1CKzF8NeLWel/edKVM5seHo+MneTKgtpoV2ZxDaUJImRN/GVZaENZXi
0shIYNkROveSOy09gmaYUzs+FS0lpwOM2ODDXhUHc2pm+jBdUDCV+5CKgo3jxzTgg0oKz2bplT2c
BtyAvrytnKCMHvlp5lguSleCI2bNmRvttaSrtq69swWkF5u1WM7DLszQepeVaPgEDGBiOZwMFTb9
JHf/dT5pHzvdoLMt05u0XF//y9msFWqSrE8e+Wsa7gpXhmdwTyLcjYtcYty4MigQNE2zegNHXbLz
VbWJpYbgn8DWO3nNhzXDqRs2KPwF6+M4b+eBcs/b3SjFlFvGasI5OXL0ACRUM3StdQ5V6PFb0ISS
4kXp3pm4PPLCQrpE0cLfaHmqhG8FJ5DWyPajuHM9eOSQyymCRc6dZxW/INBXeoDUOz2THEU9rWJL
FcDBCrOIdo6Xyn4TfAwdsK4Il/YCY3bJi67SR8ipD09IqVe13UwpDBJlUpaJUHkveUCJuQgLfr4c
tzmcb8BcDHM1lIV6fqmz9lE7G/3s8WfyYBE9Mpb1/YeS1hR8jDaPRrPJAzMTOhDt4lskbbwwtrQM
TLsAzeM/hfpnoCN/ZblZQihjWxh9MMHlqn0aoHhj7P0VMdferF9bdnw7TV0SPrTQuL/LoK3LHyfW
FNlvVULGCyGCbEW0bngjSpzPjEI800WCUzXd2VgKEtuDUL5OSNbili1c99c2+rMk4Rokc9E4WnHP
0I+Wq54xw7pDQ8lTlldH2gaXyZuGHutPoR6wh0jcLC7De2CHY92uJEXN9RGi8p40LvvJYQwVZGMk
gi7j9Lq+flSOS60EiUmt/KXFi/y3esA7+qiaXePYgCxNarcT7STd3YHNq7tzn069Rz0v6qoDcN3n
sKTWjU1SNoCck9jUmI3r7zKQOAWPjRHlsC/whZEwJMBUkNhoa2RcBYDjpyvlozvAdTYwoHAILUzx
cMYLk4d1v3TlgqcdgOkq1MOHAZHsf5jsJsk7CiiAaGt+9HZGu0alQU/F339NetTSswWctbcQR7qZ
8kjQ19jc0tpYdjzYN3hcTbjwKWNMr6R4CMw/agVhsm7DQBXsF7BjG01NXZLoFmoIF4MmKT0qsHHl
h9fWB9IDJahtEA/cLywFiU78pTVQctMubTw6xh/O5ZYLRkTTiQpMZJJwUPT2BWdAyWBS6xqJqW5F
yl6QI3vym+jy2+BoHhMLu0lhqDZFIx5gH0ZtAxaFqj4Vg2mN8PUg60F+svcAdA5PO7oMjGEaSjGl
VKQ6bMJ+Sh10mQVCXN1TSjAmYT0Ird6BilBXutc26xweEZRoLTjMmzNA6nkaXa9vIN1JRt5O9Ma2
dZn9DMmkaZhK4CSQtBIvgtFrPxfn5I8FAwxYJIm63be8dhuDuXSkf3S5LULFh6gdoZyoiAiSoyz1
Q4nENjN/+zfzvg1ebgNZIbB0sOExiOZqOFRiWj1B+l5tP48EcKHLfRzR4BWeXZvERZpQ7tdKk2ED
cYZYuemqTIkKc8efayXnkI22i4Fj1ce8Iy7TKXK9zQkk8pQqxeXw6NCV3BBsyObJYr5zX84c8c6Y
MKMtRs2Sa+fImvwWAC9JAvCzrhS7Jf7JQY7PrSflsIjGPxgaOiXsUi6WEML7yHe9vZ1nhsC6/5pk
lwrxLIranhVGD7+WYpkZt6d+SsId/ykWh9rHJwJi6hOrdjU776bebZn+/Jq55/ybjpaWYD9BDqce
XR47Fv0sInWKpPp0O4KcVk3Z1Ko+ZhVipxU6+St+0sKzSCvtZ09yX8aB+uIiH5wPQ2/SiJ2+9cda
N6agA8IEE40B7yKw9iwRyowAvGep9c4tVn4597UmupOUc8ykLdMuH0VrmrGMYx2lFUXnuWPkAU4S
pBKNvxkVV4PFuGgaA0FB3FrVKFfWE10y3KDl1aFVzBLN9Q2sErgcs5zdRPwFqlEIsFYhKlaXCES2
2hsEBhWl7Qwcqbl72QFc1AoBQWtI9vBpU4jsU/x0CeFsPjN9vGMwQ3w3weLylnat5LMLR6HnS1MA
jbO4aQ03VqSwlEfy+nne0oLo3q65cwTYOnCi9aF1MUeSNghrYThPLc0cl7DF3MS/EEGLdu16vJYW
Ry9lTnDxzTUloGX9/2crIYlvdI5He4ywvULW3u8Sm/mzv3Nwk0QiUNve0ixHU/Mkfp3pxVK635+0
NT1/LvSe74RZ/JXlrKOBl40la7KMEGBzcBkum28dZSQ+Vh4nZegTG7uRnW3H3ghBueI5lGZxqHZj
9MSGkRv3Cp8YNlgnur33FsDN0DrUmwKMn1HZM8+va8BYFeCqAtMROI4YCgceEgm3S0pmrBJ90OsS
uLbJlgzTLcHFYwTCTlAPldWWqF73uhfjriAtvMN9DklcKqjrJ1v4AJiEk4kUwZvSWrPqF0u34TVi
ZU7RpsNR1AVpaJmTCyn5fQVbtmpBT8+4F3wyu5U3oQnUw2naQlv1+qIm3fa6gTVKsNnUwE2ZeRsO
Iq7A4HHeIP7aXJ9gGBw9zFS3eewrSmpl9gg9EMl0b3h/tNmvOYzr3LZmpgnkcjC+Bzp3IEufCHzA
P60e4aFGjscPZ2E7I6+DAggium4DGYKJi23N06EqcrisSfyMvYrvwblPUvmdir6QYx0Z2zeTFfJJ
lfmfBfKck+CDG5y0Xcv3tkJJzsskWCD2SH3dOaHd2u7BXzw5vk9txYjGV0AGXYESXPIJ9IKwGgH7
SenOaitJiCnWdUSTsikgyvEAdsW6YmRsvLDemjERo4xVI2C1AVviKPdfZWeFLw8yIL/z13ILVYXx
lYwzvvvYq87ZcH6DgjvZP5mp8/2KScZE8pyuvnLIJYJktMapJ+hX9xGzrySkNRJ89Rk20ZqDYgXl
NhP9g2duaFsmSZvAYNK1tmCvKsJRskCmDZfe/OF0pMV38u2RU5riPcMK2mTIFJU+SwNrfaXaB7y5
/t2gwytTfi0trOHRbDx0QHM0Tedj/pxrMGc9/S/77UTpJZRoCAcGjD1YPDQDUl5Xi/rsz1tHLKDD
LeqRiurMIcFm6cKVSKI6I1GKU/jNV8A9l+tNPVMIoiS8gZFP6Zpzgu8W04ajE8occAWCRszXAes8
Y0VZkoUQM5PEZEr+X/Afs6ymb+LZo57qO5UfvSvbRZKwA6JRcM8vfdiVbEuJ7RgOuSAU+NQzEwWM
GJfQ1hW2UG9J3aYOYuzQBHlkf8h0pKmmyl5R+tZaTWGOAM9Gp0aGmCdF9MgSvUrZEPKyqeqQw9S1
wfbnrdlrUsKgrcOqQRyj3JUZ57Ys9uAt0Ri01r/ADfYBu6AjvgY6oYAaDocVSDeqh+uIOdCWlA5m
Mmv2p45R2l9BXyskmMBCw7C08j4+vgOHiAh/emlwt4a5WvS3klKBiB34WEQe8s2ckbQjnz2UWHCg
CkXIhtRsllh/F0cu0DQUTA8KJ8kqr6OFRP8TX6L4URNI3Qln4WWG5mX+y9i/znFB9vxkVi8l41B4
wjJnSdIMrNSnFks9MteHv3m9IieiMbZ1ewdP9lLGcbZOUoZYuaXI+Yrf3Kt6pDwN6/PRzeGYnBMR
0QRE8fSS9uxmWjOoSG/z9vdHM0U+gflQJk3km+g0IKDiKx5rJei+9ieXKhMxw1rDf+V41tKYVWiE
c5wmxVTKqoI9XaTBJlKoB2Mu0Y+WqoKDLrhlStSpA+ggke5eKNzSqC3EXkNr+FoEapMn4UAhTFrB
v18EC3LcMRNMe+bVjbS8e1RMUijE8yrj6r4ARaZbs+35ks61aG3wQsIJZcNW7i6TmKR2EiQLnxiw
n5B+g+hicgiIPSJtvTa3g5b4G98nunom2vD/u9xVAMKOyho40BM+e0D8QL6n39VpfCABA/v+ynTg
UWl+hRYC2NQEFAX1WJpQmiQM6OY1JC9NdjFPCTBAj/3hN2jUchReoLs+8bfyjDEzKOx5kaVZObrZ
fqy6czYsCy5lVMJ/gpl8qEGEKLhCLSKC3OZWMzEO37babRxPwqrtRSm0PRrOrsznwyUjlk55ulOH
yeRIGFTLkUVagateA9UI1Xks8E4hpLvF3ULgVQv8xkrckL4JiIi02R4+XfhhqKCS4erKrrXGa2rU
GlsP3NVcaEcIhI4sIvvLUzUS7bD8w5/pyRmpovJ5xxbbnd8HSpmiXY01ejJrIch/REQpZ4rbIbB+
5mUxHhiqOkTSjTF6P3o/iHFKdZxY2mj2bvY0g2relBZR/24WdTLtqB8pnB4bJEL30p7s0Njj2jfM
UnSR07BqVvP9bw5SDWTf6snb3884pGQVynmuSLPEivTvGbk7j+wvSp36AShTyq5kxKI41+7LyDZZ
1ErjjkcHKPesm/nuO6tH+Wx53CT4O3AzO4+4y29OgswkO460hTG9DBZKO7nGV/LjHT8GY7B0q+4Z
8x/DDqjFmp0znFGj7ccObjbRdkmNXM+rMNv9nyyAlDntoOfuRTZ3w8C5xk0dEoJ9o9GMIPEF1D2j
UsxpqK1a7/UDLihMXMriqSszjhJ/jw9qGukKtIHjPeKtu8TbkSIKiVVd0JVdv4SzEcGxSi6Xepb+
yhYCRB0PrnbgXPBoZFiKQbqIsAG5iQyA9GhP8bff6wKMeyAL5RO4yluwWpePsn9XpKRONgtqgALO
ZE0jTwWcE+GfYK197k1OAik5FYGAnPwutsCzU/dwTVypT9u1ku2nokpyKuCePNBRC9iJqfVaBF/b
OqQbbPo7Paorjb4PBjBs8ZM0/cAKaTz1rHWQrNLqL9m1hw7nMjjuBGMEMoIyucpw3aLjHUXk43AK
1TebWSAHuZUK82lN7SEJqZV8kvV1muiknoriJhK/1yH5r3T57O7tSFyZbbcEMkHVw1ya39GSpk5S
30K8OtAcaWo6MMQyt7FAuhPoeuPEZw8lieglcJuh3psU2iISsoFK5O6HBqRkIz9Gtt0nmxNGfFhB
LwPJeoVh2DR7gpw/IgIkDHEQIpOVD0JzglqDCsMQDaFxO+jDE49n4z/7HzWyxy98nrBETj0+USic
PuyX8O4JFc8q9Tq9PL2lfVhGL/awLoDKB+TCi7yrwRX/xdMASCWlGsdEaOKp93xA4CZBHCt29982
pxmPKDgm25TJRMIOLX3Knvc5X++QGynlzkGS1bxfIKK1w7w+3D4LTFQXBwUiKpHWD4n3DhS5yJ8U
sP29xPCL+ykENz+16Gu7h/CjZvGmnxPM/pI3U1zQ0Z+Bq+T4lhw9JagK+xfV5WBasWHJb/oRxLay
0LYWHRuOoAkLFmdFYLpvuYI4JSFpTjpU3o7tiuWYWR5jPIFEsTBbxjUPMIyG3c8Ad482rrmSMOqk
afYg/3lsYZ27M5JfJg2H2skmBeFDVSNVhCMl7DmKeWlagw6+H5aePthD1/pVyDwCJxt6QS+5H7fs
x1umwP57Dl8k/lBFg9910bwnSrpaHnUjGLnkMdgF8otobN5/vsg49lFHYZFxZWp2+bzfXMzF44k1
88j1JerbW40iJ2iSkQYd/NO+XC24fWE2ixmkPktLmqfht2+7KZiCko6moQyFXMFgM/iBNGyUoi+l
HqHI1uXMeK4yQ7uq76QyJCVhSV1A2ORNlPVw8p2COMgxXAPerxzGDbS77TJKIVOBYd2H4a48rDts
00HACFiaYoCyM9BsSPr0TGN3AulLf6JP/CpFU4ukt+8MlHOHMZqVKScuia+dm9iwtxHINtb30PFr
79gQX81y2Do5kY+O8TQhd/jAaxH13pq8b098C1wwPAK0lQn9byPyJfbWE0gVIbsTF01TRP3R3DBf
+drxTPLgNkQsjzCRrteN0Mewz/2DajdAQerUOhAo6Po2ZIM6CUVWF82huf4jArYAgXBRarSYszYN
5nObNLw8RA1WzdKhu+5n0FSD6qShWyje5XQJ/PK4fQwqZHXaQZRjj8JclbXOyhXsoJqmR2was93q
jbzdxtHrwW/TNlwlY64OjaJYcwHnBbwHgytwsmtGHjKWnaM3RRUAkiDJ38KwLOcpSXsu81V+/3p9
/VQR9NYnadnlMiYdl5QcotscL+4Ml/1bG23uJ2kUNKogOxukTlaH6oYpH7p+v2lM6GjqUmb25CRL
83BJ7iRjKoRsjC/5lx/kGVVSpU4N8X62QHEhPgN3skXz2ouAKuuCYz4VRgH4hvTUbMVsQbaBIooO
iKZqFHPMvoErXfVRkj3YUTVVh8QxOq1r3dr53e5FOJg6ggqLuQbzwz2Jed/vWxI+CPwciMUvYaZs
ATjvTQumzYHAAqOXzIPpAqYKma81c2oMZKCiNepm1+ZwgDStowYjaPtEY4L8xV0PX1Pl5XoZKPt2
fN3dZP1+ygiVYoMeHjYrRE1Y9ltKOPYnrZVdpiPVahX9GTlELzauaS+1QZrjoYotKAgYvp6ZrS/7
eqBKBbGv2laTWpz7TN6iDiVCl5XJr4b1pTNmeB4LMGOvJQZ4jbBjyg9OLRer7ATJ6No7dTx3bL+y
1jjZV0vXf7h6n6m8Lu5sI2TLqDiIeOq4kR7tDASCY7VdJdsXJRfOA3rI1/G4mgZA+sXm0Vl/c4Os
G7AtngpufrDqdmqorREpGhLJkz1Z81WTpr7Y3H0mw8zt5vAVmNX1uKlrZHxXyw++Ge1yS74lhORW
S/bQgqbrWB65HVobz8ouUEXlPEk5mSB7ybJF2e4x9RHjcXa4+GIA66O/r3RiWkQwKVPLPVs0H3Vd
3pmzdxB4zKwojbkMbXU3vXUTCeGojp7o90TM9f2F/b2w6ppJ76L+HLAx8j39QZ6DZ7qS6HJ0cjri
+NTAdbniBVi5rzPF3QnsSaOdG15Hf4mmeEw3K8/wR8F0Oo3Nwsv33pbFF3Vu3PyKB1xhuagNyCjI
ZJB1Jr7G8ltyLSjKQSC5+0MUa0qUNaOC+M6VJHTlm+S/iCy/epn95FdHOooE3aY1uZ9qngAZFswy
hz4g2xjcCXH80QUKxb4AOQ16HAR02JKfbTL9POo0SZODFnK7CMpsliG4RK3Tkza1bWV2UTG4p/C6
DF3kLIbgmmshZ1Nh7FOxwIFmZrwUV5ng/dg07tDXJDl4kYJEQQSSDZ9ojezc4r32RIhOc+QeWaw9
NyRdcg8RvKo911dgTknmAT+uvWrk64nPqFAofbOdiqqdMW0JLJnbPdSJkUgTxXvBiK0FCzAUJmRW
0AawBG/uRvuVfErpZA8PPjnFcOzKCt6KHWj1llOOBPoyTPWXwEe0vhDTrYshbTsF13nIMXcJJEr3
T6BarTWJ2t024aJzX5TRIkidx4DoNOODY6UkfyoKpL3mM5FiJciGIgYOvjlKlO9yC4W/6mpH8uHt
1Px94a0l3VKQ9ftEUPbSLxvamzbC+YM7QJtPLCTyo3l4WS8MwDUQ+ZzB2g5nhP2Bd/7uA/chlfli
PcjPQ7UYq4jGY+0jsEHdR0h/yZwnzd37Y9Aj/oBeKMLG8pb9iCzuXzNr4JHSoz2Qcp4eFKeOFVSj
X+bmqkfD8ZpXWnUMfFgqnVqlDuKV/W6xsmukBZD8ID/4fsBj3oObaMcriqSpGHNRq8kYIIPQjORi
U5Nu/9P5wR+M/vt9EKOjtECxZXoFj/msI5AWgxDuaEE8uhtFc55H1ekKt7yGm/MXZxlIjJKvQtzI
qmoXC5nB1lZZyA4J2VOxfd15dga/vyY4Lpe73uqjLOgcclcmHUUuWV7T8OTGUb47V8P5Kjc9mZLd
wPa5xNlmTRKnEmsoSZDQSyBEdFQOOL+3poTulxttGhIHuWpaJ4j66EKdYMTIpeIqNX0IQ54vWsV+
72al3MYgq7Z+mx7kUkrVch2asyCwfsi8KGmTuS7a2Frq8UU5kB+rx//XS1h/VvDFUsNxV44VrrjD
Y18+WW7sMCht79niUtm/GY63HVz8AtswALqvam6MGp3GpycoL7yWCqOh4ZGaMb9yIQmHQaG2DKdO
4taHradWzzotW4h1v2CGWZE1tsbI5+SG4PwrmvJGgLK07nDrAhlNnK5arsLsAnroy2RTHB7iimq1
+NJL8Ddudd4f1MP8UYN9J45EWsmxo0xtrbqMDpX/iDxvc81eLs5gcdVpiT09Ytnxn31SL8IIK2ry
hsbokyDX0XlKKBwtO/yjlHB5ddQvUj0EyUpvc7cCNCkj4jVcjYwu5zWBR2nL/QzgCA7sRxl+bi2D
R2arGXlvmTYK8O2RD2VlOEf4GZ3SjGQjde5/TGZAD/pzOkJXpHPqrWtkHH/kbOVtE8Jy4Nhfe2Pa
zRaceQbiXoPn86LPTroFnb9jBnHidYn2g8D12Z4gw581LyNfYwnf0nL9+aaRMGu4i/fdLLoKlsvu
jc+C/rQX/SiOPRy4Cab0y1gSztMsBtujaUqLaorDMl+Cdm9xQDHOn2gvC+vKsxPEdZMt6OFGKgwc
OF/CPNNppelTzXwvXs0PjZ7o64JiT6z+bmh/lyzlSu7WXYMRY0x8KwDjCT8v5oF9UARUGRAsKj9v
y5gwxQb0RnjOznDddzu6FvNguMW1UkTWbXHOCP7NpQTMVKjBDI3SD91pf2foxSyB34JL/V2oS5Qu
0Hbuu0wvccdo09iyVtryod+HeuBmAnfkKO91WQxHTUb+O6mYUEwt+i0o6h9S11pEqL44y5FsuEwR
l8W91UFcBl1pKeQeeOKOKoO5CcI+DoGWqi7gkZYs2eKfasqosh6yaUXJUTDSVFcKjoys+9oGpYYy
FkuSNsfJpHd1Z5N7fWblXz9MPnguduG27AlpZTVHl+dnofu7tvkgnLPpG7XG6PcE5LBCeDGDA8U8
khP4//JabnMIKvYJVGu8j8lsgPWE6GoHt1SdSwqhZILGBdh5Ozqdy2I083tcFl/B3rfBNaI9i5qb
SuGwrhCcKQwq2Ue25rpYjrqsBH1UobLABljR/6hfBXS5EYb/6vsWbzfDgqwbGoR3zHDrFXurtywo
PeI4zkFPCcOVAyjgpjuzUYI8TNOYSqVab70+Ckby2OD7P+T/5OKdQISvr7akIBH2D2KmhqcdmGws
ieUvjCrGmlljZNHZ6XVxtVtg6LZ53hYPgsc+GiJiz6aiR1UbB2RkExJYPUeaMN/altOVlxddOfBy
YfXIzveaNHC33KZjDLJ8zrbEDkjrsA/q0yXiT5W6SEFqNNbz51TonjHJA6ZFQtDtgdLP4KOcsdB0
ftc56oAWalYI5jaEfenxsw8xTPCEHwM6v/kWDRpf/O1UyO+9i82chQNig1DUowwX/R6Ke6FzeHim
dbXB8IXrNqXzCBOdsM+yJeUqueMgE3XkQ8hAeyO30sqaNcNFnq5rI46VJqnWiAbE3UqmMR1o0NWa
PR5jj4rvUTZUz+d7LwBbFfR+pLQBF9PDyBy7HYObAWrjcwYqYNfLKiUgBSaTC+OCMFyCNDN3AKCQ
+mFz9oMO2Dk/a0WbB8vr9u7IKxBvBQaJdKds1bO8GR5cGL+zhwjFZ7XxYE+9287HUGStlwy7s+Ko
vhZ7+EDEQHCN6f5sjvlHdDZ112WAGhx+IMQFXLf5CBV3kvjN+PAgIZ7iovotLqPzLQy7LBbD7bY4
1aiOrGClLwhfvnfKBkINtFTgNocHMdEarbquzKJzTnBuO2XXpT/318ixYWWz/Wo7GxrGLZNCcjwx
LQpFAu+LvpVb6YUFAhOiMUFqyH1ZG+2mgdv0tWckgNgr0Scr/qBhN5Ajxli0banoKgvrink9PsNE
Mhu9j4Uph76NtiReAoYQCaI4RvIH8gjxzfQSvP0TasVHRGsvKsZBSyzHmz1r2qf9iIIn9tavBQw5
0Og8izIbDo3BCcwcLg5zAhYFv3H1nzm+d50Aj43JgHB4EgSSeU9vB68Q9dbQNLiyltCZiB1kFIY3
z8+/HgkiI8KIjNFwkZUmi7YnWy0/BOmr4ITmsNDnEHPSHg8o++AXRaOHmigCOv2FJSlgGueXYdEa
lNp54z48vH8MDoXnVTsRItB/+xMhCYEg9muErR2auA3YDNg96PmWwP6oXW/t2IEWodGF/TVbKXnk
ISfJ/6A5+jdYPULOCCaRXBmWIJawl/gc79LG6s1iU36D84BzZHFwlK4gsYMFlTB8YCe/GFMBiXky
Hs1C6pSFduC+pj+kUSgEGGwv+kXuE0y4Dj2hwtTRj1T36jAd5byZYh9nxbhDEoGXnl8L58HWEcnV
4JCBbxuykItuVS4I5t+myWoySC3L1PHXx5nq5Pf7maA36GGeGytvz9JZkqpD99pmi9O7cXzwh76f
YcB8XTsZ+4FbtaPs3BSUXC7KB4ORyEuBbXSic28lh2tXGIi5VrCJIcvgbkAiXqeb88akWZsUNIuB
Kln/bhjMRBHLYvm7OtFp9BuryO1EADPkApCaNmFeVrkMfsKF/G1n9bez02xTwVkoz1tGW1AmQPfB
0cHGi4VXyJaRD/860+7AnK7jXdu/j/9NnWGe4F9dJOgL3N7PmRdf2P9HFiVuScCwctF43zjRGxHB
CY3uxSx/d8T8woKUOPaXtDj2UIa8WFNEvsJS84YUD4XFebiZmBaVVyq0KCc8fB+zn4gbdB3tLiMj
PKPsxmFnLr3kMbSTU6oS7IwVEsk17Tf9g0cVdiOVgilg7dFqqodsZnL7pueIHw9YqWK8Qp8zLQ1f
WMVqAikmcLFh+g8xfG7h6DfkoOTQDwG62eOk+Ge5JFVsX3ZC7HhLV+dDknBqLFRyDH8ckDPZtA05
stZd/16SmsQWRzP13qqh0NyvEr5AFV3CYKVqBTKJh8MyWN2DYN1ijVJQ5j7krDHUSTi7KPC9uByh
1eLlDqmvAOjtHTPeMYpynpRTNUvYay7CzOWUB1tdIaYuq0ZK71aG06p6pH28XxvMtv/a223Uu1jo
N0Laq5gsJBPyDCqTLP4SHDZMWUPb2rySr5Gy5+QB+mwpyzLnrTKLVFmnQ6eimYF9PTc9Fg30t2Fa
EzzDsaiznX3ozpE6Ru4N6tOSg27LQnCFtvDZYpt20XeYZ0JeqeGg2gT3yo5hFURIQSbpSMCOp45B
D6ADNqijs2DJK1m9pEBID6lZ5hlbhOTakbjpRY1Hg7l5qPktcIpUx95G01Uo/0ojpXnUqG2j8/ZA
B4EvPd4Srxbf0a/ntawl6eO02fExysiB2I5EbRTK+XzNkdQt1r9Hs7NuN5+OtlcUDtgu1UwY+Xo3
rA5zt7T+R1T7ccQt0FWwIEayth/OTLe3cMZfEuiL0qlr3jTTkV26ysvDaiWc8ouFNiwa/nzIZ4S/
Dgey0DbTS5SEuZEMWo/qw1zUAJbfck2xlEd3fdu3rKVcD7kkKXDezSLiKrvNKt9hxdgp4Dno6LVP
Ml+6ZFTFEiPuHc6WaPWHsadulTiaG4utOcR1A3CAxNswl+alvtKvrJ6IsyTq54co50dFOOF/SnZI
71Aoku0rVAV2XHFkJxqk2ZG+blBfRpqz7/O7aZfjJ32JAus0ZmmDmMDbRCkFV6RLgHS9F0vp8bwq
ZcVnSE1BTfHs5tUH9vtT0y0QGSPCuX0q5YgE9WT1N6tyqWT8HvCXlfX4yzBgnLNO+lOiX6RDtG3Z
l78UgwAEhBN/MZfbT0xeEiaPgREjLAni7mr12ZsSPoXlv78amgQiT9YWIy9K/KX1IPo8sxPd7tDu
0ljmvHtHR+jM4JY+7b/0lRjApWjMMDDZGIbrSuLtQ0G78wAAShXXrhIXmsBapHwogaoVH5DOY8Ta
11CB6bhot9ZIeZBe30rz6eADTI6DMXtxCFTgl/i9v2+o62CpM0IvKhJP8wNb7Jy5Bq1epgIeTDrB
/pzWM06UAA2pt1NhqsJInQ1vluDkxHVEc94xqKuWvOLqmHan0zGyz0xJL8KTnascFJW6Ku1OVMGW
uXJjSHl6U15bTEi2qBz+wHe/x7lPfngihMsX8HpOL4ihSfd74o9CkxlmB2G/3EzP4N0JIYBfF8bT
I+5j6vLZdzzWAtTMUkV7jWrxtKyBUk8gPiUCCfKPoLwESyvEHdoeL/irqQ8i43K4UWGvWwhezJQi
GzXFKMVyk0MGIk2KbuHaf2d+ONw0dhEEvcmDMnu1yQ4KUUzqFotCKfSrgxWTZkKxEkP24qt64hDp
ch9AwXuHBpbFX1Q7KhTwhwR4PyahhiTPaO/rxMNgCLKBY5lWGiUCcQuihTpbj1i3qqquGV1SExTz
fQE2dQGHv4rCOnRRwB0FxyJb77FS0heo1tnq016ZbIsIcKLBEB1MacIltYHwyHPn98XAu5+Eq7IL
ax3EZtAMIy1n2uN/DS9lXaH9jqMCvPRPU5xAmKIDCECxhDh6T0dvbrbk+Ooo83dx8mMG3P5UWw0M
ZbYJkFYsaXhBlhD6CSojAL89bxl2rvcJTgcf7R5J2m6fOFS2qmhPb/bjScrLFdTHlBHyfiDjsAB/
L9ET/RB8c51vYPfSMe0KMIOxOVgHB+Lj5MPERV7FrPSkwVLHugH8yzGPwqRKAuHcESzIQz8Ybvyy
x2lmGsYV3R1FcZeGn6JxEplm+NqGj0mVunu0D++S5uz1xekmGT9wZbm10TrFI+BEa45TJLoM0oJv
pUe90U+SqLtfVlG4HcNQNG4woBpiHFBT6Rz24GrkT7YW9w+RR0avGC6iIVdLda7PU4CXFw02tvoQ
xfaPo39L6hlJU7rF+oUqiPMhDr+tCLNon+vnEoDhvBixxMlDYHaYg+Z1CK3DhRoC5U08d18r0T6J
YFePC17Tx+LsdGUXjJ9OpyAzHMb7FJrxYTIHYa5W6BwV66B5Nu5ahNoQDLpahGK2yRSvPvQV2i3I
be8BoVHsYYGk/P4pwnvfmRq3V4Z1JGElcYtjidHwm6UGz2gFjA2AZ52f4ZGnqTxeR+zk5hQQeqUd
U9zWnjlpE+M7o4gfXj+uVWGdVXhXZZRO42hy9cdfw6zSD3IkMDGvelIDGrUOnOG2fsIN8/dRXddS
F9sW4YY2rwUvxRtxb3CWCMgjnuWXsfhP0TAMPetntoh4OYiP2urth2zZAjzYZ6Bwmj18yDuljBJU
ZLfVQWCpPZ1r5zGchkEk0Z0PrsiPEPP1UG+AN2uwcHKDK5fTIcrIy8rkOeQ+Zy85gunTSdnsBy17
payVLPRMitodm6Pjat/1TQh7CiKPo8OmHn+IqDV64Vb6vX/O2/ljf1EFnc8lH1DBQ+dyykeGl3kw
DwTYKOqNqnTZNzzPveGXPPl+VHr3dqaw1AaVJdQyWbNs8QxF/9YY8Gyt8CpkfY/i/CSMz916jK4M
dAywJ6XmiDAsR3kDA9ceVq3H0274ylobz96M8KKFVR8tIPAszHIrV7zWMxlPpEf6ARUm80RV2oEo
QGZH2ojhT+9ADDpsGugPTWM031MP49ejwl+oWr212j45mlN3lPwv/eE+Jc/STT1JcCUlR/HrAfgm
fk8vZ6aO2uS8p6wK1SjnyCiomCNjU71rw4DKfRuDxdvRiHbVluIYyas8lM52SQUkfecsAcZ1Azbp
iyVUFlVO2dZH8o0h3MoSINMYe7RB6X7mU3PVbYgcTXA4dVaiZYUvsHSJ6BzLW3JgalbZVkOPI5LD
2gCo8k5zNTH9s0r52943Ideb3olwnnUIDn1axtbYOcjX69kn1qVoEGGaz30LZ9frdOgTOn6WHEl2
km1Iay+Rpq/qWqHTYWypZBHdme4cFJXb+6iENApcOI0ZHaJ74gFZN450htAvBU8PGIXoAADTzkM6
6zLSfAuqOPyYEGjmOJTJAJ+oNty3m9XdbEVSaTUatkWc8zrUIeC3uXiGhMsS4HgAmBa281bWy05X
BdY6hFoWLg/u04gAm7hjM+X18bv5/J3j/F2Ya5aiAQN+YtZnsEmytjuxwJGQc9fJYw8Pndvdgy11
+yjxzZo4b72UIxeV+4L9JcCyYg/Bl1yHd2VZBCaNeRfeXc6+frHSn0PfGwp6Q1776DYWe3R6xMHm
LZnqK8EjdEfVDytzpTHMuut0vr0NFmxd75/CHKKy21vbmOkWnikhHolvTEVHrcj2EoN4eohJDlv9
FvoFm8B21WJscLO0o3czkCFZMgkcDtsJJyGh8gqw13fpjXi6cynSa20pPgyKB8rmf5bfPpiXYw81
LTf0+bjd2DX5fN2yx7UXYvPIwM9K8v1os/QNtl07bIu8yrTwndy3Rh1TcTSnEvPj1jE9A0vK81GH
yXiV1jJ4rHmI4LWUwRYwvwdNhrzh9k4wHobFaK6GOxoPA7V/UnnlBGR2cMoXeDj3ShQHu5KooGUh
b5MSzdp/Qzl6RLEOmm1gxxd+KtSXEfhMmvGfnyFyOdbZgPW09BDTkkINoJ6Art/Xy7uJd4U5fkeC
xUfdhaSbbDgk7cYah5EMsFxj6Dxv/n1hd51Am0hTwUlzeuWfYB2mSgSKO226oZdUKL/cns6xFBM3
QTtlDhtBubjXgxbE5MvPvxiRSZZ/8SSSAb915XzrWZGNLVtZTcoimf2bWFQLNVn4dkWODvt9R8KY
LpiaZFekful2LC/Bbr9qkm4LWhHDnZfYc6ICEAsZ6wI4tdQUC2Xt09TnpKeDRGBF91CCwVDwa/W+
b7vkFc6Mj6Q8ebGFykTNa6Q7ya6M/F39cisbYoYTe+H5Yb5vFXN0N9frnCqGtB4VKR6lkv/DkdYJ
jLKX1NW9FhLJaK9lQr1oz18ERasI912BuQ/YRAYswI1FjFofBh46KEW1R3ReKvQ6xlx1YDFkZpEy
nN5QOrmo+Q3xxveFLLSIrIFwDSn5AfTHIp/+HYybmN2GTHu0mU+b8Fq96E4Og0puWEb7q0kgaBQ9
eJPgZMojvgZZSkl5bf1E0g0LHBsQTOIEhaULehehU0rZ37W90L7yRKrWr2nST0mimWpY+vXGaLjz
QP25Rl/e/HY61qNcvBPNo+mendHMO0IJUuKdJn0TvZFjSXxfaJVt7igai199ytYg93/bEHIMqjXZ
8fe5DbbBC9+lcKTFFbZ3HnI8/0KuiT0iXMd0YjhUj450V1QhegczfgjJLpoIp9fApZDc5jbOuH97
JkZZ1so3BnFC/uPcTtaPDS0N1aLGuHzfevRhUVRN+oJGZy4n8A6S1d/EUbiYbtmWcYT9kueopvNr
1CB4jesWL7ASCrvTEoS/j8b5N2RShH58q+V2BI/pd7skV2/4lO11OBsg3sL5oxQi4T76Z7U6vHVj
1DRn3Z7DSO11HiW1czWzYa1L4J8GvQfKb17iFFKEmv+cwDcYdhTkCcQpJXpDENB8HjB5ToHaNr8x
ghKIJ43x6fEdOvwfclYi0wbexjnJhaK2U3OWZ34mB2+Ojm0J0JDyOUlpx+4hrNlDThkCUzpGa5UD
BQVnBexgwd928b/arc4GXYz9MlPHG3Yqhuk6NHbOjxCaU3aOJWp9Usmvgm43aSq+xdpy5uuBLpFD
Ol8b+Ac4AAvTa3MH0a8GuU/oGBpZITW+JOyO/t4/AASpkw1V2y9Vp70+bqL0fDIfp0Yvh2X8Ldc+
Md6NLYi8dzMMO7Y0hONT60iPl23GabXcrBL39+CKmUMYzrhyk4Hc+y/m2kKSgRxXNPZ72yT1F45O
sYzREiMqv8wYFfiSBsO7Eku/iqiVrZV2wJEi2f9CMP+9rt514g0BGJozv/fmxacPntGMvr0t4DoD
gaoEzefYvGVvrHzhEjv4kuchRLbq2sCNrtF1G0+rmQ64Iqm55AWeQilg2XbXsJkjY6YpTIgeD+gX
gSsIa18+6G5yOSKnXtAt1uOS9ulTXPkRNiHyD/C/u7eGk7r6NVpY1b8sLVugPiUysVae5ldaCbnx
yMoHbZr6jHXE1kTNBwC0zeEqNYVybt8Q7kM0rMgaRjRgmRtFDl5b1WT7HNRIDLs7wfZLdnR3dHnP
ybZtMybctjPWWAYyDVv+TlAktS8cWkX37aOXSnBd/O1o9aEtu959aBsBn1Gu/UzbK+dl05pdhdTb
uRX9vN8xMDG6qZ2HFlPiUKPk2yqURsBaAjfWp67+6Rxjejt0gywEHUuOUi5+jT9Is8NZzQLiAWb2
y8X4kKxlBkj1j1cPmY8orCIDqKuR6NzOW9yrTqDqoTZhxT69REuNVUjtUOMfMIyfoYTwB/a4yCWf
h/sSZnENodJ0a4mHAGvkZyCcrzax14iV2qiSGHxHuw04bPRM5KkhNFhdGg1LbukkLabTWpccSLoK
nZg1/uuFZDTqI8eWV9mSf9g3Ck3YerqI4wJJmavMRA8fPVwWS3yKMf9XI8i17zPtzSaqxXizAWix
s+Y+O6Ba2su8PNCF55fXxlAoJOZCLodn+frTqCrPxlc8jEJffWeq2Ud3640n1yiNZlOt8qI9mN7+
DnVJSCJA6BcctNy8zZG0Qq1q3Nw1WtbkK/50dhtBCZFxLHtv3U8xgzJ6IWFmfCybnxmpco3urJOr
A95dourjpzKd6VSwZycQOhkAanhQLJfjJM7psW0eBsL6uqkUgc3WvqjscJtlJCWuLYiLc82i7Xjt
I5T0lHwPCUG3oc6o8TEz/M/lEWQkKiBLGFA+8/KVLKvA0zr8tTZ+1NfxQ7e9baGC73439ELETzlZ
6aMu/DK/7o0BuJMmJjQuX8a47W/bk5opSQZgfY4LfgOcbo7Q9Y2NAMQYI03k0pj0dg/Im4/Kdkyb
h9lpP7T48sGj6C4a4tzWcQzJywSXv8/xtiBeK1eLcZT/M+8sRaT9n9J4Ft8KdzGUT5QTwd3AmcQT
8Tp9ztDziPJbLOJHnl4poLglObfyN88M0uH7qKHnK+2Zkq/Vsb5EtZdawN3ZJ2A0S70HviLWt/Lm
nsx3T1zChRKcZG1bQ/3f60D2LVIIwQlEiRO+aez7tdtY9ltFmI1Kblr+tjHRAXSuaxG5Ww3L08M2
d3KmPM+kTT71mIuUj5n28BebkRfDxKHpJ0pOihMeD/ynnKRzeeafubUACX5LF9nN1WEX18LDQzlu
ZxHQx6T9y9xUpSAEAaUH5XrccLSrjEHxal9a0u7JB9KSn2svTNVbmh96dN3HRpzb2n1qs+7hk8T7
jf5f3x2ggqm8288qdN4ZjqqBmtts7JN6Gl14JIq/tTE9v08bCT4un0hb+jTUhH7TsNB5Ysk2wfE3
sA4Nl/E8zy0sKeMobZPPtotU8Ik65Vxsi10Pe5WQBlyLeAPqo6z0KuBKcCexZEaJvc8pR3YQY/L5
W2dTOOJhrEq1p0d/wilMrF1ZXTrtNMFQXAOb3SfG+1sxDoiiAmZRZGXJ/NAf+X6+dV3D8c+Hat0t
HXSgat9C5FrXPy9uqqncmcqELGRYdr6g2AljXKohQfvMoCdIxrIkmd15HEN4FinPQyDkBlEQwaRS
LcV5+vVlFNBS0h1ojiHOpoU36k8FWS4a40oU7cgQewLA/uhlS3L+C0hesVd6xC+zPBjKnonC2XQ9
my0eYktZshvH5Gu9BXbZgUk76gyE5QlINxOnZY2NP36t1UTc8AubAUXPsYK9SF+vRUbVIP0h+Jdx
GKBhXVVSAT6+XAO9GiUv3KsMhP1lZiogO0jlK243tciMGSapcJOG2jsY35gtWZs0YXoUj6HbG/Ez
bUMFLTvvo8bHc7FZZWiWfMyazJgXfXSuZOtn+9iITX24E90o/X+dHHlwBbJpo8bClvlq0s4bQoFQ
Ez1gRDl0o8ueFETFs+5CJ56Sz17byQnE9W8fD781CPIcZ1RLMPjh8op6a4bKMOntkeaFny/feIlv
sS8HeYdGMipadkv+OXCOEo19RKwKbBqq7tg2qW3x7Q2arqtDV5/RK4u8paZvV7tE8yvCrM0eoHvU
jjQubQgC0CmFwsQfzd45kpNma6/iM98aKXxonIpUs6SXFukgDe7+2liqavOsRI4VRFWyR5cQAtku
O/iugN6oS1wJ04I/rfc3D6pE6YS8+aUzwSMmdBJVqTUBLp3dwCr/Zywyq2HyBGmq0NnTVVInu9wW
Ew==
`pragma protect end_protected
