// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
b8Jm6cRcr4JkpAQ8mwvHBrkMcwoSnRuzR2sbOe1QJuYmHDXspyp1W9kc5fd2koHz
eyCQmJ97DaJXnpSU1GB4AQII3kbU81Yy8+mOqhjiKh6Mpo3qc5L7CQDqPn9LqjvA
lSbpAyahDfis0toP7cy8pdzeFSkeUZp/sLdkuI8Zf0o=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 11008 )
`pragma protect data_block
OIuU1FzRQdcXQph/TTR5kblT8GNKWq9RMm1owQ6H0rzfhyrmio5sD2yjcyQC8eA4
3o5e8eAzAvYA/3TZwCpp/6wqIP8zM07oMzHw2yx2kfpD6s5xqhcPqrXl/a0tYTjR
xi/CuhcLGEg/deAIvnHACWOHbGZBwa/HIC3qJmA4fb1m1cQQYVtdZS/voCvWwKQ/
CBd1Dj40tbMXM5xNVIiq8I0mjrnGd3401HbAw+3TXFxdtwHopNq2D2DPTjVgy7IW
CaRpyp9G062usR0+2DnG3SwLcb8GxLa3wMz3cLKwO3zYujER+o5T5FAvs0XTWbMJ
UlcMgqjmoqhPD9rEPiCWS7HhCFLODsK7ucCL7pGBTE99m6A+gmf9V0rAicHsrGEm
tAlsq4ZJxcI1icV4M7ZW002NQNYBENVjrqazkGFNrDFxCxak+pZ0Ec5QGLNMY400
JjIY2n7BHBh11DgWImxJ1S5sh4IyDxvOz8KLx/K4udA1UTNZN2gqdg+T4CUr9pXh
7bVkPJPTS9tgZTQPlyVYJlO3BEs4yBCJ2VYrHbzfemX4rhYiAyzJqXQcGnAusH77
6yoTyPQFCp6sgKufBaLzSoBfK1/DQi0EM/mFSmmwmpeN9PJsftoE+Dnd5x0GiFIx
xi9iEGRCabzIgNB7Of+YVwLq/AiBaaOztKLMfqfxdUoFzJlqYVNvQk1cZWW9YTes
IiTGkZQ2flaTIF+1mLGaaXfi+ElT5FCWfrTY/ZpbiOYbQE2fAGjsQMzSYTzY0fCj
RaokBOIep01Lc/NG4jLVSYyF8m2YIqDpTk0VFrPeFsEUTuaItHuq37PLJHpYK6+P
2bvSmqRjH3pzrcV1yHBn8L7Wmg78H4tupNqIxkSfK0PTArlnR45ea8y3s3YJhWfG
W5HYR/jBuKN1RiGZts7w3pzhrgwNBoxx5u8MFnr2lr9cSYeMEzia6VI8gLDzc+Ks
m00e/zgi+ZIuN5yJ6D9hXml5u4kP181v6HWlsBfvNzuu5VhaBFBnHbpbKPw3SEc1
vT/53BPgoIEXUXeDa3SPjDub4eyzTVteHASogt40bVoJc0c9uOtVxFPwKb8Kbg/D
HLbG5eL1Arz9ONfsoMUda5UPCz1LefreVeU5UFFAHlI0WjQXLICKGX9sB7GacQN6
eCnjF25BmebyMylr/x7Rsge7QEJzWLh31cGEB/mS7X1l3oWzrLUUafDHkqb/oSh4
zHG76VtHhcIPJ6Nn2rUrDg9crRbqjS754/X3uzEsp0iJa8cMi/BrYNS1PZ8EFbfV
iIqSreW2lwBzxFW1Jf7qbrt5jKK/RExKVJckRDx8XAvPKHp5tjnlthc5IcOPQ+9Z
V8Jx7W+9b27RITPUnWVbeeGyFEszT31/RRPGloCAX4KUpdT+NN6pxuudSiK0Kkb3
fg98H36vzmL0BkH+zaFjXCMb2ytZvNEwHfcXorXW8xlX+cNy7dQFXfnWk1jRvR+W
tiTXJVsx+XSr4IcwzGLV3wMNEWHPcRFtnL9gGHYcmnD4OB9+w8Webbyvwkx/jNTC
PhTl+6qTDzoXReMxLP0BZ2kgY6xGtQLONJMuvJpCrbZ2BL8Q4iFb16asx4UeoRpT
56qZWj5n6T96sPFLM/gBk6sJ555SQNyrTC2+A1zu00ipoCRhhBZVlTxvREuBcHmQ
GYOechsCj0BU6ti4c3E2XrGYnQBEMVfrV35o59aVFq3s5aealGYOj9VoPzVNfYr/
EKGRX8DEYLdOTDjjzs53gZUjuYFx25/uMJATAEWjlP5gxSyTEF9OU35nWtIaWnI3
8VkBfBalstbLNkww32EF7sD1RJCNlK+cTXyFKQJ2EyLqfQDCvcMxe/xdgHJfUzpd
qnvaqNjHFRrge/pJLK1hHl/sqp1L8+PyJGxzBEnt5025UCLbO5fOE/v6RnIje8wP
WnUlhKu4kQve3lSIesgu+OQQjIR2sjVFGGmvuh5/DSph0pJaFjxyM9ttok1X53lf
GrNOyQ5Qry+qCeVq7DP7ex3CgN1LP/G8l8VDJs/jhSsS3iRsS6bvADJAj0ZIvIcO
JsYet3UfNYosVhSo+RwCQEuM0fxkm8RFpPUgM1PYyv89aTb1FgNGa0nf2sIwlGSx
faqWyY0Z8xkjt3DxzZWTnan3q4+fFWIFRcFzZJYptXCyIND6Dck+ofbR2LnUThJt
TTduCTLEl3BmjXMh3ACByKeTK2DgI1k78hkrUhnIHvIRSzTZBaLkfNiksqVMVd+H
tZRXTTCjRJ3IR95Sngnw+M/PgNVsBm5vDUe9iy+DmtOPgk2czMnAfp0+YLg4JW/P
uUXtOyOfn/k9BqTRZ4hCZKCQ1qTrvZhsFsdeVLpeoXQV1T7vqaVgInr3h+FtsEed
KBuB3QivEoAU9ZPtx8TZDwziTOulKiRggAs5LhoMAir2+y/n1KerkrlaHEM1h9Vc
y6+rpyJhdZOxbw+EAdMqB2fgX4Upb9PwSgKBeQ1mnJaMtaNYStg+Wg3Ir2ySt4tK
fzl0kHRpKaiE/Bx/3sM7cb0dI4HDgUeaC41YTaKyjARI7Wsji7IDIpbQNKuMS7/G
oJI0LXlX/2jZGCqpvtnou7cO5VxoC2Ffh7OhIFZuYRujat3fIfiaTAuZYvZDL0ls
Tz93MpV6Oz8ZwS78C9xvA94L+Jc91E3S3VZAIO0fbg3elgUh2oJdUT/cjSGh/MRq
oZGi/mErfJyYoKL+m9BeG/RpSCIm+RS4W4RwyptmxvBLh45bYKkvX+Y07tRFkEjB
cCusSeOYMHFaDraTFJ9AFSrtEfEMpSNSUrsV+DzAKlq8WGmJJ5EH9MOjtG/kN4aS
O0CBDmUPCP7yz3AkJ09PRsaEbP0XgU4MIhVBGGarig7xIxco97+3E6enWVUsOQXP
rIpG50uQt+UG+PsY+/hY9p7hJmSKOvLqFR3z1rCzqsoLRFPVjnbf7mHJ50xcZZ8l
i30KPTmuFtgpxYTsDhCJsvR38JSc9qmzrpQz3Gm33l+guqdZ/XbIPrgS44xC7UjW
CysuPxQSgAePZoDVRyDMPejwVaYUd9r2aUDWIUdytMavyBFH+ZJMX4iNYrad7ZaC
Qjdvkdboq+yH+f4k3CywZx0EF8lakmk8lqGcSSodZ3toiGvEN16UP141qno5GYAS
hTgQBcdP9KPiLBa1SDnlkUphhIcWv+1TWCIKtQSei+a5+Jo+UWmltBzVyctV9bKw
aLTZeGQckaoa9514OoYicFcAjcuUh8LnmMQxac4iM7rTq/4l80xpX/P34c8ht6On
PTmyZUCq4NDFj9bAhunHnYwVPtxY+UEYCeByThQzKovA8zKUBXrnv2grV27k3vbn
UIQdPQgh+tn5ENeRtdNhXmtD2+NNXHQq/AJG8VuhWNqMUmSDywZJj9jei8mGRELG
Uhw5BzbziGvsxZc2QNvZ/y7BQSz6VuE48nX2BysIjLj1yPMAT3Rp9uSKhWzxo4BP
RgajkMpv1LrTqhq19AEd3jA9D4li8MTfO52OwCZTbrPgGB0Db201PuvExo+4spB6
mofUKoKoZO2OJbeuaGqjqybVw0SDXujtAy4YMM9/jRR6F5g6fbeg96APJgE7tWvU
eb5VZQGy9S+sq2QnlUgJg5Uy05DpnqXbAtQkjqzWM6Y7ImgKLPSLMxdMDLFvGwUV
UF3DrVEPEjSg0YhNmFHL+nFTETl2P37uuGdqlBV7iOFCOt6EL+L+oVfswOt5ad6z
X6F0D27BX2gN7HRRrXhHaEKLGz6Z8nPmQNNepIWkAG37FIaMJlddnc1d6G1nbGPN
hqdhRIHGUotD/BZ2HaymLj2o/R5kiZ3YgWp7UU8lSpEUdrjtWpNeMl914OTqg2fi
rZaaGemKphI54KQbnuzNIpKNkZT+ZMdzyWDIl92g0sGK8EacGpjIQzvRtghMaQDg
SwxxuYaGfuiPzv/CB8AmxeL6YGn2I2gf79NB4ohyKiFmyN6z84WdWD+GeKJDw+Ae
E+mwhbSDw6hgEuoO+wPiWD2GU0jWr+op7fdA1Oxn85+yFi7oexbv8wtFp0Dywz8w
mlRedDWEdUz0Im9YNM0FXZhbPD/VFzLOnDwRxywQoRr5j4wymridSAOxcRhoOP9d
oUfLYPy7wc7/8UTae4Ua1/DkAiC59aFKqQfd7aGlaOEMkhASnTHKq1XjHKDVlf/7
xZ3YduFMVS/zA3p76d4x+hWhRqWNrlGBfB+WGUanhE9ILY+sbeHRtPUe/noE+yre
eiiWltt4MBI55Li4La0vm8A+a3+s1bbOVQKgUUFRO0iPKG1WSPufECxQBv9raaJj
VvGIppTwIOy/rQCFv5v6B3sGv8iyD2baAtF45fN1EpieSxje4q3MD6cqzQYW6veT
bD++z3pZBwjtI9WY/EQwZFYmdvPASjwo06TmTlkkxJFg29vFT4+zveWWMIzL3oNF
+56E/HVKufEXTLKHtYqu4yorx1VVF7qStbSWDARMss+fnF5/jRe1weUby0L8fGyl
DsxeFeQLo/nXQ2T0OsPzz+zIYLXS516g/WmSj5YhUj1iWBTTjnPJEzaHj5J3jZ0H
NHruav+cJRjTI1+oKAdVGuDVsavR0yEkPzhPKzrB4odWT2BV1EyB7Lmqow+C3JHf
slE4jf+wFe89yqQRQ5ngvDiSrcscFK0mNUzfhNTYDTkZfKMEjPWAsiWgQkKXrPuZ
NIEHL+TpTT/b90up0JCYpchY9QfdK9DOTv2a8BNXu3G/43Br31E5h65P0aK27Ufk
8a+Xc8nmrLQI3/1fP9AaZBCge7TIWzXhHmEZPB+WNfbwLYKISzAWuV0+WW0Am386
XjR8OEd/gnUlia4j3r+m8X30T6H4KxeAapc6iCutyASzJ/8scU3OcuwgdCZiDpp0
MSaUC/RvbI1NiK0VBtlxgfDn68bNUQ+1jE6gaHCLTcqdOwE571RlJFOaRsh1Ns7C
57FXmDvHpnWjvizMTsQudInMm09tN8cu5dsCHyJ1omu5tr/QS/S/Q3gSBGTckflA
r9r38XWelZTNQAzu8GMvBbJinTeBbZcWUHwjVbhbWPFFZqLN5ASsf1ZSGKVEJrZ2
p8lIGvYZD2P1U/UgmkS5vy0CUYHOQNu85qe+P6IVDVPjeV4HSkCQ4gMgFgrA1Bh/
PBszHe994hxox2R85CgclqC3pwvFOX184wI7XfR3VoRC9tXAIFCm3jAX8iM08Vaq
66MuHfkZTB7WE0vgTZ9gDzULfVQ/Eh8eTNBFHSPiHuvv1J2POHNsTd7V+8erfQtu
hbIzEMhBAsMJU1CdxwLdT3Dif604v45kEbOX8a+/8EpQMc/RckQQPQ7lb2p5u034
+CjOCh1FVdbYwi3pIlGy7QBbBIjB2XZqUlyRxcfVQCoB94oG7/pVATY1xoGPzDev
NR25s7R+ukNwNtfZYdw6D3tCa6An0Hi3yh/W+6mt78MA84Ab8LKx2jFYIH4xRDWe
NVhUUWltKHp4mpADlCuHFuIv0cHN5G9RciiEPlAgsM7XGCtaH8fMiCpz8oUv2xMK
nbzLTu3CR28wQpuAunLknBK82jnMc5CQbQOtWKEy9GUxTz8WzWBD7wbNe9z9npF0
y+TvhAWcfsypuoa9V4GHKsil6Q+NTuKTDOIKyPOz9AMR9RylJDBP9Y5menbazAcN
BLmoiOBf+VRnyX8gAQS+odgJvk98B2zAB26u5relpAIWOc/s0TEl2g72oTHxgTZ3
/7IwlSQhCJRPv7dsRRJ6rrZKQZ1GKmzBi8tvkIat6yKf8Q/+BBG2NRX9xw8ymfGW
88+7/d2CWl6e5wDzgLkJQG2Nju0fVfOeNBdff6MggZJPcfliii+bR6KO9eQWRO4P
Xqyx1e7biyFV0yd7uodz8wDWnLVvL5z57OxV5SJp7GZXlKGdiNPRIvl30ajOt/15
vTVJ9y+oq9MEOGS2nb+bsBE92i+KtbEzvITCjinJvAfbd2sBNet2aZSRhziLu9+v
zoCNz3ufO9T9Cnp/pYUzEIza+tKPyECY/MPfM0TBbxQCVzKaKxAhETgL9e5WRshc
7HJHZcD9D/B2kFZbXFsU69HDQ9yY81rcGFAseLMa8If08IsjMmVj61uKLdSt2T7+
xGPVwaFhsajrAeESl/v7IBcbVtfZ2R9P4/eefvNVWn6LBlQu64uxieoThzICG8cV
TPd5eJo2CkgCRG1cOxh+Xu8tpj15yDq63G4Mf7RXV2a3h/u12kMu3ozc/es5Ss12
Q7Jmol1S9QPCW0F9TH/Acy0citJ4yarBO9ABGnAdzaaxE4tT/GpvfhYhtdLlXopf
OE8onW/Df1h77rsq99QIu1K1kqcwPl9W3TBC5vdG3rm4DqD860W2Cszxbhq1PQtQ
VFzKh/heKgYKH5Q3/6L1d1wHZHam5HQeMp8513WkWUv/CZHrQsr4gcOPyq5xqa6F
cSx6NndzXk4FxImSLB+5jUy8UYgB6tt/WLJyFIVAIJ8lRP9GTObqtWYMfBC3i5rK
bUIMRhteXa8iG+VtqCYnGV6sFCqJ351fwEykEXZmP5etaYOqA9WzieWpdodq8dxh
NYe8tr+menLgg4pAIdABgOJtLUaKnkXyVPqRV791tnwQ2cgOb11q+9le8DPTqDfh
9imRqAe7FkjxKW9Bxhpe8VUGhcfaa9n8kivBftCjWOY5YY+KMLGbrSEtilWAxv/L
69E2xeQc5gMsmca4zY7ngTTE9IsKK2CAD+jdKzWPnE41wQvuJ07ry0hQJur41Cbe
RH68m6eALkLQh0gymN3uacFGpVr0db9QqZ29S+j3E5ILGBx99bnoQhASK1SOpPEc
X7dnGzRU+pKOkU/77r2HMmkklcQC8RbRG0+U+vuNutidh2ioRuNSHydn9+IM5XSj
PvxUTEtkO//HI/PhWn6pR0xcxIU1A/3Ly/OPzWd3knYEHOUNiH3U0roNCRCEYPlb
anfzpftgCQ4r3gAUFNrRTPjMvE56R4pUskO0nbRzkt0KMY+S2Sh6aI8iIuhJ80Hb
SgxP0tdNL7kL3avffY2aCZASR/S66PFqleqQdLTUfFgnaDN4PllyQtWkFwROPsZ+
sa7RcG0hRhKONHvL/UGgzbtwzLUQFf9Eo9Tc0fx+flIhxAoM83PBDqG8mgWs32ZV
b6+XS4G2HvZ4XWbRnK/wiQEZMuTkL+8mL6nZXtjPzvAeM/2EhOJPz6T33FUPy9LD
eIzxv1saxvAYbsLat0ghOX++yXMwmeH3IK+SUcSbE662WEYlb1FYgnY1rkGh4EeQ
/ZysLG3sUYG0kFdcfzXnMuQRm8lUPIC6jrUTeGLrISUooxMm0G5ylpEP2bbd7YuD
VZZIpBVXXPGBZh9+oJ/WWqlQVsK/0fxfJZLCdapNvyGlPpVfdHrWOXRsfums/p2s
VbJKYOfqHDAEb0Kt0JsJUnDu1qA+xPpmGzPcNdkeXQE0vejIsMgzcKnomPq/4EKT
5ivVVNy3ietnsTuZARwdCFNan/88w3uNe0PinW3p7E6vRsGvfK+JRoWZ4Q/liK9T
J/GnH+xOooTcjDm4HhTFYr26jM381kWTQ570kSyQGeOjMBx0UBjix7SmpD+VDSWW
PFIa078T4dfQVa+kQpk77mM9yICcyYsCsULNyC0g0pLvAZmI2ckKbM8h0Neq+g48
BXF7EDpHjwRYnCOCYwFxQu1WwzMuWGh3kyBugy6BkBiftlhscsbQQa7faO2dkAL9
f4AqPE1g1U0/jsi7qADykZop8HG3TtIcP5Nfy59b/VIPE65vV0Ms1yGt8cwpNNcf
iRdjVYleBPpZJEpcYgJgAFLj0bSMmhFRfJbXuJFOEC63pC7EKXuRj+ns1x90dtLJ
yoIvdzo/GI5cxhAh+M+AU8BWKZ0GsaRnqkgQ9tv/utxyjVevZQ8zpndylw5Jf2cf
fpHvoDU+0ch9zIBlsGHmnK59jMFE2lc+g0+qiyOkxtblB7r6ZVQQ2yeD2mXCAcgd
udKvlHi8tiwSyyTWyC1qBGsCENpL6b5B0ut4yHkpKDf08OkDQF91LPe7tadlUNxs
FXBAQ10i9cJ4bukX0mJ1w1H2Xen0DzZI4R65GjLpwPflqV/P8/YNwxY5JSdUUjQ6
eLVF/s4nM0gK0H62AdqIy4NULZl6arqxnW/6+bmov/Zj6fuSzuFN/yCwhFnIarIZ
yDO9Tm0xgjFlS0l+ndf/01sbTIMXNEn4+4XhGCVivUJoo9eFaQwb3U4vlWGtFpil
H8knqVHK2PSLlrFp8FVWKxuGOnnL46kU36CETVfp7CLuqdRZOo+zbNhIlsHlzZTE
uQZWT+nJ1MNilgw2Do89eHwGGsXgiLkGvDqqkb3zErEBtIQgVJORxcOobRwPM577
3eFDon8nylNU1l6yhY4I1d1IjqtplRBTYWZm7hki80K1onU4I2dvx60dtK2+I1Z1
JssXmRRgBuKes5bGureunxJSXWM7LO8n6K/CJ3HNNa2uGleWSSlnH9/4sTbAGW3P
4Ywxwq0Nl1JWNgfeqLjsJQh+aUKt6eb13C5cT7oisSivfT/nMwMDrS/+XmsgC5EG
XfRGRWBNb22/Z+Aq9/nS1eG6Yng1XnIGzcyOfnIY3/cfthfxILdPZxmfvMZ5GWDq
fAmjQLglIEs5/nGPW17UKiyqLWmyUTdvbRd1Um5gPXUCqB+xg9dMVwE1YXjDPTle
Zt4Ho5pgO1woczMfIYA2PMCyC/OyyQ6foEUl5yywDXDN6gp/vnaUYEwakVkrG32J
5AYNeLasERmwj9JJKRmKSF9H+5NfhPjFNDexfVZvWtqSYX70SB3JDfJsyfDc9Rrm
vKiUBdL4W/nBratwRCm+DIvbzemWs7GL7+YHTwCINeGSaFyycOPLcmz1nRhvSYmA
FYZy9ZgA7U8zmehjTsCxayOZulV6kfpvcOGrzn7DlSH8pLXYP9yDn6wzlD0x+/RY
UcYDjdN1bTVu2neu+IfJYbqdRKnaMtZyvPcpx1ulAGV9vLc/WrMADtDSRbozRCgW
lIR6n4OoiKxwh2aoZUGrrIxnOBfNx2BR9RnUBU9FObB1zoQEq8CBfYbSSaV73G4+
EU/JM3SeRvOC5E8hJHHcuCUzARaEVKidwW/ZJKg/hpip5z6WVSHgQM+yf45aq2E1
UR/5giPKU5opLNGUQN36gNX3eYP1CgHTy2U2V/pmYOOjfTSd6tD+DsrwrVf41dm6
9FdWeVVAlMMk5jwPlE+KknZbPOanKZseNDptTSYT14DobMewkLueWMr+kGcIqV7j
/W/91nVrL9JGzmEvQ575NYFMX7Qv1Pf1yP1nqeDJLqeGKvPxECikcGX/nbEW7BU/
IW/TLVWbqf/9fatakgZq3xrcRMN4VXqZ3RkByo9PsNCrqAhqKvm4k0RdiuFfDrj8
JvolH7hJ5lIofn0zTsdm75X6monv4386fmtbu+vAv8yhwJU3n8ed4bTFupU2keuC
CGCGaa35+PjeawougE9CO2khDaTQzLWe3jEQv9f91XeXeajh0++WF180Bj6fNqYH
Y5iGp41al4GiRsYZ0sxeFOO6l3eYC4hPYsJc4o6KFOcYPpkec/LQ1ptHAiF7QyVA
iCM/NhoZ1irWSsVuMCFTvSKfFVB6GfHS5qMziLcjCvIFaHcBJmbdeEPvDrA/aAEs
n4IQ0j/D3y+b0u/TZu/dhJyhHlGZJH1aZewzFIwelKB+Y7wODnt3D7EW+X2EFtRz
KZ0CYIB7woqDdhCMf3sgnmmLyGOAAcbXMNkgl2ydv8phTK/5Jk4nJim3cBPFHifx
H+F5oTViR9zU9cmHDFCVKMIeK6a1oVgN6fY9x5igRApj0QOgQKvwdr4oVOgXFPVq
9T+JoNSN5ZCWNyNKO7yf+KY23P4KhyLe6/ojBZWcLF+QRSpm4CejDhpCX+y58+hJ
9qvOmUHv+ORgYw8AgQ7x1AP6QSjj1MMF2nQJlV2416nUTQRAyzxhXqGCxCAC4zUw
e5gD+O99q8Reb9IFzf7TTDYxX/T74NMOyNt/OZcozWd4w+wlLyYz3sCQcigAQ/Dn
TbSBGdE1e+SPbuJMXTVf8NodipcN7Al+AmiZob167MDgW9+ebPdMk0oNn0TgEIXH
GePDu9+fc7gkl5SxqwHtThk9hZgrMPLZik1pukLD4K+oLiBq4oVllpNaQhDsqie2
HFwOLc/aC0itBRGjcws31tApr4M3SGf8oj456KHvg8Vm4z4DrAT17g5BCd2zV0wl
5RLsNKC+7bXDVaScq8hWORk0tsw5DahUpVLP1k2RBw2Zsya/qm25+YvWFXZ1vedH
afftcJfvoeslLUqIn/qaFk1jlwXMKzV9vwcYJa4kDTwwKaIiva7C2JPjuaKV28oC
7uQWfHNAH0fmCGVyIbIut5LNAMp/WFbQH42B22C+6AqlPIfkc1dJ6HIfTEQGSWbN
9oHgGOVFFnCSO0981P2IdWs3RSvOuDTtU5iFLGGhp+uTQgWqvg4pVccapLidXuV4
VG2itVr0FpcpVZAvXz6kZhDFSzsb0ASRkVw4iADxoPwYEFgPeD45jKviFmW8BGJW
U/AaA1KFzjPYsjPspgJxlUsFEt9kX0uHp0NCMHMVIjzf126aEkKEXbw8fKdX8c+C
oeVN5sVQYZae8RkBAlrE1FxvyIvtkNgiZ30KXlB/JLLee+Fz+0OD3ll9ope4QWFX
1D1TZbh4/Z+7uwyJIfNtWfs8DEKq2DndDWhKqNQAidqUHi+2/mSofhxmyx3DLBpE
vpTNWzV8QSXMNzpmxelNgNsmbCBuyi7FcsWeI/LTRpu1S/JGAaO4fpJfhyEscgZg
kM/ecrYj5Z+2VfCBNXfBg8WCufyz0nGrI4uQudpwQJP2qGQTVrjAJicBgQa5RQpQ
Up6xDFIyY/3AWmP38+Hf0cmYjObwfNFrw/mZMiPqstj1fPo11jDns21tP2uYf1IB
HR2aoNOLSmYHJ8YWOKQ8C6XVOw2K8LkVL8P7kkG75L/rb2QGmOClDvu0udd4LYt/
QmskEO6Am9ZW1gOAlj9ivwFzkFf0E6uFAgkw6RTba1FiNM7iT4KDqrNRL4ph8xVe
5gqhXQmI++pl3ifhTv6sHvHO1vaj3Px1dwo+HlRzXs+mR8kF4ah8ka7yzCeY/51u
U0gPMIhmJGLA199Ynn+TwocuGSfgPGRZFy/I9lSmLv1SdTZztwH7B4oF/ZgTl2jU
2LcPQSwIlCdO6pfV/cDhhcHZ9PVFk0kSpiEHTNXdECS0o/mw1pz2E4mQYgWMXx59
UqpRZZKAhTUodnLsA+vhW9iCxlNwW2Cyt1ReiB9j6XcTwR9bCr+lFqfrOHJOE25X
coMLdY+g3fnic4tbuSg7SaZd7s2gAQSU85OFsAZHIOD4p8yxIn27U9mmkdDNG6H4
ymOBoIYTxOHwDoWBvSJu3zlkUbVc/5vqmvvn3g7+L5vyV/caBUvPnqS3ZHkhVTLE
Yr51pjkQMhBsh+dFQ7ZSUtrC4S670IU6hbHsI/6Xj4bq/lO5PLV8eIt6groovKC/
ZqYKDzl1iDPx/39DPFeAQtexk9R8FVfxTnxxbe8/TtkSNuh+lOfvZO7U7qaqFTLl
kT8T60dH0SgDFu5sLgJ/pvVD5kwGU1EGpyKK+U1apgV+ajK4d98BYW7KurJujQ+Y
en0IIibZQXkCTZTqAVr8B27IPWnT2ZMnVfCCARdndNC7+4w38MA1MTmkvPw+KKVW
gOHiqlZN55BUmShqC5E8eueutGrTKQl5jJEnejJN9RRoH0b7OrMZrY0+jfIM/GGA
Cccr8qFG7bwnyjO+XM5Aes/Vk36/bO+cbV171jUTzicgQmR65skSE1BLyD+Hph8q
e+O8W1pohSDDpOpsm1sHGHIsZM66xE8ng0qL6nPZzwxvR1kmQFJsNwYHfIGP6mVe
jZa66b+XuKvKGhIl6yTMALpMMERRbfPr0JWvQh+dugEaSbq3rcxIlNp73tjTt3tL
bQ6QqkllDepNFX2xLpR+iq04EEaThjprD9XgfyJFycE9up+PKb0iT00VVeozCDOR
e591CTIIih4rEDTk+Eu54ZBlgTki8G5eQOYFlBuRfKYQGahseqw2HA2Qlv4/LOhC
leBKdqMs3l0yb4dmtpOg3EMX+YgYSPrLUB4Cdmy833KZYfa39tcU2A0Qxhopd7K/
q6eQIEBIrA8XCCMaAINpCSer9YV/gWhZJv6eIvyEPJxYy2g0k0P23Ta7xLxC3aYk
YLSB8yxZMgh3LArAMIzB6l5hQeoYir65LpNlfhuXmnRpsQzuggInjayzPMzSw2A4
CBjf/1WDAg86OiIE0gfxUaW0YY46DDvEy1gAQLBlYfIaF9TNjRXuO1NcWw8SzQ2a
4QovzsJiCd81qdCyanAxl8Ly+rC4QhW4+BlGFC49r7K7vnI/pF5KX13BDxmbbGpb
Yh/GjmO00Yxg090ruS3rX48RHldWb7Snfo784VlrifILfd2wOleBu/A1Ai0ASb/y
PdcMQXJqH0QJW6jYq1E/17x5fXxdxvP8/y0Vce8sZoqgmxYKUQygf4U8t6pjxXGG
Ac2yLfWAAHaMd8jK43CzIQUV7hEPyi0H7waESMUiJdY43EFRY2bHDtOlzT7VeR/i
oCqZussWJKUg4eMPfYNxEemEMYHq+VQ9a5mgTyA6Um06sepo5nCSLZnUCxCnQL+E
/VPrH4YvKcaHs84lNZcTKK8AJGG1KmrtFqJsu+g5ymWDs/aVBMavGotHEFY8wGRk
tICfP7p6HuSKbXI4DkjnuuiDXsSZXNvLEeOQdT06D1HWJYqcbf2J3o1B8pTzHTSG
Shkz6FKj/Aw0KNj+m4kA1FRRfN8smLng6QsipBM/puU0TKonobVY5NwTsbdDhsI8
L3ogXqUn17d+yDanJLnCwdCon+MEWgtjafjKYQnX8kNeU8W2IZVWQoQCHpgFFVkj
9SMo8T1SCfoTYnvcquXRk4/QAZz9ToavSrHodD/OFbgcSck00DB6TJ/AyVDEV0mJ
W4ufSeteCzsgl6+Nj8OmdslwAwexMpRf+VY0sGT/NGrBGUvlnfvwfFsSVQ2GeDZt
aXrOevHCKAWBKIqg+9UFUuCzwzwcO6JDqVILFinJCahWWpKu9TS+XUMzLG2JZaU/
4voAQOs/Ej4qAQMSPRQg88T6BGn9blcckqvEngUj8TT6MnHSIKEizmxI4TBSAWso
TNsaTGoB01VqptMorsSszGJmw+ubcSvnb63DUJ27vkHIEjxJ7qA5US5BKxWoPuz7
AIMfey5gQltcVbTRJPXktNaNEuhV9Zsp+urtU48xyMPx7dtu6u+yZJOFa0haGzrL
dMXNKRbZsJhXFLlrrZJ04s7ryhAHrOfhTQIQ2vdwtuzE27HSUsG0U1AmjYVAcpMl
ndjjL9v/t4wpnxOn5G+6JNOHirzJLVHAy/PjzKliQ7ICpIJdwlidd9ow8mjJm290
pyyZ1RlzKx/ofe0WAnYTPsq9FsSIG2D2N4lRuP7GCZcQ6rRa6zfgCmuJpQ+YtWwf
ECVZk42QPqR5MZL+xMalarrK/nO0B4rfSre1Q09G2HUmH8RYLRDsshn+HHTkzRaS
TnS9F2pY4cC6JRWcMQCcDFGR4bWUrLvJm0JiRdlp2NG4tk5pB/Byz/vYiJ4qNF5K
XKRRuf5ZUQfPXAGeo9ZKA6B7ZLGOy1n0u+M4dR169y634DcsMey2p4QKu9hIrSbp
4gVx0EEXr8xYhcWQcc783HbhqlO70T5JHGty3pCz/NdJat50R5wifRhAhQpFFprn
rGaS3dNvu9OBNAk2WlNQE68u3PrHs2Uqldn7fTeDx2KTMe5LKXf9/RgtvM2SEkI0
+WaJi4c7vcj4iUAzjDgW/+EqTWEBtU4OaOp1QhyV638dYqjM6ZEnVaEprcDM0jOO
vD5OwwXdBYT9xEShQPMw5mCx/NJ2bsyrRZ5hxMEmlkkwSxDP2A8eZ62w5FGN2DPF
Vkp0Hy37m09L4xXmo8WRcMNH2urOzMZwHaJKt9aC4RpSE7hInWwqLwjvDPjcO2+6
y07iWbhgSjxdY2oPhgPKSm70R6vT7ditR/p2X14JAITqT+IFulltOAVXCgsaH0jR
cWag+b02iK0ocijtkJzmeEZWQCjbAkRzV7gqv5HS8R7kUpIw9JyB2Yta3rv2sqV3
Pf1wpqcQnP/Bu58S+HpSqcwYfwRm8o90UwmcEUFXPONC24OqkP7wd8dyaRkYZhgl
2Ox95vZYsQhXtaskqyyCurrY+FMl4HGoBY9d+WKLIj4Z9/Nijx89L0udi9RUGzvv
tBoCShR9b9HwpaLDCZJyA3JJIADQWane+BUvmdYgg8eYUFcNMtPjV04cURpLswIQ
9klQzgjVlVNy9kb8i4sW/W+mQnORVBPNG6m5RqMn8NyOIi4ARGxUQnYJsE13kpfp
hMDq6rtrMhQvaLkMvE01Hjhh5qpgCJVLijCBFtjgPD9nbzKr6ai5ej8F6HLPDwTb
mg8CjQHSweKOOoyNWl9aUp+ZTfDn9rj4hlB2IsVRyucHfOmqPeCCrvlwSwInvcP4
qCtheiUbk0VaExARk93k63c6TvhENgQ9Gj6S/deG/Lrgo2212bhRCviJ6zrrT8pC
i9yaNOvC19bV+t7p+wpRZ5P9f+VmijdGEDhD1/JQMjk4AsFEX1uBRS8EU49uxCA0
rOOt+yd8+3pA4pLzEMGMap9d8xWrcdxvL0GQoZz+VPG38YfVfloXoLqFXKvBVlcz
yqun33vTzDEDr4AAgjRdfw==

`pragma protect end_protected
