// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
C/mtzLqMqFECH3Rh7NDU0pxJhTbRE2/i/p7Fntur+XkqSwth7wSD1AUdnXsUD74JDFwvrC9/7gmo
5qmiWWmcEmTarPZQYktNmjieYlZeYiDgjodBioRLWyIXaYe7SlnvJMbH+3SUY/Jwhmwbk/e1yojd
FnAd6PSagi5Q8ZpVALFpmxCWVwncQaNfdqtxq2UcZppBfBRdRvyzws1SnwcxKIK03LH/Ca1xoA5T
nOMBXgTSV0Nx+h5OeNC/vxmNb2Gp8hZBOwKHk3ETDV4MTOgr8VjMbaerkFF53gYMvFcpht2w6GCD
5Fbu2S1aTrMwICI8Ksp2k6VK0hw+cnqDhZg5mQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10656)
hKRqr+ii0N06VfT4pHGnPgEHVGAZcfgMR0dEEWIGlm2VAO7JBLEz+SKTUnzbT0YcbuZ2z8jNjDmu
F9AJJaWhVA6x7pe5JoTQCXGPKahlrV+D/7+ZTsEi9chdj+owNJvUe/3El6fuvs9Agkgp4pL5awSP
Bo29+1ObcggtLMF8opT16hpeh2kNkZDSTHI/yUBe5NCCuw/PRKr4GugE+cFb76rwHepj6OXfolWs
KxZLacu7AauVj4qf4QjwgYHeI23ks13OL1O/7pVkIhLk7IQk6FZAPq6wHN6rWZx8Xmguekhbjtbh
LWvIMYJH4az1uIRISkC4QXSwG2xRYYnkljjiM/mlRieA0TiHANm215BkdHYgny6gFHN6fHr1jzIn
qoM+HldDTb6WsyTUsVt6IzPzYcBKEx+vbqWS5uyqGfvp//Eh2zo6OL6ov765u3k4+o2AuqYXKTSh
J/PsXU1HS8SPndWT5TNjwh/6a1eGM/0CfFYxMPZ7PxhziGkA3Dh3z3VWKEw9W5he9iTsUCgfOOv7
6WmmL6FvkcHPbJZ/SpWiVqsujIjzEa3qPiQWiaSjCtISTO2ZdnQ3oykVt8EH98Uyp31WGH62wEjl
i2qhqaqBbCGIXcACze8Y+6bBmxvIUVn0kOgypYN1YdvdS/eqtSYRVWGSZB4v3kTFqOT2wRuo859j
jZUfTT8bf1GIsJP3PS0+LAsDpNoBP6H6y3V4j/cDpsdki7XtLas82cXPbUz3e6Ylk8VQNdxMQinx
Bnv/5qNz53tHQy8nt7S0NjMwCOPSFElZ/7sh2voH9GeBjleJA0bR4wHrIyz63oowuYXaeXVLgam/
GAQjQ3PcSL3g1WhPoknQviAzsb3QHMlKobcpJ92D/tCA/VzSnzgzca0r4YisulJqTN38JSVPHant
QBqt251Pw4wx76ilGIgd0/dKoAh+V42m9MUQn1YVnBVaDdsLmpNf0IQxr4kviHExcOv14sbyGMSu
64wwEIR6VdrTW1vyPP4IrV+sfTGjRg8L0R2CE10tURd/3EDoxZDdtxme04ElcW2Nr2TZk56IiY4k
HxCQRYwn0n4X64MMCU8vEotkUikF5Yq1BzPbFVWXk3gvNmwB5j7lRoEv3iArj56uXL7/6K4FTkEu
vHnuL58oTdif4GmtiLdQ3WwN++NOLnLFoxAAQLfDilUf4leUfNqhFIuXs2JrLsWiwjdzbETC/3g+
pXXyF2xoStaGgbxG3C+osUMKtczENsR3qbeJ17pZumj0omaaHZgU5EJLkMQRjcP1hEQ9Fnxxae/9
/mGAxzszojALWna2FE1Ba+ny9ZIICmwPTGsnXEaDrNXOM5ErJYEjL0mKFNDdDQ40HTa1vmO1ZqJ1
YryBAcVuHNZISAfsT1bhNKvtagKy1HUmz2gCu0MkFJE1VObIS7Ubd/or8JUuswYUbGy7WhfXGZM6
dM7Jzyz3GIqVzxQDU08xaD9WAObq1PXbvp7Iay90Wsqrb0vSlmu3Jtj3UYYnCAfdiuvenYHQgEmK
iHSnxGlMXTvOEdyci9YUErFrsh3aZ27V8xLfiJD1p0RiVJ/jfNzD5GsxVQxTUbujCDJDgU7urBmP
BlVZb9YnInGvcvTf+rdkPdynHaUFfXmIAP1BDUXUJq/LESL/Oemn45peJkqI8u+1UIqiKRogGBml
xycNYwLDZIEJxtg6757X8y62vPzni90ibX0UxE16GdmB1G3ainhRsaXdImbLngeiqg9QRqk9kxXN
6rY4B51NWdS5GGk3ANpTmCpXbUAvO1alFUYOLbVKvbAIRVfOyQGwaoS4sJTpbusq/NSl+oSu31YA
+yRRd487YQDlOsKJVHTvvs6m5zzl+UjI6CSWoGN/Hzr0hZfs1XXqCymMUhuxyFPJXAOycTjFYOrD
POUmS80dFaemjC96vEKZ/4GEiK51O/CZGvKVB65RQL020pL5FLSfInyL4Ix7yhVMXxhwhj8OcKuI
ncgsKnyTSS2IJL5OqEHP4QNVsnh/AJLEPgWCdwnVmqR1eclo+6JRR1cOHJgzRb8fX7gIpzl/zRBw
Su/fFaQ+6W3YPmm77EcoGP3RoQqg7n4fLEwhl0usfNfPAaXAJWY+b3x4Jc6JMBYmiFV7AX1eTVCl
svurBzaSBBTb6Uz7mkc1TzHRaIy85b7n0lG56NC9t1NiGWQhw/qUgxgQvK4HLODP2fHF5mcBhW8D
43mR/cBsHH9AX5D+TxaPRbqlIWSO1yN3CBa1t8nA/lKkWeMcPHJSgImL4sSnwbx0/F+SCpkKTTjl
r+aDC3+cW1Fzk+QNngu/oHZYUjubke12gtli4BTY4dE/HFvtz9BAmC+ZLF85dRCNqJCTmWzm3ruH
VzjwPvpW/ge+o/VZQhgptDPMh32M5R0R8a/7npzBg/mqmAAndtA1zWroF0WRKXz8LeJw4K9BP0WM
tD1jkhZ0B+U2+9cvq5jdUCxKX8/SCM2F+KYPlNWBS2uXpgKS0TWpVrwJCrav8zTIsS7KzrslaHYQ
4pstuD98ZtK5E0XKZTRg1YoQltzmFdGzdulXofAYg6hpIoP7QUMyZoZvkI8NDus6CNw+bnKtucWa
CqZx8HoRsw3V3KhYOnbIVol9hxxa8+iqB/zg1NRYKgDFDoSOkrHhqO045jy77c+MlvnzX2dGkW+S
E2cTFQVJnU4qHCxsrBDj0mbp9tAXbVLVfaf9kdBqNMT/7NRIakZBqiAIozLRV10oeheHsERHPvvA
dluJsdvjDC/r4WyzGeDRr8Zs/1hYYvk3YORKBFbPSHg/eMxlOv3q+qjMEDEbrlIpJ3yo8rSMEEgU
P/triufTcpElxrrlfs+F92DuE/ge3SlIFAUMHN3xd/r0sTMAUCQM36+sbWxHqVoixMWB5nvkJ0YE
8wCyjN+k3l7+CyxCRr8x47QZoqFh1/XwET/Bh7zixDDWGVbulSXy0IhufB2RmuRb045MRH4Xlvx5
BoOTMr03bb9MHdXUGgN//If+Gy7OHpvvGSwArxIgHsKLNCEc1cNAMEoJ0qob4FWjdDnbAa1xx69l
Nl3LHZ6zEDFynye7/3H9/6DtKuLUEUoqOYCoUcx2ExMWhGfgmR8blKSzwOsLubpIbSoCtbJzRAkf
eSe18dk7LklAfB569OSY+oRH8XJ1EvXURMt9/DgqJ5sLPk3vxIGCblsGLwwQHgeI4gMABUCKIkvA
eRtleuz3f8uiJpcb93IK6oHvyreQRApyw4Ktw27aW3BIR4FOcIwcZUJ9czpI5Di0ZuL3j5z/k7M+
ndEInf/5Ug9PmlaEYrhYOWhO/34XluSG5hwg6u+8QhvR4WK6XVAXymi5qpRMDmIafntFd1ES9TjI
4DSpS1rmG8QVwrDfg6W5a+qCqwkgOa/dLVluc8aGXApluspD/z3lisWySiRYGp7lvlJXSl7MgFUx
vw10Fp03hCZSH60fFZV0+ocZbH7Gv29wQZMB/NevLGJL22/9LGIiQe7Wlfi3IN4VQ/MkXsYj8PCq
3wq/pzekstkWNCwpuO9xnEdywsvO8aj1sLNbyDj0S9LGZgCO9S9JokPt6eO5ztrC2tnUAXgLIm4D
q3tDU459B4KutqsTOgxJADRPTFPMeYXZ1oMoTMg9D36ehjJdpQpHSzZhl6Ic5HSbtrS+54xiIi5S
ZxK/STmgpfWJ9xQNW1+bzuwWOYgl/A43xtC5l4Sv4kk7CIgzFmG+d6kA4OeiMjRw0y+zLwI73oAx
HBI0cpEwQT8lqg8jswwjcE3yrKbvUOiE1SnptSy3cLs1eEQATqFOvHhKluIxRIYdzkihXSfXabvQ
DA27LvJd3xSO7rw4LgoQpcRPO8BFBiEs/96jOuHWtvsxGPLeB1SW/Ewnz02hOijOxNrqoV89HWPM
SWy5EoA0XcDEnXjKeWYWNrnbeNXTf2fk8ScElaAMJkn5fzKQ9W3G08aGy5gNXcLvbwsu34RvbuzT
0Uc48jMeWGeR0AnasIgzj3LTo9CCQ4RVGh0eHAlNBZUJBhwTUIE/QKjFrR+6YeoDXZvgt5iD3oJJ
h9+RuXxWWbMFmPVA04PEk7bz9LJ/FIbm9h7st8mlOon0i6ZMiQnHxhUKIkKZKghsisXPhLQr0KUm
3xhMvcrwBMG+2F916QXXdPGQvXkFeAH64LD0kd7jnaJHZXQhLQwTU83Rg8/V2QRk/fN4GQuYbcCW
gOfvWgALwgWtLUA88gYvQTVsdKSAPAc9MJHLHIs3nmZ704QYe1KJdNs2bJ1c1XW7B24dLA/AMObT
+HwlgiZWf0g23c6D689WTgdWr/nrlwxru6HolVzgoguyxwdlQBXjxQEg0jTsFBJ5/sjjl1zZVJEc
iEChufIR4T2SbjsyejJc1zX84AdFsxKlFvxOEopEt/6qhLgiG2DwSKENJa7Y+F96Ob5qo8ECnFn8
24PV9E49s9TYsu0Snzm+Y/IQ/Ab2Cg7tC1N6Yjcyx4jyoNe/f/2Drc5QL/Nn73eJqn9v3/jt5tMf
r1AtyG1+bDEZqqY9hzGsUvsJw+cx3579xBVWLIVBB7yZfOkZjwYaxrK2lkkJ0xrrs/YDHYi8OuZ+
WeAzK98yM0Qe26BC2cAThRrC1rRvGrWRsDN5hnOfbuFdmDrd0MhQRouEypS8budRvA7V5o2yczXR
eiR2mVxAQr/XNnSfaYhqAmuE1ul3RZFZy5TRkxSFtRyQqXrhqYvJuuKIsPUvHrTQZcCE0yffG530
Yzbmrp9RPNIWvHkuNY+Wn2g9r5DYdg2TdEmz0E5Fmq4oXhNlck8P20eeP52f6+lcY0z08u5nVQDy
vpW7UZIp0LzMLvSUW7VN/oyDKyQrv5Uh//1nyBgRbdlABYpRRr7LW7bu1azDq/jaoWZDAB9xdOZU
PUQKn6ahnJLEGr8jFyio8NzxmF9qAAFlovczuN3z9vvYP8eQh3d3LfhbAEryvtT4I5m58lENWmnu
4+7LpBiOh9MYPmVYp7E0it9OFbvXykz2UapmdM2oBG31jLOQm9nME724jAzoHrZfRfNRDr/jy/mt
5FhJyoy7iaaJBN2MEEUG63WaOHXJe6ZdvNvjJJpjL5eQiJRXGR/witMVH+LyoiS6HIvn8vEP+8hm
VQ3KoAO/J+9f+JJVLaGDHPvNm5AkO9giZzsFIydMBEGW7bnLg2FcfDoXl+WBLAVwFC5cD5mGCI59
px3gF4EMuqyXccvnTuRHacWSVAxxJS6lvBlauIy9yk2xtV8N+j/W2P6vYWQTqLfhr7GgBO1Yw3eZ
SPZkLZp3GfWuxRW7nK1Mt0RsRKViP76++h7XvTrRgi+LYil3/sIor05zxuxhMXkhAfBvgoSYY1Qy
ptmHrVSDCwNYFneKk9kHQW9MeoJf3lv+Id3FAqU0RFtvuAnwT+qLjPNBL+cTbGo+G/9Gs8hgv4sj
wxucnAqddoaFc06lK5yinbpJf236ylTOEwgS0MNpVSshPRb5ogMpT81dm6cFreJ5KY6sNQ8j+3Mr
ojHhcnRTqaiezs/o7VU7OQ46fTqVBgewfbc1GJB7+SZdZxA3ZDIDQWfvjjgbNQl14mbabOj5wRAv
raCDaZTHNt+WTrS2HXKbe22zqG6j+og6EFqrp0JpfmDLBirW5K+ySsfxKPefv5j/jYs3+J3V6H6f
aBn+ivoV5ep53IU0DAfUJtlGyIix/LVbQlFXjU/5Wdk2kkUruITywErHtN33WYPLllkse57vzbvL
jxvKLgugwQB15ROuDejwBMvO6UlVfp6QFZqKLThv840iHsC76pUy6XKz7abld+XfXHlwDW86fZzb
nyFOHgZiS6zMsSyqCyUSCH8Cvf6U0Egc8VyTg7SLqVF/Yqt+qRihlIXv3r9ssn1J4lJXuSq9+xp6
FRsnnHbIoYXLOKsGWKaZ3sXGs29Uvja+Oqu5NkeZ7rffSmLMHJhDO0DYRh7qAn2/fpERtC7MRSn0
jRUSxH9n0xrJpZJY7pli5U+Y/X7rKjgiU4Ei8W8O4+cgzpB2p+AHtBOe6/qYy+thzCnuot0YHhJy
MPnkTlDaru+tj1anEIJWSBQfVFjgYgAXkcMKMG76w4JTk8Wi7zFSd2AqBHJMO5Ssx+J77UXzl0E3
rIhqIMVIE+3s6oX53Mtxly94O8LYbrecTJiLvMUNI50vZc1//FIZuOfvzjPDXdvdr+DD8t1sZG9w
XCy2QXcx8C3OrZpGP95OCm8eofNjbxuqZXbyoF+0e0WemQjGBxn4GYfKhSPGpSq3Bcj9kCcBYDQQ
ah3ehczqb2ZOQVQ13wMpLh/AV/hMJFvbcYnJi67f5VyVDnFBW1mD5NME3rnm8/WheBmOPjCUWAH5
yfFxpfQ1s0HQZh6Bk6Q+Lp/zlbmAg56uPZ9Pc8bb1S4dR6LGDS8q5KoT2KLl9aUggsl5FOg/a5x+
whGZQ/3JD1EHUgPME4mOXsGT0LCxflxJvjJ+F6TUkmJIorW3J9wYq5wk0v+Gp3d6IS8QSrSUZifS
NnPMOibMyL36sXH/iDgZSfInE8149T0jLWXPl/RkryIJnnorCWYZmI6LzgaJvP9pRQfPx7rrAxin
pODm4BZgpHc95V3ltClmb/yAG/SuG5e4mKMZMz996/JQ8sPbFElWRJDlPwtG/6JvRhreRuRJzs7i
DipY6Q1T8gb2Rqn9qs5KrluS7vjpwTG7DaZE9N9YDXqpUVHIuuyqC0aXTwkCuawOlhGHkziSR22v
y5NZ6B1frWVpUFSqEHBNJGtmWGSqNgI3DgmE9PAeWc3nzsXIyZnFCCvGnvACwdJtXhpIlYhcFoV7
kpmw8mPR9cPXEJWS9C3GzSm4aVTEcC7EozFMNFxDJToKO5zibRvK+ZWQmGPuBv8fahOSoxydoctR
qtH6TIzdEIqqCxDlDiXYJ3SwA8m7Xfy3xL59djBS1WuzN5mb09muR45KLFk3KhUWH5GnZFIDpGoT
zI6C24jD9UA9u+bS9CrWT5RuH71wztK6JEb+FTuJ7/yNwx7JlTJVLifp/cpYl1phvpUZFKyrvu7N
Fn4quwvF0TIigS+Sa4lMtiCpc0cmr5d7oe+1BzfZd1D+o+B/68zZ6gcjoSFkD6AkTiwY56bl/0Bv
e9MrO8roaJ6jpmjZa5umflJnVl/i2cBaft+lntq8H/HzYhSbS/pHPZ/SAhf+WrpDhr5BrZ5xTqCz
evrWVSvjF49QEbP9KALs6YYWqe5RAk2xvkppqMJAo3xQvnp3USYi5xBXBDFskHyFUNabchhuN2z2
E8iEs0MioV+Apa/gVl5doct+LvxR9vFlLbu14HfOjNy8Wj0qJwfxA/q6BNCzG5cwV/yIjjGerbb8
1ybBZ1ZWY/cN/EiEdSu+SFe8uhs2IGrPxNK0GXYoN2bfBKzgfMO36gY0ln64lC7zJ8wcLyFk6R1c
eCjedmQSwySsTKdox/Sqm1lEDRcNynf85WDbL36j91FDlw0IRH7mwhhjQV86Ece3kqq53H8C9sSn
Zjz2bEyxBT6Hx5d13kizINp9yq+lZIkOi7Dd4MTPWNw0RIjMXrBnXUFZ6XTWcWD2T2aJrE/c0bGw
tO7EaJ/uk+R9XZ3uj5oLyqSu9QDVwnPSlHWFcWxujAsqBxwXMPHO7G6hdeRVFjCA+d0Qdgrs+rvO
NHK/leInoUypMsfiIyaGOzjwBH+mkTanxZ3b4+M7v35kvuwI7J+5DGhecQ0DFDTntP1jw4RDqfbv
EHEZHGKF0CQ3++SmvNAv3ku4fD3Z+sVFG5XULiWqgeo64SVCz5oKL25IXCw4dDG+qfcvaDVdpZGe
uf1/xSEVy0pUVeowdMkyohB/jzDUyrsknedX32P8x/91O3UqFqGvGFQhEu76QZwRqA/5Epz17k/K
2QOOgDgLtFloOR7iEwLGMtEnfGePrdOIaVmgUUSoGpLuGO0m7TQ5QLoCCQ6+30Cu5hMZLu6B1V7u
w1TVfYzHUAvZUdjM0jrUIgVz5yC0nFFZf9c0cGTPi7fijXTAuchU9OU1ng91dmhJ9KEFJ89NgiU3
gOvN/T+ZTyNEcPwpjigscMLe6rBGgUBHHGWA/PzAkVxN5fi5l/brNn/B9yfJ9hXhn3hK2kS9hi4S
ZMfw/GKOvOqYfKbYvAXY/HmW/lNY+actd7dXUTP1IYp7Ufb1xYBLYTcqxM6K12ZMwURW8wHqW2bY
AmtlmgJKZxsF+9/6svY+X53ndrYt/TE6bgEfvrbK9Q6eoKtGuI+lD4lHd0EpjymOeP+/WHsE4B4U
fNqVb6cJKruvIyKZknEnWKsFrI+dk6WY5UjG29KtlT9rW3q+Fshxnjr61jcjxUOzzX/pyE8MIW3Y
4V8LuoL+2WKTw0XnbMNbr1Gaa4hW5T93wLd0qCjhRt8Eu+WyAAQ7Y8QC/LjkCGO3o7BfRZE/JG2s
1Hug0Ao8ZrCl7o90SE/SZ1rWnlnD/ZNFGXTpmUzN7Ye65ohkmedzZaYBQ0UZSxS+ebeZHo/mHHw0
dApwaNdWhJcZnYa4wCBqYEJ0peooBW3ZID0rtOhSESPfSjJb3NlXhBOvCHwHczCo4DiiT37dMlg2
s1gu4AfQdy0a0jTkFHOkUX2H7BfqftRsKOGR+zCJ6iEIv3krYnGRj5QHHW22ORifqFwYz5J/+k2/
XlQPRMk9quFfDKPz/vhEPynj36St4EOp+tnCJ+GKuOqnqxm63jWcBflGTUfZVaO0S6v3D0qaxSRe
fjs/+WKHUQ8rEaZNBDoW3oMBqtaTbKMT4DivCKDfhK3CJ8/eAPCR1iM8GOh5FfY/8JYIm2K0Kyy/
sSHxICxQ0ReD+BomSLz/kVZrlQqauA1I2aJ9Uaenk44Bj9Y1jTxdggvNKMkY155CDgzYE9Y0qq/c
q5ZIzzP1F1lZNOcATOoGw6EalWjMx9k8m9CJy765qMflNduCUL2cIpLBPdZ+oDQyYNIVCpOVq05N
QAoK6iGzBklT0dOdSXvOAMVgV03dRADZwlDfraIN7FLrwDQkm4o/C1B9Dzss7OgDZQfGXVI+POAd
g5IKYR5v8OVSUrjTbSsAd/Gxv6kTEYMxKIVACl7qfn9p0FVxTW02xWnTErSDJ2OrWEL7dXainwIt
9cWIVcT+DUE5HHi5fkNxZDMwoCNY+OGNTag2J65ze6ZSWRycbdwu/RbnXcCIVRxHwIidEGJz/Xrq
ysu9gqeDEJHN/CnKVzYp65C8ZhshJAH19ON1337rEPi12/axQMBaGzgbUOHmAxrxdCFGNGTK3WcC
yQ63PVZrFoJn4SV/5T3nDOfzEbXqFYU6hbFvM1eDkMpbvwqgG9OOy9s5T6/1ohMwHgOg3KEkSJ9n
8UZ8x9Z3uIoeg+0Eu3ZRdU5B7GSIUTDRWgqPdPTPuosAx77sQcZcmwcm00+vUmVTCmJsu2jL3BZH
5dyL389refSCT52/mhQwamXePr7htBdwIlXrtLYY9o8NPG7yKJeB2m07+L5eKU6vpRx/Igc0zMIW
cdKC4jqeySVi20HqtHJzoUyat7Q6iBBnzdU3rmvt9KE/8jPXxuS3mpPu1IZEcjhWGUyLZ6V1c2On
+t2QGGem7K5yNzr9H3OceHlRJyH5GC2V4WuqQ9f99oSkRL2srh8RweJ3feGElDi2/0nyILOVHOh8
XmUkYcQiXrdVnDC2Tj8I/Ci5yB+dATaYGtFTT2eEkdu+/GurJcYA52wapuR/RFUR0Se0nGAtMmhN
sVhslmWxBySeT3ADgLLt05VhrNQ0NSleseIdyPwfxyvylmyvAEOzJzMKY7xghxmfblRHuV/KeJG6
f05QH/3lHztkS71nUy4HgkvhwsugSbBqXMK6kUrraGBwsdOveuLp/6Lck9NFH4B/c+RP+9O9pyOH
h+267MgdBM0b8wJNEsDh4c/emC92oOHex5GzgK0DOQLLLG+UcJzAxh0wKz0Ur43E5j4i5sDPLCrt
2DwYhgOGhT/8/ufcLUmS+dXFTn5FK63mTaQXmf/jnGwxz9GXwac77Jm1Fvu/mAnevZeIUi2rId0/
MshJIDmSduvc+bkFwvKH1zPVgTt/WGoqFXD9k0QWOblPHq5KrhcxXcjf6AMxQ+Eem0A924KOLKAr
ixZj0t0V80egHRJWCJRCJJexvSJo/tRp+slR6dWvvRgQRmGxpLjatp89Zoc2mFdhra1A1QCA3v4M
FLYyrHcZalqx5kpOUSlvowp6W4UvqJZvIcwcc4lrD9Mj88aBx2ervwCdl0MPKVPQaF6zmpbQt9uY
QMnJDOEjtuXa9Kv1bpN98jh/LWIhg4KhUvoEmt8Mk867xprDaG/2gNnhXjOhn2WGujDPbjNdlvcz
MCqVSuBVgdn/mDAz9N0TIzxJT+Dg75APMGrs8+2DHR5Okt0Fgvo58LTPDEiNmqv6cL0JpkNMp6y2
RHyR6r+Zm/lP3l3/PfLgKeoK1t9yWDq+t/p4SlcAdEvM1UkW9wU4TbnDQYjWyUclgoY91iKZ2BzR
QX2awe3gm4G7X3xOZSz50qYIYfgkyCIAXlnKNH7wqL0CBwSXtfOA/rnBkPf4lhlBMTsF+IluQwun
Vh7glwQmLRGFysY+2v7ujDPaRnMk6sC1GEgIRi5Qw1OfzZTXCcIf7HyvaWMJNZh0V7UemNZ6MSH7
ZhlX7aErpvK87rYT0gDEiBXFQUqJl6l3BzKILj/R2Eg8gr88L2G2jF9wDyuLMjxRSaYKSZooOqrA
PFMQw6mROo6tuvAEbt5qtLB1tz/3zNG7ZXy5SdQ7SkAkd/yqUZrKaE87+oOeB94jFTMOzkLcN0p5
FJ6j7dTn5NtmyZynwQY7RchHBpKoaCcF2azrGp33qUhnEYbxJixrrDr/ugHh9ithHgjGqRcgrw5C
fcCLjsnkx/lPB80y0qGi+tvKQAnrcpkcVW+u1D6xz/lq7X6xN5SE2WtXd/5Cuv04OddslRHvRz96
hGz5xemkMtleSvpbde69VmSDka4/Xe9YpMfGr0sEaQ29vguy7h6T8kzXjrrd5xQX5XDqu4IYxnQW
tvQ7zMMPuXHYDLTYB4nSmrhL59cR8M+10vPAaG24LNcfVlNxKxAq/yvcJSu4UiW2cEE4z1gKts68
aQqJYjJ0vrzTKzXODNK1Fjt14UbdUQ3BknqSRXKS7MhQwMk+z/3M258PZF8xCLSZz8td/T/CzNaQ
+p+vcTk7YUEfls/ChEZPNgOju71TOZDfg4+msHnfc0hKghlj0YAgicF+BDjh1cT7vVcSuXfwHDQf
1AxQZlfEHUlYPjJZoZZDpFIjQw3HwE/cQ+eKTi2e4RIVzGCEob4bKk7hdYMhCuO/xSpQGya4vfg6
AEVL/V+yx73+JlusIs4a/RuhCxZo7Wm3nMqosfJdU/3Hncug6ccbBVruditEOosp6dYon7zhDe2N
AIaQ77DImGinYZ5LjnTa0WsbkopNvW3z0jRgA9a0u6KyDueqpZeGIp+ozT2A+hHQgnjAEEhQTZ2O
oYSMyaPfW+zmxLhl45aVss2YzIK5iIyZqNy1Eq9gV5yBnnA11icVwRshEXz8/UV0mYyD5I1LESvp
caXXGFLW+SmHMlsfAudqnIHv886u7BKXQqnBJEaFL40NsfjWhubwa4CmRuN5aD90eb29DA03VDmI
Isms6cUuwaKbGjAShAmCWUm/PQYse3GSiVZ4z/e3pv16l4OsdjybwHAGRnHEjdJJLkYF0UqR8SBQ
9C2ayaLvSpcbUeOkFzMU9ZkvDQvqhQDx4c89jYWmT15vfWpIPTNNJiVpsV3annZCMKcoI9RfrxId
IQND51ignJ68vV4l5s9c+uVaUTbai2tM61TeUWN9RDnqlwhoyzzPJfcd9tED1tlkUht5f9E6QYBj
MjHGrEjf8vbhSFKTFsiHEdI6Ge9rbdM4Hm1tAuvje9kVB+6LOuJ3hFiDBIMc/3gUVlMtj0rBuKz7
H0dwmTZrK2ZWSOsTb3+pIx47+MFPrNY9kgmxbCbKoBtXPHPh9nQzDPWS6mmP0dARC+zAbQuYDG5M
lIA764TMwGtmigqj0OeAdORF1DQ25BmT4v04BKqdKVpGvfUv87g1VOwatQRuX0vNOlKT3RvgixwU
cj92V7WbdsMFL2Z+wzSwlXT63UgVGvfXoqPBSHWNFktgWoOIItShFIbNgfUxuh7xDWDkMvagKb2A
M6afvBTtZ+Az2EOQhedeyNbrwQRjtTopo1hn7Clwaeh2V+KPslGlbpeUJRNiC7tdmBT29kszS8IY
CGQ+YYYCdC30ks5LQZYhwSx1oFwOXEWsCtd2J4nhvQIZNgluwnyg+5wUR+BhNaWjBHHIA/rDrA6E
SEO9wQujk5yZglFYfJAmr6+ocCUk7UCg0mrBsYcWNwpF4P6WLaZThdHip3+jTjpDS7gS+4yIUCQE
uHCAKq5zga0IhIiSNB0AxunW24qYewJD8LfoVgzxOZPmENsbrritN8uRHlQX7AiGDnyGSK3bybI9
ibIVJzk+16U2s7IRRpZU36CQskzEw0G/7eAKKVVIYP4rnTyw71SlASmCkdjnNvMC74TxIaCbAHzj
DnOtJwbyBRT2l8O4xIP0Mt8b230YdUqvrDmolROEeJgXDjAgOrxVGIrusLbeMpanV/SeiipVXgsv
SqHvp3t/AWwM1hxgmDiXeXZdWLrRsl1LwPRQMh5fs4QRxF6+Nvuw6AsfUIbZcDPIS0S7QWzwBXc/
J6kHSxEqxQ8wjoMbugwzwJ4NgXZf8SQiBFs5FQVYDR3rL+BO0rQeJDA1DPi0YW9kAG7LzKHHB3Nn
5H0KPSLJGiZStvsgwnyFeSz3GjQls+DamdFW0Eo8LfvRWPn1AOxPZmz/ER3JMEei5Ze2Y1PF6O15
lXu9p7C9h9U05x+/8QfipM90QTRMZqNwlBhKsbDaq1dxerVz+MzTaTw9vLuS2QbW0jRG/rndcpv6
yHfAGAz3Ep+bNvz8e3B95fSX/XnpT6CSQUfeuKBLf6XgMmHrLfHJXUswMoJP/tSixrM7cnqMBSnZ
9Ik6jxqVi6cZQyDVY707wZUeY7vmkANIvGdej5tDa/xjMnnNKGrlVDoZt0mTyMUbeiF+aRNDKdnn
b5LJeNr/vmwnrjLQcTUGwt56BihTr03lAflxtXcxRfTlSxZrsaV753RcSv5W+7N4F88zR+5gahHu
zPJqTvWI03J/G6yoNMUI0uFYYnV8e2iqi3PW1Tjbapc0E03cyF2jleQvw2q8SKpw/GsBCIrKn4ev
MUh+N4Wouu0w0sYHzxEwLcRzyzKaJzLnDQgseNwZLT3CtWh9t2puqUkUa+t+y6TlX8EkM+SN5OuD
iFCoEy0ccO2tONrcmdbiTz9lNJQABZWZF9ssCvja5xS8GH2nrudTg4L7ZXrqCQ0pZ6NQfQRimJop
Ov3yOrf30DE3FGSzcZIF6AAvWvnMRRm9kpQ3J9IVlvOOJPk8soQuKgVTbLlaQEeZdOUtcZWp1Pbf
q1kCx1EUVh9O+ufSYt8HqZ93shOo/7nxVsdx6nBcHlFYpH8aC7vATzYEOOwS1y+LhymMNT6pvGYf
ERQgkETYS+u1+JpNoZkGCk8nBJIOqZlnAA9VVnTDXLi/xnXMm8YkmvqSjGfWriKFOkPGFZX65Xxg
y19iTtBE+uKvS83Y2sUG/u5txlUs17N4Az81ijEcTeblGQXyDbAGFdaYnGvjExWVXohtENN6N4TP
8uNQ4eG3qJnP74zteWSQvhcDE3bOkjXDYUp/4fonL/yfD3w+j5fqlQI2GCiny5ipMSYf+SeButie
bQyAUSTa+QnP8bzglcxkGHLALSPDvVXs8kRfjlA491wtA5ol326Ry1dcRU2CiVHHJ3sdgqEXPdBd
1kiGzvLgM4mDcMl4XfFphOAOJ29qsQTCXmu3JVAWWbWpe70y6OfVZyl5jH+/7WJYCTq76N20Kzzb
f7YEIYonBQXs4eLv92X5GrSLLXEhktMSuX8TyLrEepiNUi1p7/VHDuwk80ujdfkQTlYvUJU0C/TJ
+tp50FjDf6F1WKQcT2oyCagqqD4hwh7HIUtcP8L1+rTZrJWHSVYUOdNywCZKDriou+EgGrPVWVby
RZ4IPNKwCoePbhBa2awCgdsj3RIAW+Bcru8XfeJZLiu1PtWz8P8X5hZ90u1ToKXRYmdYgYP05eXn
lKDzePWcJIUbL+HFxt9dTmiDZXN2XDJIMBDYTlTMgcIiIg/WtK6Qkx6axzVX7kGl8c8N/B3fCjmh
Tsr1YTa22y/isCa/UbC3g4/rV8g6kJdq89bQq+UU2bne4m/0/Qp34FXGU8ga42JRYSvlRzXs
`pragma protect end_protected
