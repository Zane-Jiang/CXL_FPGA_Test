// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
O5xvDDyTGrnu6YH3Ea3zwvtCpRazQO4wCaJyElfx5BG6/rna0jn7a/F77KfyzpSP
7M7M8rEyjmarPZvdu8jUMJto2lpKZ0EIbpDy41QtKpd58H5nFAuWMzlor7vSNW8W
SyUVGOU9VnbHhXOzPpCBSt9+ol7q/74qgq1Gl/hKhgw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
K6qHM35kLf/0QzbRPUid8TE8L/NUVe46AAsTWcwhHkPgZhln+UX/EkyUl0EnNrIA
a7ToWMwh8+/p6zwvAXl2YCRbT1rcTUFVX/IrX8Hf1Zx9oVA7stMF3TD5zJDePL/r
8niZqo2ciCqC1MRJzg7Yd5DclI5dozQR0oZ9YHSXCkYL2v6Hl7hwTv5F/jG5Q35/
FtjYp+S/3MEDXHJF7BRl013e06ka3pCXLLQjvHWt4tyGlee/3ELK0793xOPSYXBZ
nxwNmhCX1nPMQ2Ttoh4sZ36xhQCdrkcyh9x8QPauNH0OZ5jprElTIUiQOyk6ZdVc
nQL0+wLNb2x3fMkpcYYzSM5Qfvkpg4trzj8nqyLWFIzPkjATpseT2Xwua0/Selk2
LAhtg/MKdixVyWeBK7hX8IqjNckru4KaLvu/bqttGWLh/T5TyAKp5s44/wb11b9s
SkAjnYlX5fvstgIfNB4CJfR9nzTjfS/+MbzS+sNEhfNMVuTyiGX8ddDttzvKiBmf
zIB2E3et3wzzKel2qyEBzFDKezDdHWhsNFvIHQ2LcZ9QGdF644Sr06DocsZelUy5
mxqhwIDZvfdwprJSDb1K3yX6GkGLt5WNTV88vtZXfvyG0XsXRGOzrZoA6qa8xcGi
MS4lOLWbAO49sKH6tclmgijdVi+vyNQBAsJe/LUiWmlIrpYifxCooKvv6yNThhVz
jpV0VYAkl71Cr/s621FhbHXwrWpAc+cesg3sb4fkusQsekWqxxThgU4R8jTcoYuj
ldBhNd1w2sbIWqARPX82LadbPZGsASZYxIAOrEbEcfnBB64AJzcdyVgfR/g9STIP
4woLe4DB2YlEJwNUp+dETvFl/el7+FbqwcQF+3J4NbeElJ6FI+D+AgQmtOuFDx4K
+bnaKh/n2d7IDa7Hi9vZPkgzSSJtk4bRwgCkf/ImfhQ8Dlwv+nWwrvJWCN1e8Hir
zYwRbvDYnimQnGVmq9H5lLN7DvGh3kqVv6hYtcZgZ2O6vyt4rb2qJXK8wPw5YIxv
8NkPGh7qWlilfprc2Xwzkttt/kKENtcTiKiMmBPd4whd4q9I5RxMbsdXAUTZhg2O
++O8CPmobGQcYzlCbbIWsNWsVCyj1smA0BUUT3gFwV4X/wft/Q78RnPZLIHirQnH
NmtVTQbLJYHe8nsAg1X6Y/v1kaq3IyFkGIyqa1K6/9oO8vRZYvZgf9xBkotZjK4E
zp0A3zZrCm6eqZAVEIJrwModWkLwtfEHhTWltnp3QMPpTCjfnJoCpy6nZMIqUjBy
4Qrs1QV0B2duFYISq+2O2ZLvvswzdC8/Lg+yBpfCrHA4oWF3K/YNasMyF7ePxKQ+
9jrpTIjQ6qSuGmQtlI5GQn6+NpGQj4r6roBFhR2GQIJduVlOB4L4detbBySx01be
VujmWT7/ddICD86V7hIx5SkZKtgEMUorCBfaIMFfkmEc2P+6XFwyySGM9vhT7Vi1
IO/KpiuvzuvTmJrZzHS32sGYmC1RT2cw0DzTTq6O8gaknvYjvkUwYO75/9Obevvl
rB3Bs1jXX1QmHPxWb2dQkXcZKpgcRXKM4V6aShmColELRvm3eklk5ccRyGRP/7Xg
MFbciXZFULbVJ6yLxbPlAK8DtfR2UgXjlI9FPTawS+sZZxSsSLCwtL1w+MSsMo8J
X8L9rjHaoDiVgSA1LqMGGEf1t4EPSoex5ccTKwQLI9LTIti31owcm5bMxwXs2I+K
FkhRtdjJp1MPLopQlqBFHA/W9LFGDrhkBCZNscS2EdYaVM7ZoyE/+aw8Aytdve4G
nPe8ZiXJD73AFHf2UImdweXSCh1TtVWJnIGA7tuWG6BMtJ3QQdLHHXit/hsSL2QQ
AivwAdaMTmGsgP/iv84QoQdyPI/HXSo5dpUUu/NXv9mfznEQWd3q3CD3el854D8I
PiOhYcDWQOo/V1D/yXcHlihs48PuDWgZJRtg7ON9S3hNmTBS/El8TtHcM8VIcyn0
cl8X0IodanpuYvv2iSf8xSVBMbh5bltPZF+RlkPzl3Cc8/LxE4cyjcCh85xITQFW
fGTXO6IdW5mY8rcOzx+8xK9HuzobBf7EvJAEqF4fENqvGwExOxGWQk4HPtBR+UIg
grg8gZvFKIByHH6oFiz3WIWn8MjSh2/bftYKvBj1wjuSo7GbQOtHjk+q4HUFrhGf
wVZ+hS7abT5mwNtRVb1O3aaZ273NXHEyhsdhHusPlR2VmtZDcYPnVC4k26Grqisb
gnFhaKLJOfvAiMjYFRvmicHmCYqa7LB7WCy2dCUXxD4/cFJ8pHH72bQUCt1FBSQy
06pbKpaCJ0JG8LvmdnsZM43U/3LCAuovBxaTUXka4OPztibvoUSm4N/pN1pSIcHb
FL8xHkgO1lFQKkaJE1YUgEp51ZhUwtOQDYZ3rBtm6Me7v4SbMDObEFx7cuHh8kR0
atBUtfqacQQJA2uSix7mirV5sl7QsHlcdDa8EvH84193NK27Yhj6PzvGVnlEj8tb
fzTFcZ2FU8uXo43jqx8weo2EF8mzpgFSfOtnZ+mbgDXs1R7Rprx7OQfksWLZ8Qjg
R3r7g34yGJ4eBFCLTiz4lBFNxXF7hG5YP+BKOMXWtzz0nQohQkznuVL0E0/rT6HA
yWZPXMWp8z9UiLpSnAf3ewbTXdbRCYqLyiKqwEWlM72pR0Xdwhxnli3IZqSLph0B
4I7bCi0CHqbjfp10/329PDYhcPBNjtpSTikq9O+1cYotriTQDbbw/6uBkrvPw9DC
kNiY07SFFXMAl/59qHdolucdECHz35ie/PrexAvQPd292WNxnk+AOcz9qXHuQ3AS
tLboQdmMgOcJJRX2l9Xsf5sHdDHeDBqosOhD96AHJJHHkvHCJ9dSNl0iCpnuamYZ
m7Tw8j6e0vHvVL8Ai96/d47bcOHkl1SNn9ZlkaQAfjhZkvYSLQBp99t5/gEvl7t9
Ge+rIZ66Q08xingEJZKmx4vgGaoED6WjikNCsbKUtc7h4H8SqAgOTBzWX1YhbiKG
iF2E6BeIlBPiwRSuuLmppSWJp1HUgci0BDX9yFqilvRWc23UDP6yn5qZdaxxG5ht
T7jZUUnRfKyWifmJVR8jFdWgd2DBi8L2m1wyLrhIZLG9hSH5GzGucJEKA4f5suw9
meSc93UGC+NmCw5vu+BIPMOa6QzITsZL0EofVpZwWOz9BF+6FSYGWIO1jKQfMQlS
E3TkYX6eXDwr/r3uHmUL912Jnv8+Xin4MQP2sh0KFRkODXyUXj3rW4I2dT4ONqaF
Ln0QQlV5yxO7dF5c+jCWJzKnVEcBApVRR5W4GRRi/cdZaK7tdABO4tAmf70BNDzd
9H47TV4pwPt7DD+FwlcvdZdLWBairJxBafqf9l6ka6K2Y2obdR66/k1EMJIi+cMD
NvQeS9GBnWRrK54iC7MxQhWmdLIX0wIbucrjkEkJViUihNq8a3NIymAsrDqx1iQg
yETF0sbd/9adVBcM5VJlcWXzgru8hTHg7XZ1BIOs2YBObek1EzHCemaLclthTWwe
TURa25++Oh7p1TWgrOzuaWBisfUtJ5/4wO1ULwU/N6At3iMOYdLygKIKsgx/Z+SM
L/Z0X8nYm6HXET8Wa/9CW+Ld+eumX2FCCoTS+RG5SJxIv93vXHpJ1wxcF+QDcpjV
S8PHttn2kOu9Q1whopiNivTvB+fQEzbA+okVn2H2URibgUA6Wj1N0qehSDZv7Gia
P9Q/9E5X7rJ64T5FC1ioPRGwED29CRCVrKpgs1hP6qPf/gPWQlO6vYvjR71XVY9T
Y9GzbOZ/98N7raoSbJiRmzWnM0MEb3oKwdHcwn6upf4WUUgbJvINyQQb5lZTTLCq
M4Csk4r/61GA4vikJTTkpdPxO6rQxnm0mMq4s3LCemPMTF0pA4Naw0zEfVvzGxkJ
t9YfimtEjRD4YSAqgdidPB4x0X+9TzGhkQvCqA8DFCINmCUMv96KGdjQdnZFDhjV
R3jRycg/QXJieOkSWz4+PJQklDSW60q6VOHMkVBjn+ku3nPtp2qlGFWTsTEK7WMZ
FTDeVXuMm5IZGyM/mXxrxxgj5dxCTc+1bKRLcU+DDhfMvSsRf/tgykueZnrp0j9E
TEJhm9v/nwKxL1do+4PMhxVRO/Kln33spL0AQeeeyTSuAzp2mDtou2bDAsukY9KL
7pIP5zPRUo6pVV0JSeBN9aXlC/CPrBGOSkcwCImppYIHC/P2ZQxwWunhPyeWcJPk
WO48fAIUde/frXJETT/X9mHddzFYj+UVnXXefJTzhGKeiLJFFi3uyZWbzxlnEPQR
kJbKCDwiQKqGKnOZHQkm6R88fqhUYJdU3ex5zDJ2HU9/5myKqiYwFAmYqya3GRup
ZSjDeTUfhrqOYU5OWYQql2zqUrL/tlSTrs4MZHpz5s5rbRMDrSo8MaNxUfz5bQWN
O4c9ve+TBNgUk/CCIZFANnRp37zN+t/QMuUsxe8nwBM08hdebjyD3jHS38HIzk5D
xf+ZwA/MGe43f+i1agEt3DBa2Cmcon88gdbDhSpp7Rj+z/p71AF/IWY2LwjQxwIq
VAdCNHKV7b/yYuhfkNEkqIzBigKta0ZFHU+CPMqblW7HAFy6wvgGqizCKasgbTYq
nRQi15ILyboWkh0ci99MHkIxUVQ7VwiJlVC62sum71l6/ZhvGm5MQOeMkNEA15Ua
AdhOAQuvnTJHMVbP96wkpOtphPZ0nDyLtJyT5u9UfmM1YHeBwjTimEOKBbZsFjyq
imv+gRsAlopvNKxa8dMLoS9RAECtlyCx7/eMvcwjXoLA+mOGIZDE/Uzx1XppvWGa
FdWO4njqP0P7kEnLVQcav8nCHUQkhIKiOrwMvi6nV9Tl9MLQynTkUjSoRjKYElgm
fLC7gxwamUNXYsfnzMHU9nerXb89MfPEsLwlfV7kyVxXTMIgUYOmOUCzODQ383Hb
jRxf51khUCkfH2uQWEmYKgODE8+hG+S67nZcabjVxmEKE6foEpRUn922YKsQuMWp
nYq7bog4mD6vz/cj/Bvbqw9m9IlNImFZ+S/Dl7zLiwQNZf6vY68zlfeiUQMyS6s/
jca4ePbdren4i+JUhY2ipbiFvNTfCVkiJutlCt5JOjCLDiSDuwgnMrvczI+URPD+
4K8dczL17lqIqv+UPljjkQNOBRFMoMqw2DTH8Vnjry88L77G2q3Kw66iWKRAusfa
bkBQL7iTgpNOrMua7x1OZdqUWrWlMjxkG1N1aEevYyFDr0EbBh3qfOHhEiBtiXcW
l38AOPAJUWUN7pxm3HA9Mslvk6ZR0l4/J4JHOw4UP8WP+x84irJYDtX9RP7G+yiu
07ByzDmAFrHJBYZv1JXtjkEv61dl1obYs6Sq/gPazbVZkUL0/Yh0kpPwskuhpCiH
fu51ORYCxUmecwR/vbqDA3qEJ5t6EpiUS39RyJzYGVamX0scL/wC/VrhtrRphHSJ
MbOksxckmBY8AO6PZB+c/TeOCq3Jy0iGyZrUS5ElUQMyP4zfxRwYD6fInFmzRmvC
bNmXAK/7gzszV9Mt5lgxo1rX4IX6Fpj4zhqHYycgwjZP4GsF0Ej+GeKPr2vOQaJz
ydDjiUj8l0t8GaodJSBzHjD3FB57nsF93EGvtPpWH4QRN+oYgJ5qdqI8Ik1cx5uk
rNfd79so4pgZLCejXVXBY7njDn3N0R8ji7x/qSJOXKE6Ks+wL+hNe/yoT2GoG6jR
d75e9+FPUa3hwXhY4tA8yU3OHqaiT177bo93QZzrIUJrhdgoqWLZ1hso0xubO/LN
uQHGHhk1CXYp0TF4FcqBXmkYbe98TQ59Gc0ImkJTbIw+OFmtc+3LdHxVM2QEDTKv
PzcywSw5R1b26BoReAHKgy8UaueVfiHnZIAW3Ovka6hLxpKnmgSzJeAHxHQCvCZT
4Mwh2+e3Ng1/jBw3J/oHMwLmd9/ucVJZP4WDa5yJhT21qV3tqxDqbYfQppFZ38ou
zMJ/ggNztly0GMtsZIsn0jkPh/ug4yEqwbS5XNlQhwnNWnuJakUtXaPegS5Tj5/A
gn26OMDAR9x/Z3lJ/JI7W13EMFi6YH62lIvfKH8NfkZ1RDlUyCrGJCQp1VOMH/6x
yTt0wXyiYr8FVQoKuvwIxjHPBvLe9bttj8/W8kYqskICf8cfkjFZLG2wkOVM/x/j
EX66tkDPCoryDZNqt5FuaycTXOXsZWO4mChxKSEso6u112y0Hogu7vjHfnLMhwME
loqsKGwGc/X0CxuyggbEJALKfs2yUlbjI1I3UKWHydOonuyg2UFghe/zw7ow0KIf
atEsLJsL848LVGJn1Fd270ZG6hPkOJy/tRCz8d1u4ZSk6NJ9uL+c9ufCoCobyRKw
Tkp0m1hdRo6W0mHfkN2wluT85FCbg2nSlhx2uXmr7F7uudYBgKYu3aAS5z0xPx9b
2L/aYbhfjyj/7Rtan3JkdsNvAuPlnvN3R4PecvwNHp3+rlWUYLs745d3oajbt3V3
4UtftehacZi0AAsPq8wNV/TrB87/BzaOr9iBLsg7eUF+Yh7q2N5sKroFhjKF3DPR
bN67zeQeKfr81y3aQP4N7NZwKdP3kcDRL6xoPQ1nAiWZ11+Nnz4rMapOIFacivo2
ZhAWUZPTGrHaFFkHpu/FarnsWv4Fm2cU+RpCahCtGld4q2wCH5/YQw3E6k6wzKrl
+BWz/ARx61x52ahlRPvttzK3WnCrZn9GmZf7Pkm/G7oncvUYDN/MhesDei0bAa99
ysp1R+LockRjqmbM6KVsBypMkfBA3+ceik5VDoSKmJ0FHGduTPsHKvJp67aeQms8
niK3JXX7bn5e8z11voABgb3U8pl/HMzei7Oe1vjM+vHub0QZDhU7MW+0d5mP0dv6
qwJLSZOQOA3J7HcKRKNCVfNsuy2vJivAp1ZKJNrOGMwCT8AWnJdcNlCNJnvJ08Tg
Pq/ft/3VGgfngIChF8EVlNxAgyJZWZ4KnxPOc0k64ra2Laq9miyfB8+stZT8xuur
y/e4G10e32tZDAZ9rKr/61vfmLCUMHSEvSJLxOXnRtL+jxEHGD2dIN52g+RwbRgP
lMymcLr6OsyBtDLfDmCZ/uIdeoP4ge1MrrTk5y1J6hdbH5zZA8USpWoR+elTIGBS
C7CdxBozeea0m88wgTT/M/ut2lnsaETVlhfI2Zp6HZUWketCKXdMXBRmlDuHnKUU
7jr1DK7amoxkPMf4dIktoGLtF7TMCy9Cx/NV/9Ju3lbgbA3G0ctSXj7wXCHJHvXS
TUmpyBjEyZ/2x5ZpYPPuhRMycFU39q8+zu1EG7lHG5Ex7JbgAkMbmuYw7dXpJDrX
zjSVEhdF2ykrPGIDMx7DpbPymG4x58VA6mSjg8mzPWasnhB4b/LxmDSErgC6oBSt
kCXDzvFGByTzbulDkpKkMDMcd2Yjh2ZyPUi3ILeL1pOA2QfGgUJwRMtwXD4T2J0B
OELYpR20pe8gGXff7EL3QvtwfFb42DtCgBbucesEnbjYyywL+iaNhdOBvhXI9Z/I
jDLM6ax5/D90eXbPi2ieyduG1Z8XUfAVquQkATHSydTF0yTXVqzioq2etre03QiN
WvvTTptQeFtlP08Wj9d1nRH0NdpusdthSvXRMnGrrgZk6tNnubdZs97SLsVHMlf5
zb6YlZdHrh212nRrjQ5k+i8d7Y9FKSCYBwSp0tE7QGDdH2NXZOqmqqa3yoZxJIYQ
WXlFwlP5USCPjMWuf0FEyIGAj0KclVSzNuRF727V3PlScP+b7dv2hEhtg2etDCQ1
aQ7McdpER2hVfClhGxJRqe6W2hboBzx3/FqpNvIu+qoNJkCnO05u2IC4LIOm2WmM
f/zrH0sEN2dS/yvKVi5+3kLvYWc3kzzAjupsya/lLQKdXFH9nTdEsk8/vlrwWJ2z
rXFt+H0IrGEXZiQQ28qd5KMmS4/AvHRF95kSREEG0AhCoPZ2/BS2f0l5IcvNA8k4
Z2w55Ja5bHJ1SW5/8qHpyaApTPljbvkbBiWmAZmTwd9xLyy13b26wew0WWq9vsX/
ZWkHAhauOfT1CPrYMmNO7Hg7VlHqVfhc0V2J35ZCrkFZRyGQWB78mPoNkBtopsUx
sacS9NY9nsHsOvA9wIEs5t81ABWEDPfQ5KcKlQF5TONCZt7hcAOQ8bITv0ggyzjI
Gvd9vD56hfXa5UXf5VRuzw3HuVqx0UInwhoxVLJdj96NIsZppRG6JYx4ylUmBkEl
/RIngsXAO28ch0D2CZB2NuWUQtbxGZ/JvZ8teqQANHZNByII0LjDgIPo1CyQ51Q3
6pigZ7acNXT7yzB6pXvFS5Hjg5W0otE5hYWcphNtdVzl7jJospXKce5xYZGztXKI
04UOEbiCWSXqRIher5+aEu7mZQvsj5F6C5aEYobOzevXve8laz5orvhpEWqGu0aH
vySH3gf5qaVxpJ8IPMyEkxpzLEURZkFlYZIONVPyf8PQOo2f9ZmyM4p9eg+drRjs
JjBkAApEHDoQAg48vmPUq3EhPIPN1vIcNyFmIXFfLgA1r+5wqA8kEdHn07ceneMH
/NfTYQ46CyN/5KImNdf0ebxYVfTClkScahFm3biHbl8QN15tqVyam+xPA64ZVArN
lQ0LbqIzowcAfrdsT1wyOWfmHvAwtrGEWhaYkr8WQMUUeUE2+G2Nsif2q/ACIL9S
c7WvxGatSvD62/GVZOy/TLDJWxXMLwxYdT3z6c2njFB0/Nd/J1TlYhtZiUIn09ao
DcWH868FN9iRjzQTEK/uotQNW8BqJT+PA8drhcmHPh3Rzy+TnyiAs3HjWcwjhdtM
SMkrAxTeSpA74GnoiBidG/wjJW65Ol4ozejZSFoeJMnoU3WbelRRYqH/C38/e7oK
zbHEPUWh7c6GhDr0Npa/unlYRpuHASBFETT9bwEoYJzkgVcf7/Br/1Rc5qDkY1ol
EGSO6NiLwPRytn97jiAXIP6UImHczeT5oa6dQOqSXqFd7dw21NMOEqjz2QXybXkY
P7nU9Gxv9U5pHXq1QUV3Qg1RhEj+nysPkAY/s2RPS5o9+yZKGtfPSzvxQHBNYgPQ
pBmeiJpweIZUHiKl8yQ7JiNaoymn+XFCBqdnlEAmkvgcHp2emzxuAXHSJ2wsBxnS
AYGRcp/hZkYPwsfHZliBr4tK0bbb0OX55fVX/+kfdh1QweCmGiRmN9VX+qjXhmzt
kZefCtxYTV7Rq28klHERnk5u8EG33xF3bMwvkY3ezLuUAN+eJHH0pUZwPk9RlO6l
WIEjzqXrt0X8dm016J2Wh6AujKhFtXw8l6QgfDqtDv3qZiS0PFoEbO1aVb0uANy6
gu4Ho3oDHrJ4lU1Tlo+WrT8bZqpG+nbfkf6ehafD7ZUTvZMj6XKxCf7ptg7Mnesz
RRX90OtpelLCUP+mcr0L/1Ad/+uMmqabnwWGM6671Mh25wFB83srQvBWOriP2Opp
Ju2aZv5wEb2bucM524tCZzb0Zi9aILS5REC9EPn00Dq7/48HPBbsVt0+BoQdYOOL
qXCpP7rnyNkrgxGroGQ9nxLYuBqL8TTkqBN+HRBC+vz0TEf2xDcbsACJGXO3uAs4
A7M7DyQ5Y47xMCNOYoPaLvNZ+YoavO3eimkNF0E3aZUdqfiBrEfr8YzNIbKubSAR
zA7GpD/FukPvU696pFj0dMTIT/8cPTH5fws1gYxcEl6ATQ48k/DbCT/Vzj/5Z4KL
y5Vv/tD2ug0CDWps3M0W0X/pnCXzUN1q1HqysrOWrnOOxFHOHZFBrlfK/oqe93Jp
UP2IRpH82ixfSGJI4QcBsLPUZ6yeGj88aSnAO8FgWCl4pC21a78qXylNxgwAlrNg
3fHRngjmvxhCGigvM1BQv2YJQEaJwjT4n6/mszvTG75sRoLE1e9xbCkd58lNQgZQ
vWag0bJD8do7O8is1w7iC72xQ7C5+DOSdHa06PUDRxZBX20t7MuiTIhdnK0B9bfI
VxhVPgbtpxMgZfTqroNlwERMdcAXgFvyA3+SdgtMAIeNARqo9BMY19oDlGA065oC
JU7oQvvtd+9svmsjF/EdVGSI7Ay66wyCWccnbB0tWtvs1zz76D1Vt8xfG5jdOkru
62xyV3DwW+4xq6jyvr5mEUwVYBzUA4oWC3j6Sotzh38leWgKqoubwEriLEfcrhkn
LH2NwapTxxlcQmhjASqb8f/SC8vHpzN4zPhDKVwzL9hF84NkaT3ac0hgpcnkE2Tw
vQxWIC+ilhBjzDTJdQtNu+1d6K+G48FGGAxe4QLvstj3mLZPCghuxtWDh6j2+xpW
5uSMktIH3f0xGGRthO2XeJGT/TRjflVQWyneybOweVI8WYDMoPFi/euBqyW8l+rH
7m1gr1ePgxFzUjHvggCWGDUx+KqqE0f+YtgBDD67MY9vJ7/54R6dbc0zvdL4e8Hf
31BfaHrfB/nC8xJgOTK6TJiHaEvtQkKc31lVKcRe+g/6hoEuaTy7MqdD8taIaxjZ
CQHUw4zExGeh6sMtlNKnEeBlkJZN4JKkUfddAXeXLoP+9u9Ao3ODouMNmWXFw8Si
mPV2MnmimzYz4skTx9wFpe5FNbvqvuMLUEOuT6g+I7ucg8agn3ex8Rn1Fu4xkXa6
JUCPehAuiQJShYEzGTrjSMctHejupXMy+HNn/hK+ZuN/sPgJgIUONqQU1Z1ZZ2l+
CVYdzsos8fkQdyRniA82Ix1E0sQ92BX0AJJ7iEc7fSdePRzrgtMO2oPMEwSQbfKu
CgOaHlQgOhuLMTAT/PJMWWRyK/XN79peqvYC4Go6gCIGnY1ekZVG1kLHVfQl32m+
Z3kbXnVD/SWJncPgcNJrZY01o7KQhXdqUaPF5/XhjsoAG4YKulMZOi1UP8SGhaNp
JdFxjts6fR71PFVyhxXmH217YPdISLMuomHoHy19iHjhoQ52YL996KyHvLW7XD2q
FPchFqiqv2nwKuItULEEQQeev+eeHtEpmASqJnljgdp/vIaYPYcbmj9JGPYFXTIX
A0vokhubYt4lEoJAJfkbu5RHpCSOXdezv7Ynvw1iTTa9dVwaYSNdq5+laHuDbqTE
ObPSAD152HFD1GDf9pIzpaGyNpy0tY05qP1lqAmIzuaZRapMs8kasYgugffV2hfs
e2waylsQEW6qr7YJkrgRZ5Us/PdFCcICgQ6wl8/g4c7VQ/qMj1W09aogbaM+tXXv
Mc9TnicMYQOpnhDnS2QeCrDbkz+alDY2XAMWOXhTBp7r5uPmF3chrigjwu67T2dW
Oaoi8zrnSsGkC2UZcbVFyqRYwvVvVV5EpATnhOPbkndr1kR/QVOl3QTBXVYpgHi4
LNMYEwwa30niYoRpNS7wYQoAhFMIL5FdeIaYw+8pxMkYtFk5nRzB7geuvoXmkBiy

`pragma protect end_protected
