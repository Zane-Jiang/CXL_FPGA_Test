// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A7s9mSggAvv2862YDoAoynAdgkg3HWBqW43D2dliXj5rW3+QPB4FHt2fdvsE
EfQ3PyFTfr2H6hlr0p/Kh9r9EAKIbb/LLE4Obv+h2+EFpDaOfjVm7QRTeF5R
DoKY4eNLRhKwaLlIoaAsMgmVh+xW8x/W706rL0wpRwBfsJ9rqXLjnrA5+fyd
NXj1MO+B0/ZowdQjhBs9uLBfwr8kT6Bz9JM1LPgxOsPShtVNDl0iBeOtkV8h
VZ2oQGq0UGO20A+FzIO4uyzXHkPeaiHWZYJsWe42Wf8cH1guWAraCjwcNG6+
woPIkvmip+qqDb1uuIsSA3SmXhv+IJ8hngfZC5iySg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JRCHbUCVRp9eGzQLiAtECNpWvQBs5dPtwRIWEZTXnU8la2djxBKyl+WeG7Fj
L4Cl6JvwgQQ0CssWZKKP656udC/F4VHFkP/4u0R766cOi/wz4C74pY4HYTyp
hRrrYpsbVZBPrq3o2XpafZJ9UlX38bJ8KGSPqGkdWchKnG4ySLb5kYKDDol6
PXloDYfDvTCqnDAtD4SWkRyl7oBtNEsBf2+wMSwW5/T2aegWr//VpV2j+T0H
LR2ckh1KSvQsGjKhKea4a7+6zvR262VfC4DlbO6WEsCsSLJnmDQxPi+piTFH
IqfplHVdNb04VaGHzv6GbEfJUB2pPlyVsrjeaD+JnQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
e2SKVWOo7YcqQzU3jzF5C2U0MHQgnChWiqiZC5TxyMJ35gnJbM2ndgTiPZu0
OqoLgepmJLQUbqLmF5LoeuKNl5kNKibuoTxODkaolDjkKI9NIiY7jjm/U3wI
Enqu4u3KyUE8VEN5iyTx7nwhSgl7Ff8LvfAzVhhYJhKe/5mWNqu0QXZsexFX
dLRLaglR3akP2GmhWhvoclnQeTi8DbApo4yUE/LJbtkq/h8dYpzzLyKL20b8
TS/ouPG0w+3B6z+PaGlRQQvZreZKptB4aTjTYkIItWcnrCcQpbbliGr4LahF
ItMJb/OQOytHA4qn550rDwvJGzT1TfiZ6WIjhYXk4w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hc667LZUFczdxlkF44bFPC/aBohX44aJa/h+buTw9tVV/DGVvq/RMPzRwgQb
oDiS18qSbaCjNmsmOqyTF8lAj+M+l+KQUJs0mptIAw9ejt6vNNMKlRbKEDxW
mjKfva9V15aLglZ+LqIBjhYr7CYfcQxDnZNelhu40kMFMI9hbaM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
py3tWcZ9XKiSWKgwyQ5dJ8zY4iSnFDQ0OOd+VOWTXTDcBr/NQWTtlH98m038
jz8b3tvhMBQEdAVzotQfADxSjBjuIfCswqKgcOR++4dot0SCqzudkLuem4jj
+ggJzN+PdsChQgw3ikcyt8Is5HeyUaVt8QOiILqEelUI3XJo4BZVC7ql95Vm
q3+S2eKf+Kc8bbrXqcsFZIMmDbLePz9dv+t88Gw1xGXN/LnN1xIj/QVHqOW9
oPZeW0WCY3CDXJAupq/+Y4N0IkEOnRMGCFRvNcxsUjcUTzzDgu+YI37UcluD
CPWLenvcZpKF3NfFGEPX5/RD5iwu8P9qkCulqtKF3MNcy6Jnp/4noOH6HKXR
Vq078jOULgWYZxIw6zc7jDI7Bns3YcvDS7+1TRWhfhrNaQTdCCvi6r3CIhYg
o0Z2QZtRDtrv1QlYHEJVXzz8fjLHF3LP68KUXZvrBHLhfI3rer5A2jJ7QIoS
WVqmzbhEEXAtwljsZgAz8XC64sHxEf1c


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bwhmrqkHDUdL9hSJr24E4gG4YHUhaMMZe/Loi8W3oV5X2Ojlpp7l1p+iw63q
eL5wCVq+WUJXmVzablGyPnPB2keSH2BprkbmUqH3v5GRVTPlvew2jtdWW4DX
dq/0wpvOdDg8bObq38nNFg7fQeQ1LJyAK7rXCzclr/QqwL79Alc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iWL1TD3E7VuQuMPV2VeQWeSVECIO1ZulTsNGdCwezaRLMgmhtlqFvifa5nWV
IVP2dB/8HdwU5SEmgvz0dSe1zfb3cOTtHyZEWQKWjqB8xMOLPJbYuAFfDri7
MhhCJ6xUsg8ysd4Lp3OivBW7LCpqVPAKGfzf6KDZ2Cvmbr68860=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8976)
`pragma protect data_block
RJmj63NF0nVsCJAVfW+kpiPOAqmQ3KBW/EaSV315kI1FgOOvI+lERPqYxgLb
TUqKrtsn1s4H8L1sb3ic+87uwE6uIKbuqOG0++JL/KuZcxmamyEFPuhGxa7W
v9bbPzxHBgq8YW6dU0tpXfWWnTHPXYHXUy+pnCoIZJlKdX2ksWP6B3QrP9Xx
vfrGT3TRosru2IXb21vzbpYinU1U/GZww6xLurBKX5/sG2QnfpcnEDXIPs2z
mRVGXhIfvrQfkBOfnn0098tOE7XbaT2bf63S/S7iQ8lVn/eJ56bpw6q7/L46
TwhckWBVN3Bbu8iQiYPEwOTH4hWD+E0W++67AW91AAMNSPOyp2nKXzMwsCQI
pcpEpSJEEjfrdJCY2mdJ2qp0pMlfHHmAMcwOYcgBeUVj1kq5VjcAN0sG7m5B
qb3QtMlXztQqA666vwAxg+aEj4E6sCnzm7WCNHxVhy+PVvL2Y5jju7RDBIY6
uyuaJIRVHjQY/hd30maryzCunkIQYXcNxlnwOpHC5A1pOyDYwcomZVjd77D3
lPuHYsiTosqU0jiJOkHxyboHP2yU6D9AlLH8yzBrCa3TG9sSE7wXreiCJkqV
TXoNRzLqXmOyAwpzSEip/vWcSYqGe8ns2pNZKlm+C5V7peMXimzm8Plg/sw+
wcUbGPxNx80E5krAtPjSt1GCl54wgs0WmWCMEpbOBu1WN1FDk0b8I4d7J3RV
3OGt0K4OIhIHVoyMsqhostdJf15hmbXqlTNh3AB4WZrKdGxu3l45ZtMYbI6j
+4veGqiApoyUv14ksLpuOjjGJIN5eiCxRoOqjqv7OODxeu11uhP/BLdHgThZ
WJLbfsVEuYnz7NImnQrQe52Zzu7iyotffmCPPJlkZhAy8XcyFwdxiUvhWkvy
l26C0dte7nCTaVzcEe1DTZR5C3OPkMFvIOSLFAZfVbq/L7AKy6CTioSnpdYM
8kCBE5cxtzlOgNAzYXnbyQQoIrrmJDMXe2kNbX6kynKCrOA+t1QKoaYqrQYX
hRDl+eDM83YhN3JjsAdDcGDAj6bzaoM10F7aXGtli0BVORCe2yngVsFUwd59
0Equ4oYEPCSn3dbcwYtiBhb04n16eOPXS9+7z8cDnjopRs8UIX19jR1HJdAV
5znEKks0AWxys58M9aSaxy5WnJJPRE3gFyy0eX2YUlad9LGhnoEOhxxglNLY
71TyS1vxjFIoMpZZk+nsQ2Ik2Ezl1JL2GIEQwkxfrcffAGrN8FN5zOO7H2ht
C3+n7Ri8HEzyiXCjD2CYjYCMAlLFHbHaVihYfkcy9SHzaraLxT5PR1NPcujv
nmfF5N1z2R1ENCYtIYgGNpPxa/gqVwo+0HI7C6nv2KRZ2MMr0o3m93hgmtDb
yB02kOhxDAfb12y/72eHfnqGo5YaoiRHIbpN6HUwR9xPxIRZZbn3c9Tgceof
dyDe8sYrfifcHZJAUNKtY8ANlpCYyCrOon8IkGOy4s8XooLXDcSUo3MdImNn
a0jdaAXplkIHS/suCX0AZzun3mQuoBnm89QrbLVXJyFgWgFLGHP8D1diRdYg
PEwr8d3TB4buKGZC0ORVowyZOT0kYduataIJvJrNUxypZDwM0Y61qMq5OxG5
A04FhD7NbtgUeBJX0uN/d5de4qLEPPxReIyciX2q0yVZ5m1wm2ESXhc/uxVY
u39ZaLepCnElrDFJ9QP15Z/CMV21RDZ027y+t3/Y3wmPZGyB/J4j7SKum08P
7WUxmy0cigZRe2+WtxkUlQmlgtrIga1rhCN7zFIudztqLA43UlTi1pXVfRCL
CuI3CVcwR0Hew9tLI4IWJ+dF8XSR9fiaYnKuLci7JKiYMSJhLv3c5HRSwCw1
BpEtVp/88ug3TeyKmJselJUWECxA+Y0dX6kLGSnX/ExKJbFesabITp22JIgq
O0RuYsis6XEsIr7kvKWXorQZmyDCq7GWyRCQnFoDx2EoV8Hby5KnwMbSrkNr
cGQcNaamopfIO9UKewMjYhzbsirH8L1cr+1xQ3Ld+BE/afm0AyHbxwTuZyFo
M4u6f/8DspYT6ENCwfFINriDIyBNkdrn7hIcA8Mf4gf4yU6ad3bbb9qvn6p4
RLPgU8kkK9JxGuFecVYpB8Kyuv+80S2VgkrEiTmuslR15A7Iocc0CbfoO2aP
gHAnl/6OMTaBbntZett8zUCzFgNYh7C7r7PqzLR0t94JOzxvD7b1wSHhU5pv
VUQRAB6MKv0Oqb2u7EgG5DVBVAzYPEVbGh19GwMjLf4lI/xGMObHRDKdznyE
G7rDSwQ7Nop2srSghmnugG0VQP5QHUFzcYZlWH8kPiq+6tBz/1EleYlc7z/r
LHAQaXJMjSw44CXth9B2+lv9b1AY9xSABUsEJqe4E4pZLzAX0MYyNVDm6A09
TZBV2T3lBauOaa+0lka7HmR7xVQul/8z24unroZFXhPH+8rlyJ4/ESFF0Smc
MBuSsdx0f7tmIlJg/qPW9pg3SWcSo4TAEiCGB9WxERK1BYZkM+VGNS6sVKbU
FCg0Y7i53gpUhl14OV7smspVqclLiHpHdQqYu8Ou9VX35fi8QBtuY1b+psfe
w07IAQ+GTJueugF5mbJyD8OmN33PxqJx1sVz9qzRH4L/vAsxKPqrcZ8l6klK
Wk1plEDbJ/ckDKZRRiL4SjKgFYaIx0dduyZhnefBGnGivzP+aQwnzYPJHzae
+B9V5FCLpv82v5X0fQrC8CP3V4S+xLzovg3+SATzb9gW8i2K2O4O5swoTPa8
1WZXvA0o0TRYGAxkvEXwYVbxJZnodsW38W940yllUmt5yiqOceEQCKaOoKjG
7JRJk1cz+L4bOUReIVWh1LJfcwPuxDAmgNC2N0ckMtjdiDgBC2qXeDx18pwO
5oSQ/nqWckJ+7Gh7w3cf0VcahBVtiMpav6ZXNAuBC7N0JmwIP8wiVWkKptNR
hj0/Yx36xeGP1akW6e7z9BFfkUbiUTYH+Uj6i+ZLsvXRz4X7IBReWDuPbAVL
CJ2LrPTE76Gc05+ObzYi89wO0fe7O8lC1o/X2kGN4DzbJqdtSUwHlMgIxBEn
+7U+sT94x1zr43xsMFgBqN+bc8CnCgILFicpV+Eba3bhkpTrnwU1JdnpSA+F
YrVsF0mOgZ0XuYqCTeHfeH5kxXjwLg0+KMsNADmi4OsiYFylJ92I+3JwgXh5
fWtEeYBozdoTP7sZLt4rpXaa0R54RRfw1OY8Z+BjXptSlGqiK7PRCpv5TDKa
SUZsqH2BJtVtiLa9hHewDUU+1QTr9oVLM9t+3SXNHQHmg+wu1C4ctKVNTI6M
N/vP4p41RFFLWPnsWNxxR9APXMinOyQvUarKFUY0anT/Q7t05UGPmtHqUJWO
TGpD9Lc/SGtis0kGgkr/W8AL4Oic+Dv2/u+seWEbv43rPYRiTxAr+wvP8hCl
lLNWUfBHq+KAZpuQ3jdygcqPYv0msmIPqBfY016KoV2ZQ8I5OHawygCZcdlx
OMK05VhgTR9O/33isVXlvjeNHdHCw471xBGMXGbvFjAFDMRunYpBSkshtdbB
l+ySVbMtMUFSVPsyykiMlM2dKNjb02ZautxMMe6fWxgNRLblS9dmkyI6SI5r
3DmkLLCd0qDOlmYmueKmbYyb3M/WzZsJ+rS0sVQ2bUxGPCt8Kd3jwdwE581W
XAc/GfLbP7pSZhl+WMT59Wwq5eB9XdfkjZ+7IoUEGCHPBkhSZydFezmJ/K73
mEkS7l+FrMQpE2++2S81DOx4L0jjnY+Ky6KjoZ8k30WuERzyJRWhZxNNq5Zd
EwtvpJVUMs/J6GwEqJonNvBasY/NvFLWjjxwzyv18mgEXoYD+dhXkdX18IFs
9g1WYMokjSipS2oGvpO/7azzCYS0CFfOzW9VJ/h/SK8L1XXy5IfiDzxD9Sc8
/EliNXKBWNaPuDYcAyudoWFzow730i6QlzMVLTwJ4vVoqahgihx/H1V7kKYh
1bpShvHl17ejO6SAcSZ4udSVHiUiooepwpBnRjTHEip3gQWpYMH5F28WznLe
UEvfoHGlOQgo2embOj9Jv+FBWY2ckqSbFAPkfAkz72FA++XfZdNr0MYGZdv5
en3oAp05SBLd2GUrV3yeKzJo0h0jq76MAhRwYxZJNRe2R2/YgxLOZlhEXWud
jeLvT5P3ttegVydZer1qYzUdvry/JEO9tveZMiWr64gvNqp7eepnRrOMyAsY
EH8oSW8ePdh4BgM9zjEg2LnQdFEwqsQv3g7Z56RiZk0ZHIrgK8LMUTPj16JB
qqBog6OMQzJ57+4+IXvWn+z8pckIxv2VgUcIoEMYTOUrPJ7RUAsnKwuFTNap
PuOEG+PcZwzzYmyJRLN0eplulW87xAd0HCFr9m5mBlQv1BWCk3/FZs2kLCYb
zf4s4Rc5mN5uib5Iei+ipRg+ECOL+3NSt3t+lsdzrpsoHhhW8zNITRKqTLTD
QuPDC6Sr0FjZh0ccN+/poCqZ472w8JqQ3noQ0uYnSBIQMWOWkoUgw0J1aFoI
fpBHRLgODYP3DXiXJj97YeqWNnzxdRXKGNslj6aQLbz+X9vO9f4/khtwaSlS
ytJQvlB8eJpYTzApkDJaKKEFmeNNItOqHh7abpckgiVipEbcQJy5KPY8I1bK
HDSH9THVsVik/4h03D4penEpah+PoDLY3E9UW10P4Hj1GM031yINnBpFIgnl
7QewiGMwNguarLS37dTZjhcBwwNgC8jX8y/LTmwor35rpTEmYC/o9IR3UgYX
1LGhL/1MMcECqA8+ZJg6vsYaaBzs2tJfAxlvDUg7ZGabcJmPThzMfPhUHoPE
PTV3m7qG4EDovbWCB9TbYYlKT373sDzV2Y1Ktz0ac1A66U33to0oiwCINoQQ
soQZ9T/b5364uyRF739TGT1lHUmC3P0qiPRr6pEAP8jECEwK/qaALkeVt5vh
iZPtoecl7NH4ElSDUe7YHemyCw25k/EqT3D/+LuainPxmoVxUKRmc3djzAaF
Luh6GAobepsDVoDAEvD2XgI8eEHLceb7iTsTIYypzrs9xjTyDRCBwnuyDJMC
i70FdIGG9UcxXia2Zg15TCeeJ7sR3nb2p3z4AEfs5NKm5pFIGyh8YTX+YDOF
zuEiDUZ7OUZjhlm/Tjnh801FOJDakMuJm+KL1VFOVh+mvO/CFZno3cJkXGnE
SPlxw3SXYC+xFClGnPUZyCALpgIkzIJlBurQGumu8imgCuihdYw/aeE+Zkpi
nEtV5XW+QrbUobsrviNCXCYuAvvpTIVUHw/p2Zpz1V99OB3IrulYbTc2H4qe
EyoCHBba+n6GwTyiwv04vb5CsOLypMWSCpv+cDibBYST7f2kwKGT+fPupra8
CA8LR/yENDTz4uJnaPgNBsVkueZ0ZGptHkoLwCstOkGfMTfBD1CmgZolqm+P
sxkZRUNc94+jPCNWxFPxgcN87liu0u80wDiQPvOtPLwXlVKgguULXpqjr1T7
9bacsHpXijLxVUw3aXWPK3nALNlc1HGNK2Z9X4Y/lx0PlI0S2+xdrSzz030I
cE30sJ4LinCkn6vQLZmhDorEFPIWTu3WQGnqkUqwEABXTnSJT8NGnhKTB6eI
QfwsPsKeOm3fTvmHmbOLq918v6qWxMM78bXC9PMG/YF75MutvDx99vr5soZM
J8OaHDrgVSOfDgZ3fqOohAepPwxz/Nhdd2YiJWxN6wD33U+wvO60D0v57zY8
TBnzm9nB6HXh7cWY4BxOrimRz9hgeFBLUk4t04syIWlPD5zDF88jdj/DGAui
/dwZYgbiN7OxlSS/iX5yYnD3vnzI8z8sLinrbtcp+VS0/7OwUJOIEqPpB+yZ
XlYPJP4ERx6MDoRMN42YK3VsRhHT+CfnRe7LlE6KfF1q22Uu9Z6MtsEA4Doo
/MR7GzOy5L78lWXINWE9iPRhwPyZkF4tGAF0JTGBXCUurXowjkx53Ww3R17B
bpz0faQhk2Myv3ko1TD4ns4mOQIaKEqRG0oPUl/GBYYpu6EvGUeZqHO5leZu
E4tBkaWAqi9pzZQCg+g0w9TYY1HTnAcIeFw4jX+vz7XjLMGTMugKsn6IMuis
YRG8QC/43yDwaPFxj/7giirPY/T5ZTZM9ljQ4DOiQKTcRyh1H20XIyyo8a+6
McjljKDnuW7m7hmva1h3LZ9ZVx0/ZtSU5ngdUiDnr9VSdpC1GhksAJ182ZP2
QCiVl6dbGnPnpz/pCUFWV2Gt16CT7ETX+sluxLAhH0MFCrGoMlKIplIhic9j
teHYxS/tkIoQ8aLD+QrWEMmkhMqRpE7mC90bxPIJvksXa0xPsU16MHYGs7LQ
DafuQQKFN4Y+Cfn2AN5x9aXqRBUt0a4IBo/oHTxCtBiLwxHsDw2OTT9r+wQQ
TPgfjulml7MBISg6q4WSSz/+NFzshxSFkgjgOpVEczlw6r3uRgu/Q+sKfl8B
xALKvMSC+C+QMNpmB1Hm9OkXC65c8oLSYpFNy6SnhF+ExpoOfPN/fqf6LhDS
ZwZUfMbatYYLAzQk3eUtzr6C1xE9zBmoglV57BY67GuPabIMItQcfKC7veJJ
YXQABHrZWSEt1QbXjBo0q5ogi/vwLC7aGN1Paw2sTykQuQSztJ7MR6NIeCFq
pokyQ5tnQ90LIVeoFKfAJR9K1kK1Drw8TCH8Lqpx0PG/EwFj04J4b3U9Bs9T
vzXPhEuhogsppuYBI/QJ37MMHjosdher38d5lNoRGW57mGhVj/eMYfIjGHi/
9o8HTMGdhtJQ83Q44ZXFZyo2E6sG6WVa7pain3C2UvC7G3m3fm5r+6EMc1zE
f5RZs5d34givnCpVO8BnEiNhayPYN9A+8RKDuNLieKM31TTk3yKnAhgLTONu
qA8hjDWPgw2fHaSdWU70DRizviov0NwQXVGlXjGUdxKNt0YC1634/9caBQgI
1Nay41wMk9zeMl74M8EGoLilkALHeqD0Gb7GoU5xOjcUsCSJUE4UBvUSsh47
pLX7e1JVKcCHqbYclAZfCaymJqbXdDZCOMBOBg8FYO8byO5v+dXCAvYtUHY3
qqPdy18rJer2ziDLZfYVCOgFWTRkPTUGqSTxul2EbwpUQuOiEttJ99rL46O8
9h7D179d2Q+Jr6WoWiX+gQO97+h0ogsgXyRN3Pkoq11ASsJPOu+0OjHBFIbN
hqsMjoPJiBoRanKc3HILtfOyhm/A6Pn4851R725LakJ0PaMgAokqnK6m0jX8
62AuPt1ysE/9yjkrfqGBX5H7JCg2Al/5FGcw2JWpR+aYuBqiR7mECBMnzphw
mJZg1aFTKsw40aPQGqF/PoVdZ5xb0VBnu9CQGnIg2DPOCiHzAJbzq5xcZSBz
1fum0b5tskWI/D/6jcW4zo1eQiohmzEwq78kkhuTJguOm5DWU9MWOVpk+9ip
d6hb8faAfcyI4VZIGQq9wkDjPe++s/C3oMY+kj+iXzvsgUgxRG3N1rwqX+7B
DP2zADwotFdd9wKYg1yS3U5H4gZpsDNNOepzitHonq9w1dvBl2JJESI5BaxN
wycOnkWMkn9eY4gDhJynaqPu0LKyNNtKx7RepfGzQcPnaD/CvUQhqOuJGiZr
IqJDN3BGrlEK2gOkAt/NqbbYD2vwrzy74I3xcHNFgbJb0yCrmX1o55rjVruV
ipVVClH2L45mBCFWYNRDhbqmOx3AsFfaFh3twUbXuLRysIux0H9pOY6/UzBe
bwEERso5dNtsR0xSA90hnWbqnbh9MAZCTiuXe2daZlTPovLakOcN5+dYZnwc
deFDLJPdlzfYvFC0RWEBn0fKQTqiRtYZxmAzFaxr3zyjp542AqgFQvgmHkYh
FLKhk9ZtdSMOSW3/GWs1RxRd1UP07ccQgxl590uMDe0N1Y8JTd+4dK/V75KL
LyNhKa4kff4VuS+qZU1yvAYYGZELZsC4Wvj7Y8M34jExNxTrq4fwlZYfFE+C
F6sCsRo8kCApWhTUNDIKRgKCXQtqqYhmYjcusUEmkEYVN7y0ZDmYz9ZD04+T
OIeF2MpMPJ1ghpE8zagkG+mPa2mM7Q4M1YYkOnAjpoWq/4JnsEMS9HgYahqT
7qm5rhr+/+rsku+/TpYdvQPdUzVxQIO/rdeXjVOEHfguoprJlfE/wIPYVpXz
5pEYN+3SHEKgINC+afPUaolxc5M0M1GiCXKyXlSeyw/kVXyAzecHAIrh8S12
LcHwdGsue+bUKzdPQQeUEs5pXmPqe3XcfjXnZM1OcTGTfIeL1p9IyoVRjKbp
aohzhMvMoDX1uGQy5ojiyPCsxKn7Sac1RfXcUFxa3VSDY5CsqZnBYVxD+BK+
rAXce5sXSJVFU4jVfbGuGfYFapsEJrDOvFacAbD9tUuaXxGlts0xKQQLlz2X
Zh52PuUtevv/PFBNrN5NqkMDN9n9yWYxzLGRljl0RHBSew442lnJmlPE+M2U
tlpPUc3nolqWbrrj1nTqU5Kna6JiyvpLyPWyOW+TdUIqf0Np6htkEAI3+X17
to1aCpUE+lAnRnan0aABnOCB2+DZbfxZrdkVMoGTMfM7HUviH3Wv3fDuYiBB
k8ZcpXv4t3vlo/X2Ek6ZCN9jjWTytCg3ZZYAEBapQbzgY/ATC/f5yz/CsHxZ
5bCPkxXUMAe25i2hwjLWthF4PbERaPi6ExFhjr5yUwOPmkgZ5397dK/AEc2v
8Y20BSrclulQfNfcCps1U0CNv3sWFSbVJKO6TLAvLSwV3P62zJL1718TVgy/
kpQrYS9Zhzhxb3FobkkBm7R8lvJukFNjB5SYsD5+dxc/lCNBDu3LNkOaSXI0
Ia2qR4XPkjJOUCsymahoxHgn8pm9LTiKREY///OaZrLK0TNW6p8BE0N0FcXP
HmFWrH+dWtnbNiqkdJevliEB8pCJy9j3dA63Gih7KvP3ee0VT7tCqpbttmmT
qYOnbJIOAMyH58tgF3T7vgSs7iRCrMAxYWLgyaTYPk9BfKwRn77YaiDVnt8w
b5o9R5BM4PmwrgB/Gd7WMdTsxKzYMnBMuFsYLgtfLzg6H4huErf3/1xkSq/n
cAQND/VCPr1yweQ8YuXcigsG9Lwnws7LfxZuV3O7BV9clGpSujZSgWYwhy//
NMPakDHxiWjp7G8GPISg0yn4y12qHnEzCkAFx/qwx6IeKyZ0hYBVpoQ375w+
YZnV8ALn5t5uyWSat2a20zRqbFVx3ueFP6nD3rOvgtsCEd66c8eJCXY0zFnb
jeLr2DseoEts3UvgOogLOSv8jz7z/6qe4mVJQFdrImWjs6tz9RW9VawUGms5
c8mq8hmkAV1+SisdCvc6T8sAYYSzRt7u2UfOUgRptf1F+fr/W6xMF8wskGso
xYeCzYtp5Bn0UknKcrT4nuPSo+oL8YG/ATK9cpFiXWDBCP4vA5YR8LDt4/8T
FWqgjXWJqfK6rTQXnVClQjIRzxlZyQVMeiWEy2pzL/7J4COEle9bfJ4LISNI
YLlViinsx1P3qKMZ2iWF4PkwBsO0cGgFWYe0sokNkVEz5kHsewRrBhGj4e9Z
z0hxDaHP8m8l5QJu8LzA6/xK/r2pjMHH3iIPYOBdY3u3pM+F6Z7XcEwJCE/N
MWmlMCKmarVKOf0/eHF2D1lghCndcv/H7u6TYbdhr+pCE9VlKTrAecRbxEw6
CrSgaok7UhRgXJC2rdrn5r7Mu1zxh58tyIxYiYnJS/zHem5GD6YbKuyk6yIL
KZo18GKecTEreIa96nC4SnnBedD22nvHi4PyMwMvNSL4fweKAUndBtI62DMY
klpX5Xhj44DYTpl9vIs1u9OgKec3VT6OZ9YAOBf1Nwu9VBw0v0WzEeE43+ZY
AQhnwAyafUq9NIwbtNQKoXuxtsV2RhOo5OqfR0V761s+BTj0z8mDUgfG6NiQ
irll2SSLmzl7yEwH+nx+BCJ/q8C6/2nvFmbRHyrNSh/CNYWrj7CJWdaLbJQf
HHYVCBKDgavLFFrfsCG7xJqSG7+NSzimqjwruFRsR+yomPxEOLsa0ZyDUocZ
63CitKsWrL70WFDtvSpk8NT5YetZdMc5GB92u2sHSxPcjHHx28yEdzoHAOgi
5qUVYKYpjMA8EmZDOjS/fK4pEaxm8zNSw1FGZJ8dU+va4QX0igY3nopln1YV
PSMtCEWiDG71CBJg7AtgzDZRTaLx2QjKhI6dR3KF2CTO5ONCLkp5LWrZxtRb
Zd8X2WJxbV8qf+3naQwd31ktFFZaP9vmbhQiJidN0cEunosd+O8+9k9ARCBI
1q6SbIwRujdL9bwvAiK8it822lJf6Dv8IgCUriJcdhOanwrAdUX+pl2tliwJ
CbAx0TxSYMUVjxWNEtkR6LqVYJD5HrA+Ejk2IZkNuXv5HtfFLTSOXJ0ZlQHA
bpfLN80iMd6gclNRX1GYCeLaMZN/XrwSpWMNFSemxNknqUJGqUG52iNBfQ6h
uaE8cMSrBmraAUDsKv6DfDohQgaUCQJetUKVWHocI5p6y9hH+IR9ajt44UZG
TLybcjaLJVxTF3VDhwULAI3Px5769VvFTgliFXVq2JKAN0SwtQom96enb4Sd
aU/6vtNZnLJwI4MWC83P8JJ5oE49raNnka7OSYTU7LN5dNS1IQ5+peIGbMVl
fSfY06QpSh2M2Caf0wMBQ8f86mFxDaDzjt0Tgv8MrsTGUB987ikcwq8vKiUz
WIEDc2+1v8uCEa1VEw1PSIzEJSViU5Pf0Ue33F9w2mSgtOhe4XUzPpV+jZbS
4y9lKtn8PWwgQk9ei+FgclBInu3e3Ngiw0L7exRwfAQJWi4zSoWKSqZCFqNe
DydJ8FlnTZFhnKga7dIIc0sIOmkxuwF/K9KNo9YydRJ5zMg/iUw3iPtoMQcK
NzRv3H06Ib4DMfxMRgQ0QmtASljiNikc6+TyOoI/EvnO7WnoFe76nNT7Bqb2
ZjlMnYLCYb0zvZ2CWLb3kt2pe6TzzqChh8ohu8e30K9rZQfzEQzxSCnoF3we
z9lpV/uWNUUmf3ZVRCPBsqNfLFe5WvmfB8Wz22Wx80nP/8RdxbVuRfa7T0E+
D1DYLbMZwwr5bfz8U/Wxlk6fccJhO7x8GLyXzY7ykRAWlT9O4sM9y9yvNBTH
r6bWJDEZJchwg4Pwjp5uG8jAkHV7jyfawtR97TJI3UsxHC0/UAVfZ4oWUNy+
WDOEtSZyjhO3XsKH6KM6/VRtWRvURHE+dh1UXdpGj7uFTtidoIgzUoYmf2lY
LWD1r9dd0l/wx4g5tE67Rx5EOat/ohtqXVa1tLoweOz35GI3IQqDB0T+NoYD
DZiASnCn+VnX4HUktGVYEAnFlPRSuGZ1PooicGltx+Ra73/gTuh1AqRInCje
WWuZ46ioFUo016+4Y+R2dzyTgPUVmn11EmXSL9uFX3wajBTfE1PBN0fVp6HC
5bjsF1/0Zpb26uY4OzbNx1BglielZFYCLO5tcPh43xMkPwJS9cGkxjbnTfvV
Yi+6T6akcN9jl+R1wuTI7CiKrC2zLbSLX+/dQNOSGdj66KrfSbVy75bLicP3
rNE9T9881BYo1+q32dfDfll2SLjxz9Zj9mLSQdEwc+bO2mPHw3C4fK41j+12
QvafbLroCaogzXYwP7U1fsA/b7IF3YiOlHb7BHAPO4Ph1itnqeIpS1CfTc7G
V+9CP6aFTEIIyEBQcg9UmVRxtTcZ5FHwLyeTelCuW22Hgw+vs29yJUIfRQHK
Hv/dZgW0YDj/Y17UL5D1FQOByBoc2WILcOecOguvsm25rd+ks0xtCVuHb3QP
zVkFVEUhy7Kc2Fg0ZrxfMEfyqDYblwcJaHUwZ67i+Kn5d0lz4JQLL/NUMAst
pXHKN/44QmhBgDQkbkE7YEA3hWoU6wGEWnmirmVNSswOCmW8SCD0KxxgjiHx
wItL/eBWqzlrDayTntukYPJ+Amjw2Lx1b+D18coqZ6yfYicPwVx3DrJ00lli
5OR7uwG8+/ckwiMiA9e1zBNXYAz9gBnkg6En/R7xTUypAqdIMmtiVkWPPdBp
vSljszPZ5UYqYZtdq8IhoQaJt7nx

`pragma protect end_protected
