`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
KkaZFs8r0zm6AW/cAP0bDR5jq8YKED5HTIvYupXle0WF5EALwuY6ql1/KSKdXIWF
6MpwlPkcG0V9NXjUNT9Tk4U+X30Ap7EROvJgMi0mDA5RYKN1BjL6zVzV23XEIjH+
DEGGXhowMPmwczwEYguQWBm1zkysT03RcrX1y3XWW3s=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8848), data_block
V6PxycEGBou7YtL5r+3+3DmjuBoCeJYNwI7IPWJBjOUzBZxv0+z9/IGvVWl0DrzL
LOOjIDdWrcRW7WRciRo0jZ5L+MnZXl3C3GJY9yCMbe5YTDeL3hTxARyLl6HF6lD9
Eohquulhb5sTnuobJ6AfByqsvAMmOIrIuAmzxPSkaLeaZh9pzLCXFwyKAKA08g0p
e0Jrr9XjbWRgPAp2GQvQ+CmRy6R0HV7b4Do4WX6+zQkKlNfpUUOqwyQj83YsqfRw
kdXfio72WBXR7qTkbs2DUZ0d/XcTBwO9f1HQv2TYbvOvFtaZsuq/WQkFPv9f3UOa
C31uypGP2XNOtmwC5CP0yxYoCZrZVKbzsd4yfrtbObvzFkXb0kv/sY7SQU3neVVp
iCqbtt5kRs9T6FLfyR4USVtwdsLibNZnltZLkFqZR+Esz+sAxedg3aRLGv9Cbkb2
wHkeGb1dP8NDsOxD2kp1Y33j7TUp8ecnDlvURQneouBVBPAvEzB/aHzH8Dqs6n/x
auq5Ka3IHvd32G8K7a6q53o6iy9d7UDDUPjDN6qk8Wgb/sdqKH+LEEfyOYn9TOix
XyuKkOaW/0wPZTlN/fLUSptJJcG7CQplEgPhC2vWOddzcLNjoph9iy6Aib80T5La
WSVIybtgQyLqNZdwq9UqzdumKCck3cFyNDUV8bwfchEx2CyllFcksfDWC6Rpb8v8
DLFGZSEwk+BvHGs387k9lhADeCRw7/TV0IM/xASUhFWLqw8eTcaHyA+1zRNtFQt4
kPTzfhsjXiCuqLzArQ4eipFWzr0EnUt04HHAUSFzCxNRxSOHLX2rDItS97r5aC5j
JFKGjXCszBtykSCDBFpgnt60+XM2qpQLNrmNmv8S0tnf8fjWtaBIFkFNGUgv96Q6
3e9+B29v/SFOktyMEkxcsaG5Kv4EoHvvwDSJfzw6sNsqMYCtgvI3MdGne2sdRjNz
mnbwZAo/BffhZkrqMpV1HjSG4Awl12j+qcbLFxnSl7Nolk7aSa7fxVdDFJOTYUBT
uBvbBOCva8FLjbaT7jSg8zt6o68i049jEDzikDERplpdX71wvimwe6hZsd3FQvmD
k2kTwItGV/YhrB4177WsObmPzrRGic/0Pmr8lprX4TlB6Nr28ngqH0OMXUJNBF83
LvnPsWoppxjdMBiFo6mdMM66wemM48cAEFLm3YIXTzpZGkumnFHvVgaT5EM1a/5Z
o7Pr2O+Dy1Gj9UzG2P9idhSAS+VMlBinNb1c4Em3Lfs+8pgz0e4J2JrowyA0ib/Y
jFmnrwKfRN4WkbRtsaCJC5h5LA88Moawy2wGMxo2eZMZll0KACOxCSZQSYwXqljz
UTUC6LLujMOmwx0CCePIeZhkgJJZrl+d8MS+5pZE9dttbCbNdsLin5IYPPSzn3E/
Kc6yxOzehNMsCEF+P0H5jrTQHQ54mzKd/d9Z1VyGWulcQPtIr9ECoyFCwdl/sGe9
tZKMDfpHFKjRFnrmrq9y4JDgWXoyzauIqvUXnSI4m5x00vOw5lhbS2BBe5H/HxkE
kqc532zAVpAK69VJS+zdjy0DFSHjG6SbeXiW0hr3gMEzcds1OEyiuH8j456+JvDo
IerfXN4bbugJfif4JNSbH+E+x/+cJDE6rOiJ5qWbRBRXNsGyxiwm3YZo/2b3nkAR
p4aINbEPFzbzrSCtQd2HMd8583WUFmr/QLfPL4nxL0eZpujLK0z4VJDk2Mh3Hdf1
WyB96jHweB7faQ8vl7gXqlz3LQ+82JPyM8QayY3uKVXZpYpsqruF1hjuYXB/ZU8n
Q+wJ7j1a6JepT+YbhJgcChvmhlsvlazI6UuXyMip75gS1jSUfYnWgtdLiatfn86Y
wj7O+N9k4pwdHq2Diez39kgihKdGT+y71bxuLz4XzleP4uUYTHN0Z6xzzYQaiE/p
qBpSejzM7agrv/fT+3Z2KZv6EcJ/97VikrrMRGb2a7ab+MoQe3myOb4gTDyN0kui
rgCc832Fz7drC6/xc4S/9a/053eA+QtwkdmrJVHKMPXjW1aXLLLAflIiH4LGwl3f
oRahIUhRj5IHbV8ngRtV9xeBavyeORrp6YKaAzf8WhV6qvoPxEpWTcaXYxi8RKi/
QgHFpYllJCerE/CMU7iSfpPkZeMM0BfCVvl7opjc7BBvBF43QJobpPA0chk6PaEz
wMseKxJkQ1TxQTNuSxYU3Gf/Pj1IU3BjHaq7GzAju2UdEOtev/BY7cBKakhVjvGL
fxEyic0WUBDLxTcAAalD6zl2MNt0ZLaxKfrbZN+A5LhmcZk7h7J0z+I1zr9Yhlfe
k0563Qb+uw+Azme29KR7Oq7G1ZQgw8pIUI64rOqptxmc4jFpJ9uGWFvFhiMLWwZA
3PGT7YRpq/xydd1+z9S6ddj80Tf2E/V7St5pY0XjNl8k4hyFWq0hYIhpyOA1JT7q
PqMXqqUavMUxkulUyZ7LixVMEqIfvRT+zhtMxHMLYru+4+n9KsANcvHg2rh/TPpN
xaH2OBBiyDwbVPOKCP3iPRqJKxuRC6nYGKucNPgRP/RwXNQzYOFGfHb2Lruzc4VO
SFIddufXvdvfkc2/caLuE7ZpZKIAk6pTeayRFF2h8JRpKj/jU5e+Lrnwc/eLdIPW
MqCyZ/hvWtFbkGtQMF7aWCiR1cSz79YixNtNhZzKNpOKMuofobWx6nJ5QRCGBgxB
9G4sEDWZ3oJ+fCa0a1x2/Kh/PpFZIi2dRpgO/PpctgsFfDy0SHkkqIWvxxRG7EfQ
Gqafwq9/9Ki2VWoFZnmQcghuU3apkVdif04OdTWdjch4htjK49Tw75sJzXEV4J6M
r2PwMRqQXErUg2BJHypZWGX3bjSrgtMqkEPTkheib9q9feqO2tvpIs/SeOx9O/Oe
oUwq60cihl1IPuRimzikwRGjdfIvWQqTLgEml5zakbiTIJ2knhSSazOd/jSTizNM
fWksH8HWlaWOTJXpGJ4/r001wHVMet6iUMa4Z9aPYn+g046mKDYfwZL7tLv/H+jR
C1+2C3sZZb0eagNmyUM49W94Yolcze3IOjGWDttpPAho5JloG4he9pMmTrnObK/j
2Y2i4PF9YIlQ9KSI3tq6viduY1N2sSluJMOCe6A3LgZQaQnYtDYPpkkA/P/PTE1X
VRdiCzGKWgtcR6qYoU+c0PtYe2Qwpv6YaeUw2MqI5RwIr5h2M3xDJQZU4xJv+UYJ
GDjCoMXb4vQYsFtSJaRmcL6qnosVoB9crI9zBU4AbnMqVI1SDcHByrMkELl9Xf2O
4M7mqv00dtDHmIeVWFSwnfJAP44UiVSjIUZCeO7B1lNx3AKnXzH84dMGSHQpXWth
4oBiYrdnonW0ArIShjujI8aiY1ABrRM9Y0YgfLWEmHkXO5Vit8TJTo9hX8OYMUOr
iH7nDXUrQ3l91brTfHcV/lwkBOGPufQbsCay/Bud+1mUDXNUERWHG8q0chxrXiaC
Iva6xKRSPrg013deXHpfuzCu7vt688Js+4VBkGtBjPzrgygOxIsTJslTZ3A+I+lY
YeG6814Yajign0Jh1QDyyPTN4sij4LiDmohYnwbjGOg8Jb+bxKKn+qvS2cNeLo3p
sb+IShHVrrZckmXx9CFvu60Rmd3dx40OwdGffcGkGyZbvHOKMuBs4qhnMent3Pmy
JZqD+VjFTTjZ8fBcd+zWdZhLKB/6Hzzx8JmpP1B46hZ7jfJR+fDOZGL09LZU1dHV
TvG0OtqOojz661E1b0XmCORm6zjn0GZ115H1p7PfdCjsq4792YVnjKpfYtqD9w9p
RKupRDRRe9/USXXRmh7jWeqGTDhJgjpQ/+QUUHNV41CdUEwn49qKzHwFTdLmOa3e
Mh1yaQo8D5R2sSA0ofCzfI/wt9lu/UknWgzP8tg2c7wADc4AA1fHq3VSYvyV8j0T
1ie3CoHyL7xQauou8UPuV/ySHp6FzuIcp7U54xE8nB65eIEYhqnHobRWGplUCPME
nZgOujwgvMEpOyVe06rvU3A38OBnGFo9c4uJEP8RVQaEBjhgrLWZawzV3GNtWHyl
V/F5MgyHMCj8yR7MhTmDshaWuQ9mKqhBg16r1MoFAX2ehNtjzf4zhsO4+DHy97pl
yofNN4O7+BRe1m5zL4sWKGixy0eag5WBJr43yH4QsFH0eYplBIzNfImHQLGyyKi9
oZ6EBFTk3+4j2hCcgjzCLw1r1M7CkRQBhkNJUqvVKxr41RaAmcwxseZynF3TiT2X
gzb63HIJfNh9a4rDfssnrdEtdAKHz0p5lq0y/KXFwYy93diX+H6qVnAmAFyHZoG7
qNbacJz3pFCQuWt2zdYy0VdmkJi8bmghCBXkDxvDzPGUcZ2dumJRUgbp+TM65d+v
/9882vZf2FnhZDDNg9kVsNBE3W2KNIy463E0Qs6LNkQ+8hpWVl8DM5T0dYSRmOdO
IgpWvRUpH4pkbJV/T6wkv18wEvkpsTVOlV3ut6ybADnpU7EcbNFMm+9wJTTKz+jq
059UIHT7WDM370zsUPwkLVkOapxu7LZsKaB1Zbv4xioNsoGyq+7T2DM1NwYVSGTR
oEZNqRC2SrDA3RxAo9P2fVqsLW7le99Lu7tfbUiovz90gltZktrGND2vbQE5Mgb1
96dxAc4geNeNwlnFuN/qbBNBtQRcp9e3jpiPeGTyqeWE20j0IYaDSMOwq8UrPCOn
SnbD57m8qPw/x7L0/teXfioomD0zPmQ+rGK0KQaRxNBnZDrm2PvVByy+OQjs17bQ
kb0lelggFPHjg+ZNkCFMjg25MN8Su1+ogkej06i462R2DUePAp+UzpCmCBMY3OYH
deHjxWzMSfndTxigQ4UCyMOPqe9m6d2AUZ2g0QL8yTA2FJO8+YMZPMNOpGEcTmju
AKlnoT50CBBXoiqI3MVddVerlAWq+/4xeGV9AG2Mv2/uXG6Z5kOGjnlSbYDxgo9t
93omBEmNqg6VHV7Helwr426NIITBjwQlhdaIxQ64ZbDNtOGBLJSVdTAHwYbGpb+k
ZgCOgbnV1OjYvDHxUiu7H6ZJld5YOw1NyRGXBmA1b75XAY44jAa0WhVzTRzGiii4
vfaWTPyS7jGf4rR8Mo48TKJ7Z6aw10aGax1HvQYEqupANTHV1ox/NVylq8D1pxe4
S9GKRoMXNrjIiy86PGuvhBdCGyQwc56B/rb2tzlJB1IMd/1yKr7lE89emWmS4SAh
4EmwMaWvbcoiPx0m0rQi954jcvshGNwXKnFZ9tLPfGr0EROMdpHrXmexJ3ndyg+i
lG2K7MRFxNXqBJ5jCN5PCDuxr1uGIo23bcIbQhxpBjZ6JtgH7HUpufxmFvYnblnC
4RLqZx+8gI9NWVC88axUlq2EEmUG6T03vx9T4u2ek1+fqAnF4HnrIJ1CTmYxwmSi
Uj0ZwGStNrKCn6GGUqbhkj6Cvkf4JUs7AOdcqNoI7ZgoFDUxTOUbmxs16YMcIUW9
Xyi5UNcSB/Nc3jJXRwAWwbmkP5j+jAUBqeEsY+Iu1MEZYbizLwsjgjYHUjMeXRme
BJQRVnJLH7BOnMBo2yKE2CrwVIC8/MOAuZsXg+R4u4pjWh+cVpji9VJD06WfGG39
jXqrlR9ErqGOXKH7Cm5HDuifuf03sKpkjfw5X+AZ8G5H4Hxr2TbkIQ96uh9c6gAU
E8ye65FcE0Mt4LH6XUN64IsoXrOXfaTVd04sWSt0vUAzBFxT+vV/uRHK2LTWetfI
RrgNotvycq43+At6YGFXTbee50P0zZ+EjEqZUIxhbKFutkVfMJ76NWmK0nPFoHPV
cWKf8lO41K+TRMOdzgi9C1dJpGIV3Thpyuk9UxrDfNBAtVUoaaT58LfDWR3P3Rig
y++2/c0OpF/3Mlua0MyvZ/6yiJzXRmyoq2KWEz61/i+ooaHE9dUxHiFpzBkrb87O
telYa7EcqG4xaJE4TSrMWUebfVAokKjmYZx67C9XnAnPyJd2wRcbTLQX0geiLlsu
896w9uRvfBCoQv36O9QEiLkql0RuWORx9GDOKRiGwmaDk26JW9MZe6JWDqmiPWCn
TIuyGViQMa7AomT9vZRX4zzuYmgoQbYsgCpL4CtnnRqVvEg76RNkjUpQLMIk1R6+
hakbgZH2rnZv3kD1GxnO2gKhQICvSDPWCBy9OWgo6UBMHA/9dxm4pyo/7C/PQeOq
aB9bmwfXSpnAR4fPJZOYVO5HyebXpa3KtCILQGh18ubmmZU0RuCrm9jcxNNzcrsr
D2q0F76Bz1SaTdPBexbt2jHweaj4GROGvLJ6Yn1WTlI0RhVIGvsY5bTzcpImsvXi
Kvm58rJUMSSP/4JzRgpFWL7aXGs7IL/+f5uLjMQMM5q5z1mZr7tksF6uzz3do3Qe
eyBurjrc55rgfxg9eC0yAg2pa9KsYczRYMfHrNK39ZSFjNdYFYBQyByEjNR/c1FH
parqU0Jcam8k6nxqJpf+iOuhDVuSj+2Sat0E+8RQKLZCLVpK0p36C0lvjcTis0jK
G5HC8RHXASCKFP0ORz/TG1Un0h3cA3Q/CMKVvxFCixMLV/WYPH7ux9+T+t0KyzL6
SHGw1atWlT/VzigHKW+6TKTokkP/uFYf29PI1N72Kv3hCUgF0UCJuy+YOrLyCR5m
J1gIiaQxX097XE+g0choYiICCknTjZxFoHVKbnTf7J9G5iJcpuBLrybbpG4DV3y6
JU+9Ee805JTGAybVrySDJP2thbCCPg8kkouMnw2O19Vvawm/nQdre2JvBvZAQa/f
K2y7c2VmkS+ZymWxXcGz54sEZUwSuSz6odN/t/mPJHdczM3g7bpoGRu6Jvaj14qP
1ag6cZDDTvw8wMnC8GcXY1D6iHBPz46QtA5ihK0dIRC5da9/KtGCnXa6qzPi0qEQ
TwLBLvwbi9SU+XnnzSoQIp8aauP3Sq0GFts0ndYoy8QCBci6w3IhrBp/xLNGlKrb
2LrdKMB5byGW/B8mUlnaALVoHq4prhaq2OOLAAgWe0panqswmIMXOgGBlseHBkHy
EMmmVBqX8ObC19bDOM8Jlrosq8wF7FUx+a+9c52Td1qnQFDbYwzGBq8Kaz7uzMNK
M3aO6A97eMZxw0TSEXMHHAcKlfVkClPTVaUSweN+rJ27+5mEykF21hBmWgQtxLle
io1LO7U8pKPes9S/UB4NKUAiL//1QprgRCEtbizKT4a2ai1UiNUbimx9Z2FEZBUS
9aBlNkpIVUjnveXU/JbS52IxVy8EazXTSsjMDVvBtsrkVOflqqmlYMlfa5Gq0OkS
DJpafcXbrJGHdAOEBrd5yH2CHr1CJwiUSd3y5GNYXkpwFOF+/xyQp+D5ix24gyQ0
O7nHBQHvUNm2LdufS8y6RFeyb0ABzUJ9KzRC7gr+ErIwiYtf9y8FmQrN29nGfW6u
0Erf/IidO0xkPSjGkpLbLGCEqBJY1PmRkIKMoj0WXtBOpLkUQ//u72gKV9lqhmR9
q+GytZNv1Z540z46Ioei6YL3absW1Mo2IMsR1K851Rx0LsZWWrRUkULNyc1VxUEm
VoR0wYnoFYU7g3NHO6sLFZOCnQ7Z1DxngzLItC3epcXJKL+NaB3+ljcXXLJdGbcu
+chrcfCvB959B+nGFVv6hU/OX/5Nra7gPg/2Rs4cICJ4X8uPvqd4CG46BiJXuH1y
7uzIHUFJF2ZOZB9uutSMHG0fmo2hcsd30Yi0S8x7PU1ndVv8NUoszEVB6txTtOQX
J82VtsTVfrdBCSn6ZJCh4dOGfOlYAswNRpyOaQCk2r7mgIgkWVvpjYsIK3ddchQ9
nTdSuwqidagDa/BmhS+178jZqfNsX9zRja0TEZoAoOKudlGeQRWOZfsyQxHpQ/aY
NB/KuuSzQPQR0GywylBvckVcSIShKH/aNY1yFNaF2vEFnJAoVN28Nrx8rL/vVRfT
PJOLM2Hl7jd358vVmtVCPWCTeF/1ySpLi7ck9/UmlnMnw1f2ZB6zD8QlYMqN11rc
OkTRa1jFWkriu4xb5OAeBRBh+nr0Be6A4rvoAmT75VBvt3qT0PIARTdJXVkJ1Uot
livwQ79j3Jb5gbi9DLO6v4S6XaGsRBIyqr2D36RmZuVNCsTL/1K1P2sI1pRSK8BE
XnBiF2jUlLbkPKL23VslOZSRhEksDt+JZD/dgw6ihqEom1f8byKhiP4Z3Zm5RFdI
dw3/Ii9xDaAl6H/H2y/Ga9vjRbjd99QGxjjvZ8Kkb24wB1aTtTKr+WIGAA2XKLjz
XuwtBj4oPVnEHxu1YdxTdgwGn2vG0cUwaqI1hPVzUH/c1ymbpw2gHlJB+7KmfL78
2L4OeDjQ9IzoFwVWv/fBqRC8jf5JJKLNszIAGhhAc+hrPxKl3a3yHm2BgQSt5Yk7
Lu3ZmrcQAEDp6Oj5qg80ZZLjSnyNIXWB+y4cWuzVgOBR0z5VzZyHKS8YTMHgsaXM
q5LLZV9YtldniQjC9n7RA+lXWZf2gILAbbsqWwEZZ0O4M8r7TDQm1uLxgzYd1nVa
16W+591KjOuZPZBmsabmiyKErRXRb7rw8KMOWT8Mj341RnQASR0bzlobVTL26XsW
qPQ5EgRYXlolT+JZEqX4kEzbaa8JUd7os6iwH1rKhwScAA+0FCJcm2OZhIDgyP1Q
4aWlF8bbSb3/rJEVo0FDZFf6oR80WGE6QAxuVInJ4OAdzivEJedGyai77ejDulVa
1aH68bDRS3W3LlOd6bicE+4FUP1cJ9zk/a4+B/s5xiJSunc/v376B8ELRQpxFaqr
uL2tJJA69YytF/+m6Jyq/L2TVCBFwtSIUxUaDGO82knFanI0WUawNShSYrqw/H5/
nAmM5wmF0gjYBTWnLrpPi/uyisnRshHb+/dMprKH7pUarU36mPXemycZQb3DdTVp
xyZCkOJiTxo/qTNwufzPxUBbDgWbLAVsfAD1R/2uVdnHmxO6K56634Ke1kMy5CnH
ErsK6A45jlIqVOEhM838G/djdCDixJvKBN0HdE7nZx+yvp6yER5Q93JIITXBGp5y
GpgIjM5o834G1pyJwnlUs+X/2IJgUCeHTEWgRn/8XvlYc7B+5DWB/PN9L21MiqTI
hpDI8ezNT3qelPchMknZlzzzN+uktKd7Co5pNwX/2avm5ydxWRuuV/rgRIwWDFVZ
UTnC+rNFPC4QztMI8or9RwWIvzne7msJBqRMGmsZejMzUKcdcFP6CxRPgt3Ubqgu
NbW+ITyE0TgxGcu4ToFy++oBFP3vLj2P+mjKA0aTr3ZYDUygNW1eFYo4b0NluH3O
MMtMrwg6I2Run+FJi8hSuKmPrd42nseuuZDYgjiP+YC2EOJejbi4csfVtYox5/Km
GUt2z3E5S3jKbmHymi7/STtdQAbFHEhKUeQCU0QgrHDm2II2ZKBL6yTyOTWfiik0
92luIWUj8wQL6IKuddYAVfWcZNqhsXvdQenUXjrelMW8qby7dK16FXaIsZ9VjX1M
9k2lLt/b6Lkv0T96FYKnWgIzdrZXXOVzxiWR+MS38jVnIT46gMHtBHXoYwMD4Rdy
pb0hHryIpCaZU4TFa8usmRcNRFROu0SMowTcc8vwnMTJvuu+qQZapknQEn6dEvED
Vah/DU4KbQvURaVOtZNjuFsDgJZ+Nss8div3EcGoHVaWAKQJeMo6yO2Rqd1axS80
KZlwXNcs9gJ0aPnQ0/tHhxTKOFlCrxgPKbWJQ7ZJdjl75SVfr6fL8hjav/9FDt+1
nHx1Dt5MdTn0EVsQxDG5D7uNwIf3yeKKWj9RB0+F2/HmtTesfC4LWvu0GDBTthXD
36hlxRgHrppUJc7nnVhD1JwwM5AplOzH9SgqUznD2cJQGHPOcZPmjgyFFY/srAmS
drMD1qCfAW4Ywy32CnCbjDvGzrdRcojo5LbNxHYpE8Vxrozk5818BPPFvl01FFKa
7bKGZPWvxkfvesbajAs7uhNbHgAxibBs50FFzIxGKFXhtwzLHdNZ1SxZgaG2ffa1
IYl/wwjOTTsHj6uKtFjUpYt9BEi37sAeVgJoKZftf+SRf93Iq9ib9zyLH7oyp2Xf
aJU9E/1FsjBXQYwvQR868T6pFu4MUJTMxjiODZ3te2cCsNhuoXh6rU1eAgg/11fs
sakY/T/tP/aFxhl3TUAC/xvLQF1Zu2O0HutypFEb0LthwT8XpKQmHYqYgpqjx5cQ
LXIXC8E5S9jvdN/9KerI2MyiwqIoQtr1TPz9t1JH9FiaYQYvJqoflOCSupmbz0QZ
oBWZwclTPlSX52ZUOsIKjZmQTi7pA/a2TTMby3LAWC6Qa4Bhh0HvnEEUH8tjrIO7
SnHQD4JmhE1MYbfqMpoTxGr90rX5L7Syt/20azVH0cQBjOnhZUPCvll5+GD8iSkc
x0/EJoEYCwT2K9JMF28o5Vh1bz2dAADlWqG+BYt+3diJuxlFBI5+oSC3+JWjA90u
R5za4ouDsIV+QTKjGF6iyWA94biA5GGfFuOok6sl2inVAy9mgAkhY9nq9RazeihH
VpQ/ZQZtWsF3NTMKSF+3px1Z5t3IYG9EB85i9ffdVA8F97tHm1zRXdmUVU4GeQSI
3dABCcz1ATJVwWwo1WAtPT/zaGVFKwtGgn1eBM0ZNz67BgdPgIVY4z+aICCJLx3t
gKbwQ3wMfmw/4kBX6XIU3HDRLVPSPnIfin/DbPz8mSE9WQBSEp6xOe8DmtJPoE8b
0TMMpsNf0zpOKpjL7xo+8ZJOEHcm9djZDRiJgxt0qNzfEOJJjWndmt45m11xHH+8
kOdx2TXMNISSAVDEJI/uZP0XKdpjMI+tZP67TFXA7pDdDgKj5enM/SZki/gQ9G8I
00DpvC/DYAn+muKx6CcYIuSK8xQ3rnB9SxGVLjbvPCem0eAsLOMbhuAtWGKhtAeH
xHm9lXS1MwgUC8ch9ay+8FYN+RAFr0fwKcq6hQEcrgXOOdIidPEASXHqZYajq245
a5W+O1C8bktIj9yS0lbQYnbY25xlYx7zZeVjQMHyEZ6PnAM7a/Mi6eVviBN7D0MA
RblfgK8hunar0X1yGT3w3axHBLcVoFSS+pDW+qqsMItHxplm8kBF7Q5+qAtMB729
elZDG1dGT3HCruscT/KOGHNvYz8m9Na8Ku0HqqZW2F6GQzp4r/e2n/k2oHcGQiQC
rSYvTZ2rdVdDhuWtYEJX1QL7wm4Eea/ZDG9ZlEPt0YrQZVJGAs49+X8/MuLl92XW
Aq7BOPaHsP7VbhDIHL3rntPIwIWspehMmLbtpXeV/sH2WluF0whHqw7Lq1pFCh2V
b6jWqIUVYOoCfFyqeYdw3XA/18dtcehkWlHOnP/u38ftw5nO8lMutmBz2y8/YpJ4
TLmEcscw0KqEAgtjyZn1nrO+PDA5yjOs9nt5Fhy7HKiQkr7+XhfeOAi4+rHoEaej
JTfCNn/b/MZfFPY6FI3RqcrPW1+monmBX3LvidJg4WrrUhssdXXJYk5mATzGEg02
EOuBQNd/wlQeiGz5sHfg/Q0c13taG0Ftut1Ik/lW+iapTBMMurDUZ0Wf75QbItUF
+zRBYgizn4t10hTEOd8XQ9x0NDGm1iXj/9wfxydw8e5At3Xty/fDroJv6ij414ik
QGN6vJSqRhD3ElDCzUqQmo7yhg3A+v/r1nTTdHS3RGqpDF8DVPo29nAcFvglQhwi
CApaZEb60HSakI9K1iArMSmdhsc8GQtGng2rQzEkL5vlyFLT1BBxbyEmgtS9XmYJ
7sOJOTHTLONyQYG79TC2gQYAetktjlk42bYCQXak99XYZ0j+14FwpoRmQH520pHz
swGpqyQ4nbP4Vpzm3vb9fO3EYe5CK+Lb0IP3Xq1oppIf69j+7MNGtxx7okWR83dd
TFnPOYs49/p81xFwaunRFQ==
`pragma protect end_protected
