`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Ag86Ahw/ENdVrIZHmSjI89Ur/tyqZ8ESTyHZ3bvtKb7MlAzOVGvmeKPD7JFMa4vl
dXm8qefd/I49YJRJFRbLNMbJ6EjIacsqsX2jR8dWvuxB2JZvWqS8EshJm8Qy6+PY
8YTejr240MejskldETqspawWpKGlDkAoH/sZpsu1ptE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 11360), data_block
gkk9VBeSMJ1iUkoqIXXXGTNKfTIQ9wQpxzkoMWeWIY7rIR507/JKcDD/tsSpCx4S
ZnIjsOKqswjcw1iPjmkUAW/Ghj3tGmaaLmIr404BuTY4jiTcngA5NHccJaq9p6P2
8KXVdIFpoHTF1HrT2B1zCKESJVlpul7K9dOMTgGfaAnya8ffGwJqDrvBbSerw3fm
Rp2IhiNTggJll68xME7HidLhOLAVxd/sI8b0MQ/74CyNb0aR1d3XAd1Kj4JQIK7n
Hf3WTXvdQsJrsaPt6c5L9kqnAPBsmEK4j4i+YbJovRTRw/55az9Ea8RO5c98ozMg
3VO6HV9VrW/5sez977lQGs28T885twa1k6HoVhiiTZdgDt7IfR4rfUsaRumGHL9k
4d96w1ZrlAha0bqhuW7VjBoNNgpNaPulL9lGfPVa2xTt0VuKSTMadmMLIVVcpnw2
dIs1GF51IecnlJx3MTh3yXha+pUKwrdUV6hFbG+AE4zlpukbbdKeqWqxMS6gfY/M
UQrd6SRckhGtsJMsc2XY/78lx+NMBirWdMEvSaVmmcGS6DY/jpH00MSNlNpML9Qd
tMc+IQrqWE5Bfcr89Bet9r5OZ/WOZ4tmfLycgjgsr5l4l0D8ojmiKVWUOz7UKsNj
Jh1s4UHNZ+8RbmxZJ0X5htPLT4tW/i8llpXTPLedghfNtS/gPPjt1RcTY1+aVo/9
y4GUI1RtKtJTi7QyuGW2UjX3DbgSdpoalQLrPNzHyYNRQOYaeoPu1iX+Vw3JhvC2
rKMCZ1Svg8JPvoOl24qy/gsw08i8QQFM9V+Hw47JUlVlLRUqQGPiN3vOE4ofuNLU
uotODw/YvqiuGSpNNf0i44I3a1p9E6b+nL0yOCGt/inzQozTPuHBnyaoPiqg7uCw
yFwlCm/E1XOn4wnYHot7roazXEDk6v2NMHbYQC6mi5I/u/HL+vIjDEJ2f1Ku6ZhQ
Q79j+EkAVdl7GVCi3H3VZkZYfFTiPQrInejrV2Seo70Zl2Fl1XVaLOSfpTO8aKZ/
SZYKuU9gcqbGdPQlahLgSZKMV6OF6dQcVwfgyS2gAnSgU/MXPMVhJfSYOLFvzkyH
AUK9tUEfdx8zzzq1/K4NSLt54S/e7IDOueiEwkRnBvN0DYzyos6ibpU2HDTM+7ww
Rm3CdkncQF7km1J30QJxMyTKF/bQvmbVPz4AlNw5m2+6iVHe9KGXFpBF/E36/Ars
Kkzm7OneohgIbnYxt32ouBakuHglLtgtZEbPo/YBP+fCmb9nSyQLyEoGy6vb7hel
TED31VV+iuue/qRlLp/IsRekXjKE02RAIolCiYn49NYa4jrNvxU91euvveqo7Hfq
JHh1DRk2E3K6BwbNbsaWzsS/0XGgk1XXiN0C9CRIeDn2KiatAVvkXAlHojiRUiHF
JD4blhX5xp72pysufjATMif0M5ZhSyJbASA5ns1dQDbF0PR1itJ9OTMSyzCHyRX7
5BfYoOv+MN9pBHJxdbLaZRyDvHe0v8mLbQ37p+j/x93EsS8hJkmpp2i4SQRp1IBe
IioMcBAcluSxJ+RpE0WochTh35vpPi7cLBSQnDbiKu8/6SymVbSK05OEqgiROuIm
ildjY1ZCpDOPpSH3le7HzNMk5sDneH2aLAV36h0PKE64uhoVT4x23kc/kYBFVdjk
q6U0QudbiRapgpJ/lM8PjcXet66aTHDTYBF9ooQPnhtcbTfFG7ZPn22E6w3ITkpD
HYd+Z77ZD+J72e4lPKsvabJRNpcqAmvr5ocUlxppAhF/DfiuWtf9bEQIj6d/hrP3
lR71kfYoos6oIs2Dc3l0d2Nt4m/exRDGlITtmXdMXpBGtO4/6GjM5B/1LtkpgtFW
7GY025jr5ITVF8NZVcaWiTwHGOjfwTsKS5VWzvA2XuERNtcpKVS4AG3NyaWq+1rU
8MSmcAX6euqdQ3CLqcrXQJgqNVEIKcgwpTgDQ6okXHYjYpBOx/W1A4vWgZmk9Q6L
xVOwYCWu3uCmhaDH+plPodnIcm50YSC9Zr+cWwymIl9cvlPt4oahDpUlLZgVputg
h9APETpvKEoyuHCSsin2Gnqcgl85n9/YA16vzRiy0LUPQ2DANGrrdMQxGig+Nsd9
bUuTdY4EGkHY7kjfir2e0DyMzWikkJ0IGYazk7yXp9stq2ZY85tzO/eVquKZIbpj
YgXy0TAFKCebdtWLuJw9BkIL88txecvxhHELLrkz/13QAYShM2fiC3m8v+GqlP2o
v9XdC8uv6YPR7mQ4FAYA0MticD44V/3YQtyeDsIUg4PD3I7BOHQIUPSHenf0SRA4
RxHX8u5O45D/RkShbxfLTc7PUcEAb+jBQojnofH8BeW6XSLe1Fw4fjB9KbothMCO
XzVb0V3oovUnGIiRjURypmqg7C94Kvbh7Q2L5ZvvOYCo+BGE1KQlmRLxU2aVnmjc
9fmAWpCOxZF0SV9+ESY1ALMKde571BD1pEnDmsOwkMXYe+XiKR6uxygRVN68ihn/
duVtiJNvvt+AG9eLnltuztvfkakrS5JUG4X2PYXnyrNMiOcoS3rhkKCu7PPtyw/V
KM1nRsO0ov0HQ5JR7E8SrDnaa5PyE+Qrvz7U7Q9afelJTrwSgnP5EiZCfcQJqoeh
EbBE9RCmJeAKx+0KhukG76gBK+86x9BkBvGARHGe0IJACmiTPu2W/C+wMtXEXwdb
JqjMUqEwxtBmZL0oH3FKLVWeDBYEPbDRdEAByjpEpJBqM+pVBuBpyMtxqKA5+qDd
2C1/Nwafp6k5WfKI0JcUPK1+wIn/7X1AiSVkghIM8ekbr7dAZIy9CXaoDZQv4seB
Zyn8vSTq+oXI6PNOaKC7DcgZQv4LloMgqXYiVSQjm6m+1t6noTqjURFT5zY5YkFc
aJWFcWPJ45bL4Xd+wynG0x6CT1VWliawIzSlzPfu7wp3isp9MG+a87irxhnp9/z8
EHyuIuPAgrgVZ2SXyDEOu7Bd36tkJ5UywrGgDJE8wlrpPxcwZLWlps4FoFT37QZS
wvsF8IMVQxy0UmD074UVPpz1/LmylyXEzNSKIH4p1+FoerJcfCw+6NdsI3sWSsKN
c2cFESkyvybhajGjQjYjPe7qw9JAhGMr4coxnYARU/f5NDYcNzOfmyPy+7CKLmt5
xT1B+BiTQ3zXUXq3R2Uonh18M/ws8CNR+sZqG7chzhvyRxsOcrz9FCCZA7vb9Bfg
nVlroUa6hueUiedhk1phQ2cvL0ZtY4ZqDuHO5QU74lLUKbLQwXjyGEHnvmd9hihd
c/BBYLM3mTjwcDT2bjG5kJTumLmSqLC6mihqQ2UvZwqP8FjbFTP3w1zAM7HjougT
TnIu8xtJTT1g4JXBhS3xeWsi7i1SQfc3l1yGk2rhTHIDoLf3ttdgCzGFJV2UaG1F
qM52xPEsmTMKEUOb+XfG/It0ata38pleKZKH34TX0JLCTzVj2nlisMVyF4++YvUk
mZb7lwsmwhNGose8MMrCT6xPkWMhoAFayNsRwvEmlJrU+1V3smHXKu+xUxFn9Inn
ThDpQjuiae0tP5GCVr/zZ+KFU/yJShCNnvqE/uTgRZ+iMwsk4qG2H6G8F2ky+4ED
I4TKyGe3aDpQQ27I0P3S7GrjvsN6XkuKttIqEu0NbAYKiL+7HSZlSgK9PAJfs8I6
HtER2qVGclculHT3JanFwL7MaFrfHE2ACW3biBUuYyzQRxTDGqjacH5ptl7wovov
M92dA7obcmlVRYNLcUs44wXz/D7MO2NM2sfXRC+fpk+wYzAlCgTgxv/y4QF217vx
HtvxsGNrbpGry6UtXTT9obh+j2DVmVpILYScs7BVvBid8ZfgsYECZswP5hgO7nXp
5et4yeyeW12CgZav4cv/adV0yjCySiNsLqSTCUNv647cDMo1NkoiZoEcc+KpKVcc
9slOPzwheufxcdkHogE4it2WoywZwKYGsJU/dtX1ivbw94Q6yYFqyHid63fBuFPX
y534Ms8vVZGhNPyqlOnHGvaevXWmALWSLfUs1k7xJpfzu9zlt5cQB7bZCEmjsYAn
6mZU6O6w2wY6MzcG/oVdjoAKYB2XRgxujXcspK0X2auSb05NTTatfeI7FDxFGwv6
ik66an/Sk+uymBo7btUD06qQh0ScCnGLcBUlLVm55kbcdBDTmC194n3Deqqjlb97
nJvqiPesVTCwLMz9BNzVePmE9efThORjP3xSoA2RnFYVVrPe1Uh/C5HTFl0GTfos
5PMbSwI0gKPrUYvsZb7WHz5FM+mqKey55Nk3SsTwGH9vf8RKJZTHJT37oiceVHTn
fvmLUr6wLA3uqiWXid6MK3xYpouUR0i/AwKzVs+SCieILwseRVHtFOaLXqXAhysk
jM4e6Qqadmhv+GWn2ipnKaUPN6H7+/si1bqtSsFKfn2sbT+m0JOrg5p/ynEm9wTx
ucGTYPvXWOVZ3pthVfEr1tmkW6GvdTJSFPOigtRbYbSpKvY3h6sK5JsysS22SX7Y
fxk1JPHErkb5EHC1eQE9ofGjk3mmPBSdG2ORJUJvbsbEvQeGMw6lYymS1ZkigE+7
tkqYBfordWXEtH7ivIbWtVn/B/zWBzkMFtCH0ffEMUn3Sj0DeDd0LFquD/23Lo0L
mdhOWabZrmCjyUVbAcm2OtdXCZwJWPQG58BEixmOZTl+4hRVbfgBVoQglpiGlVLh
9MQbYxu7Mt1kkJ3TfTonhIzOSsAeL23+raXRyWyGPuVIBgygGnHyBWh3JM7CSkt3
mGlHLL/qE8Z6vy5+LJYhD84v6xId0Hk/Zf669SslUwmFbvPrhW9AoSk95MfUoy5W
86Snmk8ATq0/4R5hNwSBe5aFI3CodjY9o//F9/qYgIhaG7h8aQ7smF1v/DVutii8
JhgetVnLkwEW4q9AzQ7T8dzsDdqSwXJZRlfTPMlx8RA12DMbheOvDDgdKRuPJHsg
XERoX97ieGti0auwoSkEGYw+V8rM9BAF8dj+5xXfz61xXdYZJC6prH+DAGGzIcgO
UYhv7HYyhFCEbX051l+its1KDU2He2RUsXlOfDFWfzI19r8GGlgFtP5CPiOGOkfZ
jSqS28v674s6k6EvtI8Dsvj/GNkNlIzkUCUe3XQy6Z0zh6jwsJI1potpmtmpSdxp
eSe8mL6jVsBmh/htpEbwLkLvcgeEvrsGGjxFu7Xehj4xMbnGtEl9h8J1M76nKOfF
86qkltv/2Mp9p5z+wTJc9IwLc81fakub32+BGiardudsnv3+jlvGTb6bsDk5kD1j
yOPqSHqsoJeF7kha0CJF5piozla6L+oy06SnXhRmVGfTACXmzGxVmnDEQ1TalaQU
JG40DJnpCwSl6cD1Uwe/CiNwodJ/YGf+v+oMErmw14kC6uK0VPrX5ywDfBRacEx6
27AYPKnOxsT1oqEZEQ7zY053ItXHeJj3V1a1jRmqqk4cK0EjBx30/WkZnVAvaxrO
Lz/EnlITQUruNRWdR7LcekdeSBnfq5KwtOj/t4FcNBUhNdC2qHTuMY0OC6KmRkVK
+EWE0mtk7OGksvOSl9M0EMTol00vL7qsEqO25LOXcLFFlCWufEuUtJ+V2MgpPLhJ
d18l5yvEF4W6lrdbcs10oo7dbv2zb8a/Pf+w14UoL8G3dkxJmEUFjRgCv3SBKBZy
ZlAMRnU8xaQjmbq2x4VJ5lfYTc4T7RYuo2ILh6X140KB0PjhrBumVfLJi/blKCUv
XsQtT/fvxRT+Y8+xiC6sw7Mt1ZhhyR7ag0b+VfagoGWzAlFarLYjNP5ut58hN8u6
65+RAMqPxFqEb7+YI5R2RK13q897vXwHOhAKGIKq6+9WuBF45szkeC8OQo4fkMTr
74JIm4RGVrOWFwV/t/eWgIwRAlwQ0Kuj516n7pYUR/54tPW2u+AggueR3R4ZyHyd
5mGN1JDkrupxVf9asJ0ZPuIdLFxpfWXEgTHUKumLmWvePNYP88149n844ykBHGL3
fbHrsh2ckl8bC5+F4HQxdBD6WBkkhlmCOZ9deSCDEKOGS3GwawSYNUd2+yJOSr1n
PjOGRZcOhxJJF4dQAjzyFwSg204UUZoS+YKcE1MCZeinG6RJcoV9gUepRrLsUeb8
VKtH3XVTuN/t+NHBderEosaG3EJDMCHkfPSxVObngUiix9XIEervcO+ISq8a/+Su
IJ2ARGAAhmRaMMjP4AW5X9VR5rAesrFUjP0Z4Xqx5O1kD4wSo8Ox5HcUy0QV7Lsm
K4G0B2VY8rSWinxyqKABtpgWCmm3oCNtlYWmFGiJbAoD26ReURpnyEahHv8ZozZZ
v97MyIVtXNUxxrXo3JFC4cbXgBvlIyHRA7KsyWZf90wzg6hawoPqpE+JG9Ai+ap6
42Iq+LxkM1fPY/fvng8ddYBNlu68oF++wKr0/xrGkCaQqkSxTmKjDn2v5SoLBs47
DaECyX64dNxWq35B6/91oB5vKnDm1A/r00Y7gAFznNa8WPM7kEMT1OfMZ4k+xPGh
Q/+fWE5wrHh4ULINXgQ05u3WY2e2OEz1i7Xu6tPiBtg7fD5x4m4fYxurfUZltJyR
Da2XDHe2jzea96Hrdx3uS54wA3+Lh81Esm6n7zSzuNbIL7tpdT1UGQ1bBdj+caoR
8RU4xey8uExL6Z1hgzZGGpQBGuvWN2tT5EyL5f9HiRH7UP+FgDAk3Mbh0EV0KVOP
JKOGSqdM/3VqK1N35Zsj0bhztqBU0EBSAmQv563RtPzZ42pkwGtkJLMLURVj9tqd
7iq3EKmMyX/5WZJim/kLPeYiaWIZDiwrtXZ17ozofKza8eB2fwUV2NlYyhYmTpZy
0z2E9GWGOg+XiIfiZxid7e2IJljn2OfDOKIIzgrwxApW1+HWnCxcA0Px9cRkE5C7
03O10dWqzSokDy1Cfc+i+XWyXSczcInVSrV4fs6tzBknFHKH0nvZrhhkzH3NWdnB
qKSd1s+Si1xMWcMZnRPitjOnYc6ZytwueLDbIwHRkHTJVzGKNEmsRERnVBOg3qg5
eM0qehzCDHlJ7bQ9tKKxBZRGP9etPZ49XMLYGosYWyZL/caK/muqvX/XnW8Sviod
kOvkqxMjCti4PEZdf9YNGiqWSa8GnH3vXcOxcONnjnt4UlBYnsXtBpXubNEBm2f2
OWk9Rs8RsCN9HoKxFsAyS/XACUWscsFIhGhe6Fjy1xE5r2um6TZNpqUYUB6F3NkG
k8yR9XY+Xw+tYMZDmlD7OgmJhO/FVIZZR9BC8oGCTb2zZhOQmuCsymI/1AANEb1l
3fg1WEyfmCLFABYvCxGR3N1KLhsiybhdJfAETfUtFPLDfj/obGXk4w/kNQJSMDaA
r4ArK17gkoOK7IHYrWj2eLLMnCrnUvTqwJqE1qv8ws2CJjuZUJLzQrNUcX1FY02y
FiUT+2xhUff9JiJFR2fcSZ8QMqWmfl7pqKjOwDKK2fK36hTBjJCqHdmhKozh3gXe
tQKJB0cYNnm8OjvjVzNJ8xl+vyZN6LdhwKDfQqJw3Wi5jfRnvvlzPgglPaA8+W40
BDnsvfQ35+np4J/++ndfQp1ueuOukL+Dkio3CnzjMO/dnET8t5/MEuSYfylG7GvB
D++zwTRhONChSdad2JkDTANG0wJJY332NksVAcyrjERGmThxl1efK6aobrsLUXbq
jyG0HLMeFLaWlc9JTeYzLjiyVrjcLQdFlNTqLxohldzJU2v5UWnq8faznnlkFjoT
7DOra3XS+OHkqoU0wOMMdwUjykgszaQa+PVGRhQhGEYOjzdvvFqDSr1NlpyI73vS
BhPisOvN3vEzAH4K1kH906p8ZKBj4HywF/w3+o5bRd1RQEwWhzkFhaOOmaDhxj1o
xp7W1ycHQlLYnJUNJ/gYa6nD8/iiM+JZuJ40GDkmLonSCuvl/seD+f8kqwZc4qKt
lBCT6YoLlxVCDWWpVv3lOb58golyhoYN63qvLOfo/1kNalT8Nk4G0MJilGN1VfrF
IELobHByixZhRDdDQwUrXfYW85Gi2R+dXSbRjsZ7a8VIuSL3/h8qrM5jxWveDZZP
Up6d9LxGuOaah1spH1aUWpDzuZsBFFmeAf/1vHuXjA+0g+w0ro7f0xe3iDI54UH9
PtmuFFrZ7LAZ56PKsOEGJPwuKw7wC7ZXtle4WstSA8YelZT/OrhqWQKIwNjKGtCk
oUDAXe6ih9LCjKxZMHf5hHbdwa5cOyi3JCAa+tEaVlZfDl0/N4KiQ50PcAlQwQ1F
D9YD7t1KGcjNTEKu1+S5v1DBuY6Jxyzzm0vPBX0ApX4gBtrwLbIzkxDi1mExOzlF
ZyZsI76iaBoU6DhdO2i/utwgq3i1TbBnbFZD/8GcK85Ods1cj1GLunWv7lBNiNxT
rD/QdwoTUiwN8gucrUeDHc8tL9ktU6I4CNoOEvWuh0jwW4KL23O5rmU5vqRPkmRP
S91kDd6UcUpZ7iqk4hJ9E70V5ShiIM2mXJy8nowwBSbqs8bCXKlQIQStJsAmyy9/
W5u10FwXlbj+ad3acgpGGzJLu/J07gtq2Yp9dsk+WOIfUAc9LBfRwGI2JQGJy0Cb
/078GgTMqibGUZ2SnwAKxeQ3wE7RLJXUtHE/rpvCXcrsTvdrBoiL4M5U0t4jIItF
Fktq5FUbllm87q0IN44NY/aHBRR5ksBbUKzcgUXKnVLLOQDyxrhL/6XSdM918lXv
300F0mysndmAGzukCL1MQe5bmgmQw9jqd8ps2j/mxHMtLrMoKJ/1Rqs80WhEr2MK
nvMrbYXwOTl3jxiIK+ut5HK78DXoMPjj9yrcNFpHr52D9QqKsdIF1pzQCgD7+HG4
tbqQjt9aVxHYNqtVKgrny7C6W0oUllHIA1DbyNWKdaam8MXyifWlPfqAURTXAzVL
N6AWjMqvbq6Lt+zAVA23ZHFKfAhsJThzbHH4tXNWr13O5tdReXcHh8v19Hk33xrM
Krcn32cr+73y0P79CTAoukt6Z7wHqJJ8ueXx2pSEEZqBvBKYoLi1iocxlUYId3tY
/EUjQepXIUOoP6CKhvG6wLZyR0R7io+Ds0iaWLUMmmB44Gl1O3LVUsxEdaLJLRKN
ViRWhyvL96c+nHEi1D2ZAqMhg5jA+X27dcqPLgs4dSk7cF/29GFC6y0wGeBCE7h9
qAAlzgXCpwBU4PT5RskFG0deEbPNngj4PbZs1Kzk7C2CZhF6Er+IzBihrhrExeiN
qXtnRAqNNP3BkVxUydAFP3sNBJ7bAKnN1KOwdi96Nl18xmXEgKiOsjUUjTaZxd9A
TKCDwW3ECFo04ta2GR4D64A7uCzxUJM2j954z5/p1/64ixSn5Rm6oH16dOtRepRy
JEuE5vZbwkrI1Hhsyhliz7yJoKKxsnccvQnXv+X2zhzsSl7i9d977FjNFVcwgvyP
lJGk9FN+0A7tCJqTZChnqtWlV8VMjLmGs3nKmjuShah6fOfEAmqS2kYMWbcBCqlH
oVzl8XPmRtI8BiiJfGBV6o4pjyGaz5pVRWct48sF67ps3josUyOFG+EJudX0iKEk
VnBw4cbfxaKBa6tRFI+D6RMX635M8qOW7v64cgN3K+Zv+PwU1U9PF20bwPTpXHeD
pPmA34HS3Ib9PGIjCvQcRkgAcPGNhzrK9+Iw9L5BY/iwDvMhbRuLZPwbIE+XyyMz
UXojvqwdPE6ZhkvLmug8OU5mIi0nsB44W1QXEmzAxZlPSJoGba4n2vxdp1iIiJAO
fO+ozfcm9SV3FzuMI0ai28/s864IyFbFawcZfR3uzfoVw8cxCU2s2zXsgOJBka2y
M/OnB19kCfGChTtfQ3OlrJ7aeMwRKeuUWSZA3kNqGn1Wso9jV79QKMGBRFew12N0
HOLHFcVTqjLbRWoUUrt/VXlkC6jQOplPVY5vAy0wk9EcXh2KQ3/yRAmL1lHJpcre
qSGDp07YPh6KqjzjvpyH73yNYVMeKZ1Q5+KZBsCn09RzyG4IbU13IA00UVUImbAc
FyGQYUyyy1eBwisPhVQfvd85A6IZldKKcOFxbOvRW54UCkby2cRCK7gX9UPCd5T6
wM3fxA6suZ+WwfrUoDL35WAVTt0x6faEpefhKdXDq6mixvIYAKki/mTcT5IY/yb3
GZ7cZ8L33bBgbuYU6QFmfR2F3tSmO1n9fdW68O0OrZUIrKWMdxmf+D43P96aofrg
jQZLs/c/Vh2K1EBI1W+CK/li/rDXLadaitCuuyEKpUitxBOvM7zZf/y5xzfgRuU5
RIEn40yGySeZsUlTueUhNSG+Ff3vF0G7h3JjWM26OtvZJQ1jYyu/z88Wb8hXq9Ef
E8dyNg2kjDZ5I6vf3W3ASRIEBGo+ZqrWAbl8Bbe07saMxg6omcoAaAVs9z5q92tT
IAFIuF2dmJGzGKfj2kCPxNeYDiBFzwo4Kiof9kycTpYJ8S2QzPaXH1IqAHQsWbs7
PXbl7amGDswNI2g+BioOqftkn6Z+1ZUL/c11MJkMjxt/KAJJBVkCzgxBrz4iRvd3
eUcpQnXY4eRb5PerNkD4scly9tFew7VbHtytOgy8VGHFuf+NZ5RiOcWYL7ApoUeZ
3UyJSPIRlKDnjDI9IFZOMpIjok617dGLpjpuWUYDHptdFhBqAaq6NePIxtOVoul+
i8OA4bP9NHr/EeErInz37ZjPWBvKbFiNLhD1ZrGZSrZ1IOtG59WkfStHwfncKodP
3kzEZ3Nl05EV00G2ykzXRugW5WeBOf14KgIb/MAqxIdCsXMfdozJhFBOfsS5LfCW
WOGsSQQvQISGk0fskYeCLhiadZD4Mm3KEG7/pkxXOsPFz3dQ32AEQqqQA/VoRWcz
VqFOh61rMFSyS87KLFyGHPCB3LELE3B/qrYOq/tkq+R3i/+FJVnAPiOIz1wvGlID
XFMK38fse+3aly7pooAHAPmWu3IRIXFoZrrbBKqnOYE88I1/YZndOcFtjJKwHjgP
pFbOoIbtcyZ/Zsx5CxwIe3XvYUOyuv2C0VjVgsvVJzoHnSCfdZ/NFb8oqtKAmle0
Uu3rPy/EfT2Lk0PXDfP7hMt/9AZAH6x8isxFLnjW9+FXpjcO6a5qOGJtT1xIMvqh
RlVy0rv+UeE5FiFPlx5SNEXMGEqRbZt2CjZY/hBTp22Q4Ge4kUtYmxfHC9GWFpth
2nS3P63NG623OnlhL10iH/Xx9ZRehS0Yoe80GrLLzqj2toTRpv3j9hECL6hkGGjG
Z5DVGJ4mm2dxZ3iZ9Cm6LlTOZ4SJ4MTR02WG7uSTmnK2SwS7LLXsoYSHgJhr2QC4
PiNzVivbatFZxDX7J5atLBUe8wC+cXWO04QYpNcztMU/RJMH7geq9rDGnL7eGXcY
B/wIkMHCHd+4L7DazzbG03/OuSjor+diMjyf8uPTIjX3+qEjygdHuwSgPJWpM84o
2p2YyZRb4X8/AHhjG/0/74C6GKK9+JNeMzIGiE4hNe1rK88nMJkZLVuU5XFbpaSb
7hnul36xeRcdCJxHNV6tNJggicve/2wfGR0V3n0ANmAy3s2LlKVT4ISPZl5z3uM7
ORenQm7Kp1lTZn2RcTd+Ev/eNvKj0r+2nRLtA7lMbyaPMF/blYJ12vZpcWNEE/Xo
yxD3r27x7F7jVV9et4oli8K0vjvn/Xzr1+yk7sDLd7DLB5wZob0MjQ6ZAfQd/csP
zM2h4OEtXoM/dcYNzzD54c8RQS+b7SM7gAj2X3kxmQzwjRn0eedEf+p7nDueMBSd
lqABUocohq7VkSWAtgyDpFUlKgORqd1NXvKiEfIt7t9+tDYaNUU5uUhYL//8YOgv
6M27nFXPlA4olWMnuNnLm008Uo8f9/h1apo29TL683jJeDIaJhQuiFUM8nSpCQVI
/OSVtpKbZ2ReCUkztZ6/cCmYMT09ynkIzVFu9+uAA7H6z9wMwXeN0i+w4H4VF6u4
bufciRGuUt6sGXhkRmniUQIwBEzf27ZJkcenDQK3RbqffudxhY7wERlNcetDMEE4
ML7BiRQhDoNkb9m1F7k2XBDYyB0tHZGsw3QM7+pB10r75vvMJcQJI1rH4Mj81auB
pLrL3NFzFR76AydK8CXvyt1idOappfglDx/UvJTsJbYMwjOe2GbJemeL9WPCBbZw
ensd61/0IAG/1oDD24Y4HXPPQ+c71z1zEV9n262wh+lbBwk+Pi+atSDn3+a/tGPo
kar2S7BAVgBsEeJ0GLYfCnJPaHJBrd3gmyb2qOjK5u44/mHNS748RxurudCgdzbG
JH1qOMpw23Idk3qD+0/fO/b+sCsT1s/UUtGh18+Hyiek/35gK1P8hwcYtS25BFmW
Q5WSZo+TolPF4rEHMaCOdoTUKNdMXwcBs9ePeMmiybRTb15EwAsAvbKh2zN3aN7x
tjNCNfP8c5PVz/YdycaDrkG/h3eKSikOiDQlmaFAHEOZwAQM2uU3I1cOIORJIcFq
pB+HBGT6TGIqj8fAgOfH09r9UJccPJ9Fp50VdWn2sqEAJtMltPElRhm4KhHsirpV
xYv2YAU3uV4dJ99EAt9DuxPbD8J2q6idNKFLe9wST6uF/PPEMayrdDUA7caHc6ll
Nrck5zrTdvTCcHjlz6g3WvBwsdYxPpZ4M4weur7omRqij2sYKSYf0uuQfORcrFnb
UZWW468yNjka9F+42W2wjD2BlwU3NTqDkKN8x+nB+VLsMvez67hD8kqL/B5u8m2T
D7QxZ7WB2D6LDa6Z7KdqLE9ydBftbsrB7G3d1xu60uz5cLWAEqAdYw53DDQ9+6z9
t2VTx5YpUt+dDKu+6dr7My7TTwFx9L5HXmzOxiU4yOuy46/nIlNVeZvQDpuDZ+jy
JaSLy/JSqmiD1yikuzgS2f5/AUE1J59CEpISZ5F+qrJwXjipABXlEqeQcigLF+4Y
Jvl3D/kADHuAvaYQCw8hKTcWwuBstMxr6BQP9i1m2JlbojMWrMSmetB5BIdph+in
cMYdkf7oN9eqbyWFMEQp7O3Yk4AVg04Xlhia1mRX+64bY/ePzsrHtSM9GJv8KCiE
1+bbnSywKVUVkMEmlXfVk4/E7I7ICvS25+wslXFrgBmNF+nMcFfucXVX8HKfh93X
WO1LbOH+y3Z/yyck834+y5sqbOLi9jNrhlmjeFgc0YNPxLO/Ixi2YvF9Bd6/rjM2
pmqnUaul0g+9h5dkLYnfhRMHEkyBa2J5ExQ1rqjkagaX/sfD9XQoq+HdYxa/m8BZ
r4GpN26NbZwrTcqNSsv7T4jJPcW9soA04hClfsnw0xBPKX8Ke4r82E7+/j7ABqWW
kzWD6IwaRWoB3QIY/B0H+WUqJBHxSk44EQewENUC3ZYQsoVcDwlkx9/Xkn1qcre5
I66n8t0WyvNNVGv9rAZ/tBz9fH1lrCwb9rQdxTbcmUxTFu7gnH5Pn4t0CoBuSp8r
GtssUC7189tfazv0xkppnlPwEZE01EQ1LEk7C88H5iqB+KtWbdwvB2325KQIMKaj
HpLfq80FVEqHQqtPY8ivc/+BJGechNT0xOGGHBamdghjNxesC0oowQAwxyya3kM6
l5FAOFLlIhs/F23qzJRRJMC2T3c5jv4ThNlMfS11FjMyKrQgwNAgu2kgkYyqf4as
RWPVeWaN6Pb8Xejg6vHqgzoPezLGz1G0PRWzR09xlhcQEKI4sndYqWDi72EAIM6m
Cpoa/pLpTD0CNneNl/T3twl8fowiFTtgXB0s9t4Gi8yjuvzuFrynb1BGfse2427K
msdF1MM1TakQsydx+Uor+v3tNNoTNN5236vKabGYwIuH3nyHv3eBhiw6hI8l/sIY
PyDzIESycstJjTlikYarm5XlslcDl9AGogOELaA1eVpR8VlEmks0UZZ7BEGioiMC
+wFk7w/ha4Q+JQLy85MLlt+0XrHM24KfrUtR0DaFMKaRIIv12zXKwiY7ejRuASWL
/0bWV1brGsKQadnNM5os2urObydkIVD4Sbn1i7dw1X9jIe8W4LK0naskPqbB9z6k
dFyXtyqZZLCKw6y+u1hQohXWQForxa/DtOZakM5YbEcbPkHk5d053DmReaRhxRxI
JXb4hW/oldDVPAujPqpuGDJ8dAMs3fKwFZeMDi0ObkfJ991yocSDt6sWGOv+yyuR
yvM5XIJsV9ZERPGUU+UVyP2F4VU1FcLbZPd0lwfO81hKQxIjuHmo7JfTP2qliFuX
MWjwlqpCl9XjKR6omzhednJqhWcmtRhs29AcyWU1V6JIjieSQvWh7s4fIuO2E4G+
41BDJXmNIJ2NHbQ3gmW//sNekbfrAgbZHg3tYh3H1XnvxdupIMFjSbYkGbYeRT54
pHMSF4n91SHJfihauZnPjLVn2rpIFJsMn+KGg28lEumOYnke96epV0Mrz+2kFyuy
n3Q0ZdnOWORipW70FA/yqE33t77YrMnNK17c1uwDzxZrvNMrZwKLJNMuftq4n6+t
YQSPGUXuZ0rZdIvZou6YuYBJeECVdFmowxhXtusn7bhByfgc5QR0mJm5i17ek7fX
BxYlOyMZYvIsxLokvcZPCsShMU/Zzb9q+XL/A0cuddTso6agdlfBKr/tp3ghUixB
bOYRRoHi47plxsVRZ5HGaGixScP6VU3pwytZmMQfllY43KWl3jObHKEkppVeaiGk
Tcjo363xeY1NZ3ILj2JcV8n8XAF32acKiI04YwjAaF9SdQQiThzponm/A/eJog03
AmwN0DFJu58O9Yab43i9NhzAYyBFKS1qb9uJ8fBF2MJoX8RZYAnh9KUJcuAOgxjV
xEpnEU1imHmAiJbCyJoY3IGdagwtv6EgxxFej2kzOnfKnclFoViqPjVWGAHfXHDH
em8cI040NJwox372XHR38ovM4Lnv6U/Hy+hwFiVAu66APm9nQGnt/ZctlR0k9XBa
KwUW13EnYNEZks4QmWvC8uOjMj5bXAbPhs727EjP5WRJYj5XsulnnhvVI3HHzs6/
uAR5bTQO6+4quyJ1yNulr3qkmKZy5DmbDXfL4bmCq8PZSFoSTBmyWgU4SVCm1aAx
u8Lk+/X4OqYpDEzlpJyCeZ/gSwy78UmZUm/DEfWopHLRMhufRlNASLO1frjp/yB6
YYKvKn2c2FzjrT3dH6ZDO4kagEPV23quvrcKEVtJPoukblKmxuTEp+l+zYoNxaqd
16Y/Yrw2xN3/rGQYBQYW1uofzveuMb3EKTb0sGbXqumPKZQSZoEeG7tYcWQhMxPZ
uwOaIdTZ2mbOi5UUH5rzM+ljLsAf+FRbNjZSfLnPW7w=
`pragma protect end_protected
