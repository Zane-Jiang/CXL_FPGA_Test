// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
GSJUTpqqSHSt1qw+soeKokahrP+gSxzQEsOhO/9Ne5NvTaMrRZ2IHLXivh3jtN9uOTfAwRXQjRwZ
hoUOhzDHuCD9Fh7GFBI06yCQ1mN1wSLq3iw1riJPul6lBnCn03aBU3GaoF0pXt0b2IzI5J+ogB2v
QtdpNaYk+HCggogU0GZHdsOc4vDaQP8PBez0Zkaynb8qeBFvKNLarpqQCU9yEyc3U7l29GSk7SJY
d6HWoOyAWUi3NnGFthc9Kc/1ZeHuupd54xTW7IVaedA0+QL1Uhe9E9F7HoTr+MXiIo21wUz6b57l
dvrhy7RRXT6WJ7lFYpdWOpF+7ATDb25R0/rX/Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5472)
SxtT6m5uDxsqIYdw72zWhpsiLhY0LjDzGNpncTMjzj5yrSW4BYSPSyMq3vqBqbMU1HiwS9QLdOTo
49FixwSn4ObRTULhak+8CXFkiJDVmq0+PpZUkkfpMqEdGifQXSt7MKqcpR94SAMmk8jn5DvIuSL5
2AH9dK3n93s652vnuWgsLQOZywb8w0dfys5g828qqkih70rZjY9qyPLO7hDh1thgW8qK/67uCSoW
IIh3jYR+F66SsLhMY2kDeoT/wQT79IRxKwSUt2pJ6sYTsi61s8Bd1xUNjLzkk4BGr5LHWUHRYqsL
yGFNmEkUysXv2/e1TVnn2hWUJFGwlKBtHMOCjVMhKxXVZigyQiw58GMnwGivJTExSibMxdMRr5Mg
pzGLyyx0ZE9smoS8Jo75EWU3NX1+Gv+vWWh2BHOYZKc4D/XLmRhQstwdsERlzGGnUlZh/gPjaQMq
Ht5y2jxnwbK/WJf0RdkHueZKKof5tss9XlirCJWMgbxUgZBgMzu2lMu1N9bHXcmQ3HmYtPI9bbnM
sxqtEBlRRVV1h3IOqulcFHjVfg8UsrGdl5MerXr9t4sqB6ziI1yuJg4XL77Djs/3j6sl3nf/t+zq
GP5j3/NgoiQXaaKbZWOrnWCb/STMOqlOq7Ue5dG3ZXSmLSjx6OlaiH69JnZ6293K2YBeN71b+52y
tPXsp8jDEwTarWvrzb0mDyQ9+mfpC4dSGy4cHJGDKI4yFkPJX4VkCEcxLv4CjgTs/bXECNSNBcyq
H1J8tOb6R7ijoAn2vHWYBpCOC5DK65s/mJICbEIOEbIORX4KHTY1oQO3EwsJoWoAMEW4E4gelsDV
cKtm7j2NLjj2I72cFgVeZzQPuBXJdby49IwogeelpZQ81ANfmpxfnafH61axQVcdpHni9Ih6kTSR
bJvQ/BmJGSfIyh0lnf1loXoc8275uLjyVvsycnZwZAIEfGi4e5vuLicWIkGkKdJ31v5W/uGw23hw
/Jks9tGFOwoyxkI/VCZ3IgkHHAOOx7pZuxHi7Gd8L63/ILvyFCR9orHE210mGDMtenPn5NK2LqBo
/lM+ICOqX7ZiMJLr8dMvNY4UQ2l74hD1hdR8lm0N1MboyODkBL2efcrIqtZrnkczw5a3FaUzBYHF
4sSemgUZCUgWuBmmtbwImfl/I6bTC0DhmWPicxWO0U4ITg38A1UA3CgmM+vFqmE+H0nc0V7YRD2A
+8RUER+/KMzxlxTZiGmwRN9fipSwkjW4qZ2zc0yjmXPpPlPTPRwHxGvIbysd3pbbEDeOVuTmuqPA
fX6tT6Or1GiaatdkyM6TySSvQ77yHBxyLYLhf9PaN52i+QMN+VkhSZOEVpy6Qanmh/ROUOlGT2ql
SUAUL3q3zTFLmT9BywEoj0oRNgqrJS5le3VdT/Fe0xa7Bg6MEEFlIYycbQoGiiLx6BzJZuuaMVC1
FPAoqMljmeU0X5e0C8APmjhg+HM52zDcqaYCYZedoOTKPDB5eStlZFUIPmnXg3S4RX/ZE3TOzImI
TsehTjioSot7TCOkcTt2WiA3BQUounhiVJ8SXPYJCwdQV++E35/z7+aKf6f1oM2FKVdl/3ysr8Nk
bc6oib6p/4+ZC2zrRihg2fCWxoGWvzS2w+mNIGuzKZY7pT1QFhI2jgEVgKwiEFC7zJOW7uBDJI2x
s2VEH00br3Q891TZG8mJ7XvJNCyRIWHEdTDT7SABlNPFATIrhlFc6oa3WYNJ+xa+ldpnmHepS3k9
2PYFebbDjPnwU7IhE/dQgshX+lJcYRt6PxZe8Gray6I3BgZeEtXls03RnInmt+WR9oF+DLUvL2vz
6pjdaMGGmKxavxCYEeyPX4LbZhYAr3ycpGJFjd6AXZS9x9zYOJPHLOFnFurnD1F90v+p8rn7h+O/
FDW6kwjQi7SRrpgAaR0tzPRF9QBZDkpvGc+hQ34AILgcKLCTxbRfOZgGvR7F5WALL+RTTGoIRYyS
dqsNJOWMvCyYLqNoTavygTzY/PGRa6hjVKIoNfyoIgXEFwQ2PF3H/5JD56bmeLKP4XXjFPTiQY89
keMDSa1omwtduTzkeYXubWqorHaoHXyNIdT/73GuF3kve178hTj8Hx6dsilcIC83VgbJ4iLpzsMW
IyP+flK3FXnc3rUjhm+a6Qh7HKvN5yWJvvwvIdI/8+fTSajc6b/YH6IjiGO6ux4pfE4exwTc+KRz
mhbFDrA049VwpOBFlBX4Xosvk8IS+h/4cR4Yhi3YqFvmpOg9Lm5XjbGIYF3oKcE1sTRwTJdg0aKg
MLZlK+xc1axx55nFsY026KM4cRInF9nYLlSHoZBxW9TZZEWp/+++tEUFCu08VN98JIVFL9V+efD6
JzsuOKy6Kza0dDKq55ZqN5bnGFFMRrkEWGxXjW951C/kYA+yWfAmHIovjVrU3kOBUe1GqYMJDEtm
SiBd9pVJy8EC5ATLBfwza9m13yMC8TNceZFHQ4ctos/UZMF44tqHzK8V4Fu4OyG8KzLn9Vl5kG5z
vA1M/b9JwkKB7NmLHnujMM+ocAJVkrNDIVzrovZ29DdgxhjnZ7WZOfBkDC36S4bL5O4abIPF5ze5
/Xu6APTlgPVfTPzoOvd0ZUn2ajYCQB6qsqP4VnAbMr7uJcIrgo9RKjhJV0yceNDIT2i3UyRkfU9f
pFU7iY/4MJQPMx1aKKUm5mJAXKZPCPjC93J2LUrLkug0jkNmd+29YhkABqkHWZYWDJvpdbEnHv5O
N0K7nCHNfvYSDmeLyYqaRXL0hc+g1eNlb7gFEB6HwunD9SqP3OICkcWCrvXY4Lvtjw0Iq56oTcmC
0+DRQ3U3CeeDzLXT1J3x/Mh4D5JwygkDBchg7SNJgfIJVH6jQxxbmb0TBeANslEequuszz4S/DXu
KuJvcPbxeetKmuggKvUm2uQG6F9ji4lph2qyU8gJY7ZyGHFDATTj5dMxcmMFcqLFAOJjoNy5rh6W
1MlhgTbSnXw5Zd8VlNrA/aGIEE0oBXadn4Chmqv2KftrQwDw8ReDFWFayqgCjkLcx4PlVxzhVwqc
kQzfjHz+9heICBScNR25LIzBL2LeFb6i4fRTo2t+R4f2FDAmtnxlGtT3CgC2CK7bkFE1vsNu8/2Q
Sg4IklZHALf0eoXmsnuCnbsfVuvnqZMavdni41B5VKVKc/1iCq2+yDsYDVzZA9JDNvXcfAze+qRi
CNCoJ4SJUl2WeQIaSmsPmTPFxkx2HQ7+I6IX7HpG1zdZ4sgkkFEw2+sqaYQWpzJLbjSlfZgLAshY
s2iQNWzOTGtNPXYeYnJOANUjzEV9U+XOS/YwkqrDLU1qZmd3yv7vhDdi6BdOlbkYfZ8ynhDkbQCs
zYm3QOMHvcDrsRt9d3/oCsqzrQdRrP0D7716SuK4N/q5iyoxZyih2HOovMqrQSU6CW+xuqhnKlYa
vF/mkravGlsgOCcFZH5vV4uGtk/hdhQPe/T+7FUYzqxiOF2OcXIXd7IkPegPeplbxCdG1wNfvjoK
uiUMaVyrls9HWC+GqzMPFm5UexMZNrtdPiZ9ygBK3WTj7Hqxwaf1C8Vto1NOiuidz0ekjReIhoaj
3EM3/2I+ox+t2Uahom16Td4ivHkqAYtjv3N825Cn+y3F7XIPQtMTARCXb31ByXkQlk0dP+MB4BOw
rbDm0ObJllZNpeE+EaE7zBihegq5+zCB+/HsVXDUkeAbcdtte6vGjSSue7iarbi2AFZVKA3jXkXj
ud+tgpC2VYdgG4ENHIzvE6mmc1xA7e4zDJY0MkhI/UKLLo1mCsdkvRU0YbjQsS04KnC2muPHTZpm
XLxyK3sXbaJVSVKUS/NI211k3bQ+Lp1+NdcFJYiaVNVh5LO7TX34CmajrB6Ww37mu8sgq5tw8pGZ
kh/jr1Ah/pm4dlheZzbZXDnyy5TSl5R+uCCOkGfo+D0C9QTztrksxF9nwx2icJLieNWcWHvT9dtG
kCU4I95Eag11RuANUEjKu8y/t6Csk3OW/KyKJAc9SlyrsgT1Y0ct5ePHb1sjhSxfZxVzHvKNfGPC
UlwQvOAlndiALU9Oo3KDNvUPt6qppBCW6yzP2km811CVuuCx/3pJw95pk+yFC8kFwRWm6Raq6bMF
6df9SZtdsLRxyrigQmbajNEWXOx5HjE4njYg/3utmugrLjp8DfxYR8eu8cuMkmT7ymCOJ0VHvYpa
qvM2uT3W7x/0+uygpUv+ehUFkwlmoPKANBYZUdK8Wke8Q5b8ff+Q1rNlAbWCLqEEXNxh6eG2XigY
St25wEZsdKPp+efP/1YXSXZt/Jx3msDZOilHcLndWRE8Fhm/WQNcrD2ZuDf74XAL6MM8B6GiG2sn
JmpdS+KqhuheVdq4770sXOxc3pWNGbCkGChhBiGvpM1CSjrvpcFifNhtV0UQNaxa0g8ogL8Fc8pH
rMhx5rXVpTajW8SxALa8oTAi/y/MT+YWc7ufJc7fuolZBUoBsdo+zkLThVA7DGwEBijLiUShjPkU
AjBZsM7RMSM53nmfL6hMsoWz4tpTvbnxhyyc87g0r4HzFuqM8QWICCScY/87TYh4ChwlT1SiqQ4M
qqoejQ57HCPRN7d4V9aPlDSBlgP/h4o5HNNrWNJGPLdrQtDrKUphxfxST70pT4L/TM3hIsCocixo
G7tskd7TKmqKJOxtwi48kldeqa4zLA17WfTqdb+1ox7HULUk0TSXcbMvHZFkiSxrzK0lXNZApJOh
2gp4EchoVJBQbcM3EdYZ+gYNxVvfioXlB4hqLcBwaAvPV2q88BpKDvEtVma48FwJG1DyLyrwgQYl
6S2wqOKcx9R+zNaOXWeZiocd0RE/3ZLTN8ZST5YO7uqgqF43L23zfp3nXq7Yz138pRWFwCuBEnGf
K0U/FOnFKoWL/HxtzJdMLq7jHmqCmV6Sl3l0VuQZRbHMOpNJITLn4gj+MBqAVPaNWOKjGJJhblC3
NmKf+Lo15/4sfK1Vp3Kgj8N4EdSGLndzJg8zwcP/R6fUSA1iZ/hywp42HxyFvc45WWMJIKXB1Ys8
X2cp5mx4AGhuHI8GSvscu3eqM+1mdyB6xIVtoEbTL+o/HXQnggJyYxwb2hkJ1WYMMRmQiAODOAzS
0t98xObmWxC70jX3V0DejbKrcnfYYgh5a/gTrqm7xzEkNQzg6f5VLYqPgaRzOO4OCF2vxvdvMomT
pnEKAdyJvIYnLPIFaCuljjdH55W7EbkYvBrrr+mnOQCQbWT2GljJbAQ4/Ay1j5vJr/wc5/4n50AI
cj8LkVul01jXKEKHOdnSVOMt1KNxlIb7pJj4eF8wo63fHffQjs3+RrtPhOEt1yTNlfEvmz3DWD0u
70/Ska/pankfIF1IKCti02dqQU3mbRqDOPFki8ZfVUiQXcuWtDBSrTbnz4vymms08upWY+YQTGZ4
VmqiBqqI/r+uGMzA9Vx79BIeUcEfjKZUv7OvJudsI2g+R+j5PzzVhkQE5BENTfz0CAsIWqM6xCYT
UHztr48lrfh2frEiaF5rZxrzzznNZUyQAOEOydSDEH96UpNzOxQR1Cz3pHBwPem4Y545bXxV6Et4
GnX8foksGseUcrmcay45MBnsuyr5toQtSLZuhlf9znAvnUaDQtifbsLbIG2QdG/ZXeR4Eka0d57i
81Hw98a/Wf7c0TzSRg/FqdgUWHGnRYDmmhUnQTwLNCSIA+745YZRkF+kwHbS3gX/f3mCFo6ycJYO
HBg07kBl2sXPjkr5ngEO1VLJeroU87ac2oAh6B/nHK5aJvLLyXGy+KKZDPOHEi+5DlInbK51tHQY
1pvI9M0Ey0gTqU9MZpGdbRnzyXRpwKob65+JeWj8ttAN83xzT2z2+52/sKHPpHxBfk1zt3Yd44hw
WnXhZIpaOjl1yD23TcnEOBU9JFMxqOLw8BdwgRaCEEMfRd0h6JOMuE2emY70Ky/OdQl6or4eEzCi
d6cS3+UAcWtEF1iYPWGGAv3uMhRSiP344gWbj2D5RASOG2GWE/dfJMQp3AJz6q6prQZ1uKE6Svct
eOb0nJ+FAbSEesphb3JeG7S19wm4kEfW7NPVBqHx1iSt4FAdxvksrIXeW3BAV14GNEhlK3XAqhJO
kBPKrPDs4B92A/k0ZjXO3O84ykZIw9G9JXc+0r68Fp3NWUqH4bPhM4n3+uv+tKRJZUAUF1UleWtA
h6fFr+mcL5yxK1lT4aorVz2P5I0jR2BeBBtVEESO53ucTFRyzmkifqpY9Q+pfgQ+jFgpwLtIOpib
r17kGE7FBpis/1ay+JFnkZQ8oDTS/tfgLSfE7zl2o0sj7VpQeWkF2NtDsFEa8RmyZqcstILrpvmG
P2vHaFMJa2CWhnb9iC/Bn5K04U1aZ16Vr9sVxpP0L6gDuGeNtTFBHUK1Ng2xWEXNWCji3ADzn/1H
El08nUC2DbVE5fVFq22L7hA6+aygdBVb0qwqed1al4do1kr6UK0zLV2wIn1fqWo8ECl1qrzyX9k4
dbrt+AB6Y6NoTkOsKS++McHVa2eGCiDJKgQrQIRY17aSzOmGF4FYZ3GhZ7pyK1mboNO6X0WuVnj3
e6mvFExBvQhHQHtaYZhanUpUKaTZQq47czB4QLO7KyBbSXcYXAzaSwsHTwJjkdKWi9uiSJzqa1kc
ZfetwsNN14NW2NgbX7pohnP/JgaXM9r9ixbbKtizmtpiQd/eG9Z/iHNXuvpQZK+FB7e4/8fMhbSq
euNmGJFKEHMPsNGEnAtE0KGwcvrYtjgdDK8gETOn13kyYluV6a8YU04nUHS63ya4568Z7BwkyQ77
+vI5b+IMGkleNBTvQQWod6ukihKkxkRBqhgue4E8ewj6Sufr+M7B1NwTZ0MNP7SrV2fQcSWT6mmi
zuZxLJs81eYQwGjz+H55vGinDwc/it6N/Vv1+dDlmJdmswQNkCZTqMsqiDZ1UOgUoZHoCgBINnPx
rAMce/2W8IqFUa+Rkgi9JTOMNjNsfaZmvYuPcoAu5O7LGJ6uNnAboAMypoqovCAxn7kNQQxU/a+E
p9rmeUK7mGDtFe1teJhx8yeCwy1eyQewcYmHkMb6VPKRobEzJ2jhTF3ajc3Jg7eoRySYLqPm2z/t
zf/HuNufhKHupUnZ/LWpgOMpySa1R8lVDJl6lhka2t/84RaYPpCC1FUdFAtdOb7HxjKCBANqOXzV
HOPUAe9bTpgBDkC9/4bwvhB+nIaHkJJqFMoVCUa3BW6yeLFhRXpJYWebSwpHdEU52Fgh9ase9U+H
25Q71YJgJOswyi3Nwp4Oz1chJgwdAdTs8tKsT88OZhDpDHraA7113tUkx46xzVZ601tsuCk73zVo
`pragma protect end_protected
