// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SiqfVVRHf4S1u3vRZin/niPjh9HUbr6eWnjDoPxL/+q1CXr0BlLaV3qikGD0
arc/+H9uZqTHWxClALt+fu9pZkG6XF+gqJXIHiTUBRVp/LYr5dsACWgccseW
5FypU0htrsulewKnBqST4CZehaPGCz1/gyD4qfMz7gAsS1qKRJbEfEbCaPCd
dGcpIAc+coUmlz4EGI5n+RHq7LiyBVFSvEX6xucY9v4EwHGcSzq7CQrG5m/M
gG6XGFn5iqUzxUWaVd5tuG5ZYseKeFULjLHEzmHH5DQELmEWH8enZq6QNlVk
FdgjkL18FrOEB9iX83rWmw7aSav7kEMr5b1KpEzZJQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hm4wGrH/P67bLGQ3kNrEqQiTuYqDh2zbfUydmWpBNC2EUO/yMrIXPgAhrbwh
q0zhJHn6Ps+fN8pTV1G0tR+PlSIJed6XJmbqX3kmqYo0te47sZ9q9fjtW5Hv
qXlZ7LIpMjQYbSm3kQyquVSVz2NyqikwMlxfJhcbgURSTvVfzSkIMbhqPxfQ
ioAG86vsHuoN2DDob5X684IKh0XCYjueW4/l8VBWEc5dXTxo1BQD1eJxIAnP
9TVZpx+KMhlxdHKb992Mv/SF9mzrpvcCWW9nu2khRmhSSAO2IGSQUUTI0dXS
1k1YVGK9n7SbkPbqDO6VJn/cd9+xSTDG7X4W/d5Dqw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rWESCtM8g27YXMKHhJPQzf0IAjCftKMVrF8aSRkhvBOvL7iwVwVZUMBs8ZDa
Q5QEFwKRaUIbJyK/eY5AEoGW9LPB2P5ksNSLK90cVAnshPoHFqhsw3JVyixl
BKQFITnm36jmB2H/SuG6yo/jjAsH7kU273DlQLbV5cJeeHJykJb8vIJ5DZfA
MwkssYMCqRp0nbG91zRo5G+AUGpv/RIiQQVZDHgobQXCJikcLvkconEj/eZd
FBQHMX0SbgKjs/McXaLGKPlm1siNTEfw8qOzbS+sfGoalsYmmHKBia43VbPS
A6iO/6cSy3t+X8cSWLeZagxJvwYsKX/yvTD9gj+O8g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jsC7ppxOcZ9lQIFAWrhQtmyjPgpfIC+SkSss5rZtT+Cq9DH/gDgH3RtToMuI
yPbaKtRy0WD02zcRpbYOrzioctvPhJOCGlQ2Td2HCVgyCizUiayG6DiPZi67
dHDaT5WOnC9G3JUhXkQUs8yBVKy0uNAq2/Bmu9uJ6BySy3xNj4c=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
X1GLMGrR84tUP+dcwZ0/VJ4OXf9M6lBL7RKihtt8yVI2muXA3lu/O14/lBb6
++IFdnAsCvtBFDQx+ZVR72M0Y03u8iJr4HhMZsa+9O93ifNoYhSRDHKgwJ7G
H//2y1pDcnUwpYIIowascjjwU0Rj4OPrKg7D/o5UDgYN4TgJOFlwFSwkKSlU
a1VYzzR5SYU9Ssb7fqIquRanfoNpZrGaAlvmvVoWlIBNZrbe0Q89p9i4x8xI
eqyrQD8IkH6Dc1o6t5w+tx3sDsrRveSNoPqA+II5KUgTXDq0VLKORXNNWSrN
D4ZC8dBZk3MSVSJBaZGkiL5HJHLWVZipKqoZaNZdxWuYY/riLsI83117o7v+
nJkHBNqppLGhBbe0W+tammHzk9dAkgz7h/yFdv8OUCScoqHKCvL1Kthr5cS2
qyR7EVsHWWVSI/SbBFws7umiQJfdyqSytaZKsGrIYj0NxVCH2ALmOI6QrvtS
PEwXxY6UMMSCE62ZO5G5jH6l79xfFP6b


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
V6JBTL9bexCcbg6eIdLEbDHwP5OZDzgkESLQUnSm1Jr+E6e+BQL/5gM0z996
DTx158iWC0pnr3Pm/Uq87YJ5z6FtMfXqWYDn3OuX5R7JmTjxUqtu4JAxdMpR
Cn3UYwG8m+75sZShocqxbhs1e6+mSTEBOwl1NKmvnNzT/VD7Jc0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H8MxuZWfONFTI7rXShAVn9/a30glG6F6ZKGlfY2PsXXP2z14dNOUORiDyNys
poKdQOxldJkh70zo92zpXiETIzs3Qp333RLeOMK8mS+bmhLGn1xyxAW44Glb
kuFXJnMHVY/Eu34s0Uqq48UPMnXDh6ylHyeR5TYd/2CFaEdpGsc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 27680)
`pragma protect data_block
1OHJ7Lb/NCZI71gZ7bfDXvVOmqQdqJLj/X1slKwtWrVbinIlx+FAKzx/uQ62
mYJo9EyEGfGJtOXDmGqgZ0lGepEyChbQV4V7OQxawFAz8p2XWt2MONvZ0snJ
CVksjGqm6UFR2F43abljh99zLyxxv9lrAd+S3yFl88dsqQbxW5q7sIgREZrE
phDzG3cItLsUHCsrOraR5Njo5UIBod3/bpotoPjMgaj7SiKPpYnrBLTdQnAV
S91imim6KtS2GEz4nRYrxlQQ+DSq9NpGC5M0dnwVctUQqnzdezbD6LPMLFVS
QboHcXcvqxHu1mMiDhm9I9XU9zS3lidumes+dvcuQ/q/w1RNCjyFxpDhpAqH
2ER3TfLn13+ZPojsvJAfgvVz/To9Ja0VDo3sr1n6yIx3FT3+R56iItcTV+7V
7LovPIb0viIH1oIw3oyMJ/uuhmhAplTLW648vREzB2011HByYLvBgwZ1YJE8
Zcr4LZnY4dxZK4/ttxS/GyEzuzEHDTLRMlZO4GURMOpUkwrhgmuZvMdgkfWb
5dMuwYtXFyMVYRa9lfuKGmoFVtTCZmYRmOQdAsyIoKZdCiy43u3pI2jlqWJ0
RBvnKHU1KZnobjb6lW+fglNoUAr/EkztTNQFc/PLGDthie03lZnzeJI9fnvf
snQf4PnVvKSYiIKoivgi2QZeXdK8OhgeREZ2UEEghYkwUkWoxirlD7Dd1ii7
xcvw3UBZieXmVwhmvkqKlrw9fw4TUayVLdJPJLw0zC6q846/Da9HR8k+BS0+
1XMv/ZGdm4ozrEMAjLy98H1jMNIBF9YXngF7EO/6PbmB51teEKPk2vVgr6iE
AwxQR1HadjfimCpmr91RxC8ItvLvch0LfxNg8vp1AMUgFek9SZ4O8jLglmRL
cdMkN05mneCu2fGNu/mUircFL/kcoxDGQcASRQbDB4y1cBhxTDSbYCkkxhxk
0XvKAVXeUEiScRy6wKoTOe6hU0TWp0Hbrq7J9OyUbYOfoe8oMQ0Y+L2chsxp
3dJGeB08S3YtLX0zO8EV+DkSgq7fS8QRYS2GMklfHOvDr9BmIrfjO8ciVAgy
YyGTtdxftxZLPnviqL/JkMRdVvSEQBCzGFFW2cC76VA1yGARZvdRnWyijcbt
TfnsxdQ5A2riGeHJ9bNtmRa3Y965AUqa4XnaY6d3q9o7J2iOlv/+/BV0auxj
kUVM97TT86RHfUH9MhQHO87VT6eLHch1yQXYiw3KFq387am4K1wZ7RUknXwO
/ApHz+ZgXsGkERiijYDo+K5cIlWHE5FZ0aZ05pHg4u5Z9cFd0y6ihnsMlfTE
lgnyGDL6p9i+s6rKSl4glDpEDXHP0SKUEQwKBKEyi3ramBCn7FmIRL7BN7hN
0LEa0Gu7Kc0h6F3nV58De/oeW/n/aZQtfdwGobhHOjoh/NyFXDyOY3jog3k6
YbKZqm4ONpFDk3cO24ysyRaYxGG/EBN5Yhy3K5hr5xzlx/Uu9TNK0/OuLP14
VkbevFby8oj+3X4xwh4Pz6yndau5ggdHsU+dro/BYmDZvCDRXZjEwzPyol09
PNl9KeZBaYtewYo8c04m6OxWIsoZoahsiQwWNNamR0+gcGAtQ4gCd/XoB5RX
Dtkya0llTZFe9T2PnMVQRBEFQVj+aCrNZpdx8XhHD0BXoe+7UILZKYo95VGf
WTRACBW1eDRFS0rK5obBPiejwN09pDCZThL/7k5nseceqI82mOlJsfl4C9ny
STxQDsyMpM9WgB4vdVlwNIZ/Q7jsUeByl6UOjWcFOM7ydHUNLOR12LdCGAaI
o/KuCClAz6TGtf9mBteDCiO6KuexO5peFmJQzNvizHPY5v6OMoSiDRP15/3c
GQ64uvODATOTakWi0YctTXdoJTM7WywSgh73fyRG9hILlUBxASZ+0M3qqRtf
e94YhhEYzsGD4H505lE5UPt8xYDYY35NQiEVb1Cryogc/AcdNj/kiXrdURCf
jxt/ARAFbVSt4bf4d+c5/vNvIj7naYsuGfLN8ADpuyxOO/ZEmxBkJbERBDDo
fCovUGr2x8akNRDhNAGIzN7ykMOndvZXbuxDFlUOa9D4asQr6menz7HgLPjn
MvSSZyR6nNDS/MnGsI5wfmGQKNfshh6WhJLcBJGd4w30ao+ibHT3l8eW/Qgd
9FVzlVevcrUfhY6wpMzrdQXPtFsE5Jt3MU4jRRjoZRHgX2jGfWNizbcPGiYn
bBNPhGIVj+J59jo+dG2T41RvWvbAXKEEANFUo7qkxZPgVH5CFXQzSxWzML+a
dr6QH6N25AjRZZjErEyUVzQG36S/B1IE+MH8wJWgUUNL4irPQ/ia2cEi1C1U
OJ5B/HWDnqKTkpK6xMaiTPYlcYdYwRkiEWz4XwrpoKDTQv6smcH2fChtEKJK
DEz060dXuEafNIU0C6ECW/tnu9dfbu9o1JT75TAR14rruUthBzVa6dj2ZgCm
SXjlrGuklUX/M/6tkfuIcFnUqGq86k37dKhaF6RykaPcHWA2GMTHAjEwpwLQ
PrLvYXPF3Ih8agXGE9pMwL/g5n54txRAHhGKjFMiTqztu/JkTeNmX6y0o3i5
yu7EZuuDxAzJ40GdRIY2/h8bNaG9yCwP8ZyCblVQOMlbo3ovJKBQoEbWoAx0
o0XnYOTNkfbMXVFgbKfw+cx24Vvk9+BwTTCtjojTAmCbNAcFyAwgq1VJITxY
a2w6aMbJcJ4t0jZbdBFFAgzcFYXovhEDFRHRCwx35DEaChq4PoY09sk4ylHg
oGlETDPkVNf70xjKODWN9Q94WEwPfWOfGr/lVagCvnqp7DbQSQaM6mqAVC2R
vQkCKC2X1i5Ad35AwxmxacDv+y7fI80FtOgKPIkKVhrZbZPoq3+6958hTv4S
qvcguvm9oNjogA/+TmwlRxUzcyC3+51yOnRB95vHWO/DICvH0UhQEw/w0vfF
kGdhYLIRBE5c5mnYvJEpBjkKkC8deD387hTJVqW/aOGsvOu1luhwpT+pGBmy
GfyMhj2N+lVCLEyoSNy5aG0yl4YcP/CkmRuLQtzSWiV4ulsX/JsQwUnVRErJ
XIW+zTH5oHTmKtdwI+RsQJcKTQ7hcjCLRXuj+8A/pJ7MzAJbcdUJ3FJAvGvH
uCFJKWjLRv+s9C+VJDjAzklw1jpBHA86lEwTyKAEn6q14KMSIOmYYWS2HMSs
bvkJSonfCGStEk+TnAtYjHJX+ZAhuJvnOuesaOeOPBsrg8NF7EETpGVV8jVV
3/+huh0Q7gHjmb8I4WOY6LTlnfKv9DuAhwma8Rr8fIjB+GaMaz58vVjCE4H4
h8mgtf/0dtckvYjS/Ra4W5D1ZXrH8k+g4wpKCNtB3Dkak0jZ1uFpllfdd4o5
3CLJFAVRo1jyoSubsSWLb0B4wuilpNDx9JFluvwESZHsblN4RIFhZAwyeIMj
XDPNY5mq8Vd3a/Npch5i5GxT4M5dF0RgRE8Ys9zqJNtw3G6uaA/gc+Efosf/
lZhc1xKNQ7wRG3c5BASViDysnzBt3DiDy7HX6n9nFeHTbE8kvkGvQxEcW/5Y
+Nr9HjZhb5mavm0XVkJHZtV9JxKzaKLu2SOYWMt8qGjQofFOdSRpT1MDphfN
gvngelhjDDtv7yv3xWo6J+dLPoQnUUUX3yKwZ3fmvjja7sWkOTVNxeAfGDvk
ITunXoMBzsbk7mTuN78wX6zk0XT2nc3gBt3q/szaH1HhfesD4vRAWkNvyQlX
cuEwgza42O4LT4z35CnzT5WJ4fc/D0si7Pznb+i0HcGLtkbw6ErcyHqHSg1j
NSsb9s6E2jnULGHnS7Rid9Oaq8YTNUZVs2JmqbE++3GPelfyYLsSQlI4ibvP
iCObTzpZNq/MZJeFPpTQIYQ0r9B3yWv/7I89Kdn3e6MBg1Egcu6g5SIt5g5e
PZN4CimB9Iz134LRZ4ojKRnVTGU7cTWJnSot1KDgFPzIUKw6ZQG6W+EsYXz8
fE421c/BslGJdEw4QMv5llbWVZ4kaISrwo7/zE2hDqanygvKVw0So2zw2r+Q
YCK5pdLP2Y6JtN1W5X9ypWM9k0LjYxyaOg4sDNNuHKJH7OxuuJlrWRZlFfm9
Q5W7Thz2Cwr9BpMso2UWYecPWRWYyiisnCL0ehGMV895UkgCNnWMUWyZK+iR
d6QWucPt2j+fNYjcNjSRMI52y4ZdX/aq6Zqljc3o3MnrA/R7zTTPCxDr5XzN
t+NDYo1DSjVfMsLQiw7wVDJp8KrhaSVJD/DKlNf7bwUrUGsdU6um7Wl+AvGU
qsw/9xQ2ZqNkggMRDh7YOazwoKpzPOaBq2aaXlPQZoDbXdqO6OFdzUfCuP0p
IyAQQIzKheiEXWdArR82gbStT4ULwVibDGht6eqMTasa35fkUA5p3ctaBH/q
k7iR2OE7nEjrhJVI3XtmA6gJC839eUA2zhHKkDjFqPT9qXcjJCJkaDgHob4X
jDWVELVn6GRamT5lg/3hA2/2KzwBd3CEseoMclRsnKRoo0l97mKloiJNWwVD
eKudQ7Ex3BiHyYMjBQ5STZiFHWJTMt1NQYQNFcOy3MsfZIJUhWBGzu05791K
wSLQx97YJlAaDZq4wakI2Wxc8MGrbb4n35f0SgYd92PMFU75Dw/IpxCoIKJQ
b1AmHWfE0joXMXQFhmO5d26RiG5TbRXepZJuUFwnQMYBh6p3GwQnT/GTZLoS
FCmw7T+miY95RcB0M6ldK8/vog1RcgOlnMGEFR3vFzc63XL4M2zHMl1w6okf
+9NFZw5EULAsc/Iy4rtICuVTMbPGzpdhm+HTZCrq1mXDBXvqVDgzWxSR8H57
ZRX80B/BKuWNLMYh/W0XSCKrnpfGlUHSm/t/GuJU5AKU92VH4mW7vRZnYlLi
XSOIhG8BJfUlT8cVDPycVZgcb+wNQbBTW0k85evW+KUTLiUQR/GPEkXm8UC1
xzsQdajcDWm/b2H1uURWQKVrMK87IstwsSxNUTHtnYVhUJZ8IJGzsseyQISa
cKmRpifSE61xvQwVMBlEODAz76H18KUiJseBqK1itYCUZmmEdr+f7mx6V9xU
CxskBpLJFcBvhEJBi3+nuqdD43CQ7gMqFgrKpVd7FgcNY845nE6VviFlM5pu
xJ3InmDsAyu0vtFCQTQlloFL0Yuuhn6yuNZTNT4q0HII0rUN8+dfrjhed7SY
45zRmyoTX6g3u2QqjbqftImSj7Htqv+CXrFg7vFC5F0psIzdqPrNavP7YeWN
7xdH4nDvphXzGdbtZm86fJNy3mJUZM9UGuToqZ3nCBm35/IRW81hNYP1MRqL
1wFTRNaw7oDT8yoO1LUFZo0PDKjyPJJWOQVjqBYkGlOVYgmcydhJ83vTQ2EN
F4DN0HhKVOTsURBh0nw8HkWzINa7QkXSPvtDT6LTM00QWGHXM0IWMwgMec/I
ASw5VdHX8pO4HEX8q9kQiZfeWtW8XHwTgwOUo/fTjkdjLXzOcRZYGgjbAeEq
05KIIFl4IZ/o0lti92ZFt2LgH/2Fr+38rhpUB5K5kMRehKTfU1g+hVjD0R+3
hT3kpjJkVolnaMysibeiVUjT/BZTisz3i28lqm+RLOQGZ4fFKhSn7bUWr6p+
Vn366DznwsH0vVgY1VDIVOeVSj7b5OnWwoS1qf1VkD71FdYubnZXvhpGjxXh
1m1GwfBTyROjO8//IraiBeNFqmhygK5Jiiv6CrobCWHYAIPt/bSofZw2NqCl
0bOp1QOkR/SOSB5wzg3ElTYREqDHtNgvML8oWL4aiO80ybj7G0tbX029qYkv
HSOqjfvF4y4S1qLxDD0w78tM2QnlBLnAqSPilSRhqJTIlNL+MLReEBJLT+V8
gNUwhjY2CLqc7LaMov4Su7d6c2WFOrxpXZn9xTsPLCn1tOiaoSzJKExbl69S
Cqy3ZgtlA/cDqR6e5rLpOb+4cxY7T9vIqAqDMzYArgNnQWqxS8wf7GuoHnWA
44YZuDoOPFsldqtUpcGkwkuIaWUnDk1YH/hK1fd5F5PIk9YejZmnIW424u/D
t3svt7Iw+1vX/lC7o9BA111wr8X/kg7tcbYn/BtGEed8qZO0yWDnNq/pxU8o
xkS7L8p2QJjIaAIYhIaKzFj+ImUjkvlf8d+ZSDoGmoLuhCjysbXplII3SFC9
D0cyd7z6tEXOaF1j0vygBa6EN15iksx9vqPB/+m4FRpmz9Vb89LbiO3gqWdn
6UbIkD7MUmALBT6s1NoRzCW0kNI+QNY5Ner/Rw+Zeecs/5yymft5+6zBHntT
sK4gAXVP23KGLlli5QGboIq0/EQQ9moZ3suQQ51J4lJ1h+jNBjnpJqmSypbH
wAkQtYBOg3khKF4eF8XmQzmv9Q8K204AlQK0h62fnA9W3ESfDSIejeghYF9L
ubSTBmMeJj2VSInzhLgt297YVAcBgCAQ7iJ8zOn1aC7GVbJGMQXRfuX/e/yU
uXuCRNgousLPEQpgrihn7hriPU28t0WihUrVPyxOsRKuBK3N+R3hoqst34O9
yC4xDGs/Eup6oEswRRBX+butPQx2XI8GTlRm3hYd4I3kinsbl9FJx5lBxEoa
mhNQc/Mi/rxsiRQHSIhJfqIKcPd4K2zdfJZoCRPraI+KQuF9icrYk6X4/0Lu
W9BnSqyWa2pbinY5q5a11if8gDy/1Omxna+3HlmdQtL7ASbN0cjX8LGjb0ZZ
7EmdtkCzfVGUUXcuR++3K4sjmdN97/fjR7CywvHThgG8HzTKsx51Ntk5pNBh
tOLkHH9BPcSqHC0xRhde2UXze0zmTMhDz9aJBXKgLRhJFr1iCPE524OwX32d
0v6eAJPMjkTQTWyHzdwRfUfK714vbN48YfjZNn8HouFGn5kJQP9H1h62wdbe
qxM8ObrES4yMqINMSmjkv19ehbhexDedncJoKbmYQrlTL3IMAN6tycwatxiR
5z/mbQz46IQvoyf1yvYxNVGH0kq7aLKoN2/JNjlTQIjHVAB7B+ghkta8NjB/
cNDiyMOopcjb86lCV3fO/NSHDfrUkeYyvkgM1G3nHJPwwQShu+CoZHah+MNB
Xr5PGv0nLdByoik5VrDYjE2G4B1N914QIyMWDkfn/2h34rk6Kt6LBYwEKsPo
zZgpY+5r7IpGttLtgJBgxUdWN7AsaMaZlPFSdNXMem4w/HFvVSXTCIIhZfd4
7kcRjfBwJVRpbyTr+5KUD/UTWpMJbVQ9G34B6su2tKZ/lW3xTYucYb6ELqwO
CL7X0liDQ0Cj4AJE9RpVVKgC3BBJZH9jIqb5Qpr9s2qN3gKd/Hy/dHJ795r0
cMP27De7eTUTX3lka4Fy01H5KhwjjDRmLUui9iRGuBhvNQcxmrcb23+k2kRc
vg8Z8yQxUY2B2z1DA1gmApjxbkn9RXgInT6yUc02QSldlw41szPD4rj8eBie
mTT/63Fp5okODyLunrb3wyMiHbjhahd3zyUNX2NacGeTIuA/TTXr7l0DdIsc
BXQ/fwpc0yHjEnEZKH/fkvXUXvI2VwaBQ0TZTogdXWWP4l7f87wWYKdt1cEo
vt7RGU2m/866xuUY6ggc2N9A7Vmaop96pCAxO5GkQvA7lAM3El7G3k0JmIUW
+oWuXeQqaB9myZEhK8akIvqiWRwEYAf9TPVcbqz4uh97o0oGPs4ogCyGg9IT
cFcjmbjOD+h8jvwhXUrrGXsz+LXFOkGP4W9b8xDMW1zVPPpQ9zWiGgKl5RlL
3n0CdCdtqbgAskso6JtqX/8jIkjA64+mNDU1+p1SqB7+oM20CYaZeeQRSb1L
jNNLra0UzqcHEjLvaDl4UHUvSQsDWKDFtdqwKllKQIar2h+AQxYSQk1Yj6H+
FmpQsfsGzYW9gjqDHXs2JCBTmRmBiaj8As3dikH8EErTekcr6Zrof2atbqDe
ZA6m/LmEe0tQ2L+GOGd6H+eMJENdHeh0GZbU8amAs4dvX3uWgS1a/UyR95QR
TfmJvu9HbtFyT0YTeJvzBi/dfhAasba3cqUI+CbMtb5XNnpPj7noKRRMMadj
ZZkbRZvlv78gzSVzBjAOs6uQhn65BAgcp+jaIO02z63If2oMiXkmjpDqcBDK
MwBrI/uPRpsx0nr48qSxL9Q9to6Y4PbDDpPVlt7k3BzUfBTMLq8SA163WkDU
wGpm7JoxojAbh4/MU10cTO+ALinkCLQRD/a4GRVFIJJP2bhi5faRj7PVdG/z
MSFYa5eVqO9PTzCEJS8AnN6kb7IRNeB05C1uwUk2zkhz1LsmmJg4TnPPibZN
IkxB6i1Sv+u7K3xptUr3J6Rs4l6lX8GAo+KFP2yqODxIef0fRGVGMLyn6fgd
Zqbfx3DZU4MI7ri3xdQ8MiOwtprNjxIjaE79sqKMNm+RavKPEFFCplT6BJj+
ysZhJc/Zy92v3W+oiwV6iwd1mX5d5IlqGHNwitNtLvuTk6MljD/SONV7eu14
pvNAKAzcC6w6BlRd+XBviiPT/A26kKtJAZDj2nAZrRien3o3tZh3/HzXMbDI
IfrnzYZJgNbQqjJlS7nSN5fwj9VU5QH9w7veTHLqv+sTifRLtIXlmgKTFC0/
ehcYNS4+5BmHhpfMJs6yfSu2m2gjmpCzHq5yskMbgXRdcU3RS9tk11Klw07A
NOlk3n/UJ8syWq8mi5qFCz0Hgn5hK5z1cdQDgsHZRuJ427y97pl3Z+wZrER0
PcapzX9SaFjuOZzRiP2PIwg5HlUUjh0HBvfgyh2WnqptzaaZwzEuEcSgm3Zd
XDPOIgybLuiBjhS+H6UhWHTc2WXOFhdUYT3yVu7BBQneYOHOvUaRgCSm5OTC
8dJANuUVped7/5uM0ADnM4723vW95DvEpLwpLyiHNa2bCnXYrRg9x7JkxquY
ampNczITHUWktR/BApA9Txeh5svgo9ifgLXs8s1CLqoonmniXAC4n5ip5twn
pN8q+0DlhEWxnm1573gFAyMkUfjzqgw5ev+xYV3IQ6gVlJ6Tytrt+WpQ4GO4
Na4KXZLPqTyouWCGCEC1hsbz3/AFb/sBk3ALbEsbWpF0kbxqlp664BUiJvwF
IcjqwpYp+no4DT3/xhPp+MkDlxgjShqHIvQiIThR5en1tOzsR2R5YzIEGAYF
lI9/2Cqb9xCINXnwpQL4mqo9g9NjFxN5ql7sSSHSr1qaB2NLoJv/YTwoIiRl
0NgV8BwASQ35Msr70f2ILgOBp7l1j6OY39tr7pQ99EE3GWsJbig0HEW+7/5l
t3X/hnrjPQ3iSZL4fINSJzw/HWiQG3O83e79nCY8c4TiBmOnGHsevWi5PDpC
lg2HnROJyumXXWgneDvXwoF1i2tvl2Vx/lPdevOHF631yKLV9YoANaWtt6Wl
gMh9nKPmllgu0kLU/zGhslb/Mwps+ZkksvdRV1ZGLTnObzrJjGH4LaHaXxCs
Bcx0jEclI4ooBu9xlff7O9NtrDrwZKj+e24t6LJghUgIohBSq+rjYGISzH26
QdU1ccP96hdexUq4sKVuNH0NuJcmApM1LoU/yO+AHQSw2KoAtVxBLvHZ+/Jw
RQuA5s/gpXkkjEQAZyk7ErpvdBh81d9PaTUrF6NmokNvSea70eu1gdzWF0rI
nFWOYmM6mnR0TshjxVm033tmzVUrAzBZUGCzp0W9amg5yC0mNFu/EUmTapZ0
VQP/3/8c38G5gVXRGuYD78sibQ1eGpaBfw+LEMFldHcxTloNI2KcEL5Vc89V
SlEQ//3QreLYKJD/q5z3Rg6tOKy8iAEctvOhYM35SsAf5cUd1PfRxP06Jz/X
vHCpWOUl1DDhxdlMAEsVKThfrIBnTmT/qW5YwVGcSzNWP216ZjJqXnAVlw0Q
St26rGoG2vBtxd1KdEu05phowEx90A42IsYMefzpM4EO52L6Vl2K8x4Gg4vS
XowOWT0c4acil7ULG6inDTD8wSWBiy9Gj7HmWoolLKa25XImiOUJHv+fCvd7
KIOi8QTnZ64tfgKCZpiJwqNmvn+uAROsHFDBj6vG03IBsDywcAuAhdzs+lA8
S8PV8sbGRpKAT4ItRfIbUVTOZWoOkxO3AxQl2vpWSPzxDLDacBAWGpQeR3hb
mdb/ANXXVBlE6wBBWjKUlFJZSnclZDskrE5oemOIOQwQRMCkvd1qmN4JmrxE
fvxxNR/s91PKihCZnAnwXX9UZUwVZQ+UM98D2DgZJ2KjYEHWvCMSnFVDUKyH
g1tVDrSDws5j/lAkPx4mdkQNcxlT61oiU8Zot9uhKeiTsaUALS+tkBHMbWyX
zBh/d5vWitMtlaOn2te5SCjo4i4LoqVNvpQzyzBexIxJlU/sR3PWK4NejpT8
a5VQTvTglU7dNNwsd5sO8BBwWd/Y4OqaEjooDtAq61XmcfTsCF6KIgrCdW80
6oHP/nyATgb7GTevdSctAk4h99HEtyjw8nwljM6/JBSBJ4DUABw76gVi0imE
uLI2l23xje2+4DjhggO0l5E7RYAlS454G7ZtcyU3HHEnVCX+7bEKvcIR5/OU
kqsteMo4XXooS19SStdXrS0+mEQ1UzOQfzMYZNZINfx3El0ZpE5DL0fjIugk
JMn+GwJbr7AyfXXkt4AwALCBNVSdsuBCXx6CLp8zh1OS9lImsQaN3lOtM4cU
70gWr///AkLz8xvdDuVzsTR7/EbvQsG2gRytA28tb68aegrBymtTsccPWi4p
fz5wKJud0wDXqH0mV7orNKzexTW+vaEV3J+duutuFvn/VOJTM1sC4uKcsDHd
R0leIbB+Rn3viEzIhLr2FZxHMKOEK0EpYZX3zLuN4prjY2MRs1pORzQ/mOih
Mv/ifLaE2mSRnLHE6RDJuuEU7zwIjgxQXA3EQaPTQxeC4CV5hZfLY8Uo3Lxh
wKNJXNax8NYRcN6oxZYnZuRKBYh8R6L0ldPfwf9YTQawAtH0ZqW+EsK0/i05
ISkzn/1O2RiTD5a4MgkBtUwjtOAUoHCwA1t3jsASCgTyv57e8S0xU/ygFiVz
rlm6amjH/1FUss5ePnTUhETDyiFchawZ/LpmGQtPonC8532KqDiK9nXGx6p1
u6PRySwEB7uLGvwqQR3RhXFqfiaoLUQ8hRiJArpUGefbhN5P76eBNSxkJQAv
vElhXlHc2cfDKLL2fAVkm+rmlrN2gKRLzTYfAj6f8DWqe1u9UtDEeMUxwyC/
bwyF9kOrNwtaEKXRjRSHLmH3pSdszPDVKqfWr8dvyoykwf0OnGH0AR97BjZE
uBXBK0WgwB7Wm1cohlK7Q2OMBAL/xPsXSm5wGbyVHtzMQ/gkB+VFKkT7rkhU
HbmCtKvN9WaQMVLTReSBO5/yS7dsas57BwRkiSy1cZiqNgVBVSlgkyXpompj
qiJiV8yYBPMTm6VMJhhXBhg5uY+auNx67yaXFwSb7CPTIPnEuJUoJNYCtUMb
KvXLlkt8+8Q4my6JXkqhnulrirW1TvNeuydW9Nh40Jp9Wh2ljfq8NfKV3RfV
eSGPSDd566lLS8k3NV9zFFsnhj6ON3Rk/9BPhTA3yaL8VR8CjMuILflz1qV4
Bx4IJAEYOaOO1oxvYeLeIO93EImmiQHWIlb4/nhWF7VHK5cAkJPr/VUpmPjD
emUpbCeFLmUytshl0gLXKu3Go0bYgJOZJVQhBegk9uP0oW1qRt/KqC2JxzXV
lO/GqSNruxmE6OlFx5Qw6mm56F02SRrsrSK/166c6GX3KPx4pRWY9QOjK3y3
xVdUoVTksec115t+ftq95NMgSUL//aNelFwoARWbqHg0uzpFi1aAyZhHwDL+
vOi1BIF6E48gAXsZBHrqjCh0/pGCkQ4TbfcL04t06k7fM/i4feez+XkC70S/
GTGVYKN9qR9fxsOBuNrOGx2bTj53621687fw3CucMEcCBAJiTaf5q6C98Hqx
+KigXXgfQs4E+aLjh3qEoTwVOH7K5K9W4h3NAx9p/Wr0lHYS3L7hakGlZzZ0
D3IMNyv0u5NbxJ1s7jYoUynFs47K0b40eP8FzrUVPwnNuaM5V76K64h/ADzW
pL2sRiEaYucxDpH//VmtW45fNuA0scD25pb8w8d3mm+ol+onpuiUxk3lhi8z
QRzj4Jpu889IOiN58xMPwmsbZCFBUpX3c/adJJr/BvoImjhVUMr/NnI5B9ji
l+TpYZ4ICcJb0ucOg8QQ0I3ZcC/1d5W5kZLzaMZHTV7N5zgFHyBCc8zDQxwh
QliLrTwioM0fQJTd+ERF4J77aLK6JZYypge2X8QUeNBFqdZPBwP6xrS8Scda
vC2u+9sjlzamPZ4+mHZKObHtNEEDBe6JlQ052rUkk7Xi31E4siZiW/00YLJc
hzS3UjCby2VP43943MnNDuoMGoydDwWFVUuHDTOeYVAmfG8cLRRxFOaDeS11
3+NaMl2aX+lRvdDlfd57mSFZeWRF8wGSkkioK8N86FvZJPoKVGQqVIrzP9fO
OLSu1ZsSueQProdxtYyXU7QIF55SgFMDsOuHRAsVWJNQOgNpXgGd1HphM8B4
jj2WzGX+dT9KYa7UTzHDz2T1or2c4sfEvLuagNflM/qa6li21ahRuv/Y339u
Byhz/mRDXKd6m/EsDhdSZbQA4pot4fukWJQQnEwMpBIh9PEYqhscXHdAJmhb
gSsxenos88qO741hyAhxTci0Zm/yQlXeqSs+AnrW8qgo8XH6q4VSlAdRs4v9
cHhc3tOzuqb8+bRDTU0gN2TxWZq/bqu8wsOmYFpVi2tr8f0PiqLy5QHvw56D
EYUzWnu0BREmpCM80XQR3mdKIx5LS52bp9rvKLqNp6m5jNDOGASNleyAAW8a
GCnVH1MzGoCTPYa42SlqsEPGp+ByjoeYhK2E7GQgnn/kB4dV+D1xdkNXupDq
PkOxZ6bVuF/PzmQHA65MYWf0KcVRzVnHt0N/RPGT8JLsvCCfrnzHJgXksQR+
BCSSvfUlvfp3bjPRewZsdM7LurpEZ4j6NXi88WHT/sAh9JmLqezsxzI0nYXi
F7N6QRFPO5cJDYJ+vm4Qnl2A63AlnouqxaZise1uwtuqAQyTvNBkXo4mOvGY
kI1Y7UsV1nzzq4XFXQdjMKjXTOpfiNqocBpF53WG1IvVLDD8V4ZXhKTUO5/3
R6qHMY6CZNdFeXm5GnGg60e5omKI7wReV8cfmBybOyKDI6a3ilbLBn2fVUF3
R9uwnrLMSr6LZQPvVfG+3/jSkixxjMWWnvwVRDC51kQnZUdtmqmvjCetP5S+
/y3Dcwx1USBag/Ya2sMoxYEWfwGZD+Xa9qBGRD9WKkWSmJu+dg5GzS9vqEoC
j4+yusMpzdkLiJFAbuAnKMmjPw6U9pkwuQaOBFFYSPh3mMc0HJiQlPm3EvQE
LAKO9+zM8NAB2wkfGdAfn9ENR3keTX7mdxZtkrFRQvxWWwzxrmtRWZBQ0OC3
gHgcHUu3QYzzR9JaioFQN2Sl5laCR9jdcNpMCyAcNs1JCTLCH+y7bs2rt+ui
CLCptOpHezMDu2rSXLGqsPKBpSkzwyrCsbv4/jy8gOgWVXp0s+pMEvrntk3d
se7UKZ1jxMfYka9rSzuc+e6xOgLTK3fs7N5kMasLGakpSsKG4qmbbgHtCXOI
ZjWlCxREAwQWwZlRI2O3dbgmJEC88Zxvg/X89cJg4O7u3Geqh8/lDkDWQ6gH
sK2biQDW+Krdnin7k5xhqYNfMAVKjDaVoes3mOpq5gthUpGAIDLA2w7K96RF
TIRw/iw6+jo+mmf4LogBipx2/IIBL0T5xaUP4KG6GBD5eXCbvraeByK+lVbu
1BQeW1PZ+6lrfCC+A5a1osPBr+rZHkTuuMqRAvtJlO9qnALxxjyBdXayxFtm
S5PnKolZfNtHBCjVt/pCA7MoYV2B2AvQCS8Kl4+yGtp6F4ajCYh5+JRAiYag
7CGNeQOxcE8OR6tc5OWaEt/r3juNfJDoUW7kQlw9IE1M2yV5CCZAmHCjUCWF
G1b+F5N+0b9tj8hb8RN7843lq6K58f0oPu/Lf2PfM+VhRnPjlI/1e1uP9zZ/
kOY0P8rrpdJKxtWeMSnBYMQIWcbsSRG974vYXFrL/GsLUjxcPMqB9S3aCu3x
vC7w7DZb2vEUkNmeaOmoKaZ9rXQRaOeS9xtDfekpMQN18y+BqmTc1sPsv3xE
Qvf+qpHeuif5Y943X8LFU1u5jYTXBNdEdUwN4Eg7dueBKkB327neQm19HCT2
lzN0ZyYeQ3a65Kvjv6Z+sk2uoCkajf2ORjyixQrZE79Xkpb62UfYmeMpjfqs
tlii4OPTZkyL2qmZLFXRkBEDqgZz/jGbn9izYZ+nU+5UKwH+yWMWeqaPl+1Y
ySmjEAZFjydHjtI716+Y9VbllQ+a1LKh62SvSVP//s4/NhZoyd7LT700VeUj
SMgC9uoQYlUOAHIbkjbRRXdmrRCJlbeavGbUim7t2YnDsE1gZIX3KmZCeRrr
8Mflpx/3WDemNkECXlM8izhP43Zsm/+niYFOh0ICp9k6NBWOKp0nKn64g3k3
T1sStnUl50a61kWnz6jIEBGnHY5Hzvapk+qhFRQrR2ixJbogBf7txtW1r4Fr
VdGGb5ocw+rh6iWAzO94y54BSUh7HtBT/oG1bkLfm7Altaj1pd2Nslwv9Mie
t86Od2wubFjEms2M0/ls2HlX7TJfJ1+S4zF5Zzf4oJMKoInDNh4NxXPG50ZX
Am7IuxiUY8b+nLFso+5TZO1pCBS92dNOpkp+q7OvUKcJpeT3pM4HntOTmPBP
Inv2X+oM3Cxm8Ul+nlwg44xe4ga8hKAozSaFl4kNDj7P5DzSLLlVsrDo0PvD
0Zu2v4d5C2WAQ0wTC5W8691QcRxuNHvdZsgIgPfinGt/VD7fshzBaOiuqaQP
b6XRd9rtRKqBqZsbqEzDJzfXnKl/aq3o+l9GQ1L8vxwwcP6IbIVZagbMgBrM
wOHY/tdX0M9wDVTeNn1kLPkf2NGUYzwxiSL2o5OrbMuyqaxxA7/7Wihud9XZ
7il9BymortIMvJOdNO3sJiCNAxua0+htasn+N7vlcyeevVDWdeW/Wr4/oO3w
mBQkUZTn9OcBzuHMPae26KPGhD6Tfv5kAat9MgcbLbQiJiP5RYk92f082e58
EmeFJuq4hvvWKccIq2W4GNu2qwjXpKQDUXlycjEaOqumgFEZV0rfJbTsIo8e
s1VW9OaOOlbJ3FKWO8NsJVlbujR7Pv++1I5YIEhkv3w1CeR5y605hFhCytwZ
dSGzIs3gXA8yEEEAryhx0O/UTyJtvMLhQThE/HcBl/OOUedD8KS/4Jg21OOL
dsHuIeLxXk0YIQVOREIkk+BWexBCyXe7usoq4NE9LRiitM5MIpkPT3yeZXAT
+c92aAO24mCr/07cb5fFMDmkNUtWhCuo23RjrL/9qaSMgbbtPIMwNx0BcfKI
r8M9rswQSlK+eMhgjt/9AaRx47+fLwnijjJJtcCb1ZlPksADdbODEhMrwgOs
ukkxWwgrDhe6OUiu7dguj3Vhgmn7h3/D3g1j7+Il6Rzhr29llDJ6cLAY9zwU
se4vqDOhOp4XuJu3n5jwq1JuFBvOuAlURb6YLd5mSW7wQhUiK9l8p6FwKh9N
Xs/XM8xs8bH5cNbJeRmnQtlFk5MvVc30CkZ2UuY46bXTRD62NH5zt2GtxMhI
rAL134Huv4nfNgvxbo2kV+ABG4SFVJmTiQH17Xx1aszBLJoiLqQddSX+SyvV
cHqXhg6DeweAgBAjID0Si+5xVyWTF5OjSZ/9iFcgOFli2x06nmx+IUHBgsV5
N8ptvz0hjwyMnaqR6QnF9p4HVRPZ6kgMshZvTcg+zlr3zGoLv+w8hHK6zScP
R9+MX4g0i2aiGwI1OSP2I+uyhQ2H6r+6hOGiYH+OmWyZaMzPOOPsF2ynVSWA
mLRLSywazRA8+j5rP0/SRxOZqjC1ZuNoudihXOZNPO9l7ednDcJetdfrBNkK
m7GC6wG0L1CL/TNxTSznLc4kyDJ/2LRZEFFQjcmej6CEe3UROzrhl4BOYKiv
1eEbtaZDCr8TqiadL0aIXNqETdsdMHDJa1j7mGjt+yzj1cdchkeKgDk+mtbe
B5V+9ov6VhjswP4GM4hx/ZTmHNDhS1CURs2O/H0/zqQrSV1X5KXKdffdD9s6
qZXXh470S33Mb6biFsgLC0lG2hMjORTUpjNDiMe4dcN95AHoU180PeoUz4lJ
nNhdhH9BjThTwlXPvJJRbwGQ2EFLrs+6x6nIjpRogC/wzcxc7BjyORoL23Zb
NcyyRgPK4IkmT8mDXtz3qVPR9t2YWrJ0Ms7v9B8ZdF3IUTbl19A7vCuRITf8
B+2CdFwjjx5Oe7Dc8gpoTmTiwNojs37YxYxo/x9aIM8fzHKk4fNkPMpnlamj
AJ65LQ10Ek1xpy9oj1/u8WThyokGgK0JK35ptqr9cltvAknTzTGXu26fZVSy
0sTy3TgS8RYzNKeVoVP2KHVmIuQFdUE4vdghL+ZKWItkxofRha/CnfdbjcHF
gKpmOEiLLaShb1r1OWWW+YjaaNA5Y3uK5Ww7BKn32SIPL5WAqmFy0qtvNKY8
oAeFAkwLFTf+TFpLRDwXc5l84b6XcZGgliUjalRJi02Zm+CB/2FFQjQPFPfw
qD1UwJlbc6n5VEiyvJm+KsLIb3x7e7abrMn7gG/wkMKJHtvpsrDd3egY0UIo
2iE0NdHpfYZ8yYs/F0meBTZW7s7qPHABklZX4MWRsxxM2dX28qAi6Q80j9qM
TOXoxo1q2V9Aeu4z2Yx8rTbPPKYyIQ4R4Ra8lZSY7ZVpmOZlM62OYSSYC3S9
7zAIzkLjE30PVzF2u4KKJjmYoZvDyEJqrd0MByOrisTv7OgAgwPIEjHF1pc5
g1Zggj1HndTohlg7o8bkNAdNYX+LSOYzkgoqo7LlDgQLCkHgtTbuRuWQ4Qw0
lgcVhk6nAVAMfimshzsOzqLtlOamX5H7YWFsSgNvJPsA9h3AWtQI81PG94lI
U1XBwa/r3JaA+Y4S2spJW7XkMMBO4Yv44z8mp2mZz/bfI/0AHTiIlhNgTuOF
9CTYk6bMghmpWVqFClqu+vUhDFAB62PuCGPo9UIRQQNkjPRpud4C03AmbxsZ
od5tVrOUlUcglXgAyy2+UMzhxpnhVTtSed9FuPsHC29KxZYoDemx0mX9Wikj
xO8497jpX2iSeXSd7tx9IAFS+QcJIhivGxDPMVE96BiByHa5ERzheEPELmQe
F1zEx1YC1Ev51tVCnHC8RQQasHDRkcSZ27XO+EMH0z9URRQZY0qpiirTPlJ0
+eRDhCCAXAEjLDZKQ0aqKQ4Kpo9lfXPAxVSrc7EFyo7NLExd3HRbnjrlUcqc
GuG9F9M7rimVT8ODd0T6hf+p9K1Kqcec4hnzNljb1v47PSc5+QVaENlQWjBv
RRf6CInbyoM2r3gcdByUCpc8NqtqdnPOnV20h+X3A7TfEICI6E/DBsPGWWKR
AuXZrTvqffsvl27f4R9dvbpwJs7ibZ4qq+stD75vJeWuNBdBHeveDjx2vpVO
9TwR012HYjhTS+fVlTBEjDilINP+F2uxkZ+WJwseboSHtrHtZQB14wLh1CGL
V3ne5LXauuIoIiIsTMDLDJ7d3lctFQg957Zg/7MYY1MyaLQuTaQJK7qc2zKE
dNqBQFms1O12AStXbYD3130bp8dLqlr5nE0d4QBiKazUZD4llLWBaxx/J30g
4Gq3kr3ggAyjOqPNj1DNiPVDZabI/9HwWoKjPIJAoN0+GtwM1ylVsLc76P6H
FytvHuOfplCx991FEeAFTtlVdUleSnaazOB17FM9OuxL3MB3jnmKXWhs5lJR
59bijnrO8VnduKnhjhno8DxZ4y6FKDnap/8XeAbCWZpiFAevO7nxVtfDjcQJ
AcdXr10HQ0mBSdrWN0G4U1y9ltQ9Wq/7OzdeE1PWLC3a7XxWbzuF5sUzo28d
VW1jC372DDVg4eIL+7d4Ci5IFkIMZrkmZ87PwFLSN/fNNLGdglJ6x7Y3HkHA
QzS7NY74FsV1h6hql0hegNY6A06JgrO7RqnX1i6t+BVlPPQ/17DAGmPumtiE
iUn3IzJeqO41Q+78Wxd9GUl15VvF+BWAnY3qeDmBiV5PIsHde0lXsSe6CAwY
ftxF1sPq9XQpxwkaQrBlvp2ED1O0fZcrvb9k056UjNWnmoS2+kzidH0CMJzi
/BNEWFTA4ko7X7sWomle9JPiR0w02N6kASHMODeI8wM/aEeE66/XRSUGmNPY
nDkxrs9AKLxpZuswnA/5tY0NgfZ/M2o40J7piFF87W4cwytFXDmKiMXJOzqa
ZgT67GMxk1GmPpVywErpmYQqwuAh8BMJpbvKPQiGZjDPlLG5QmsWwczcWlzA
Nk1dakx6gNsxTRr2XlisN4aypDrWOoMy5pbo2lXkHGUlDyZjdiONCc0kM9a1
84QtzaFadk9qpfqBrYzy287KSPcELyrwdT650dWQtkJCH8f4mqIFsI0kOGs5
muMiFMNPZomAPYCHJImFckPxUo2zDVi/4KYWMiI185vY8lb0WTTKzqkf6A5H
dTkxL3gMSn/ZV5RTrkQGQ7wtsSLV7ZXU0p8yEnv9QenoeZ+w2FCDEENuZJjS
mbaXhNqyOd/CcV3eb5DqJ4II9lHyFkzXv/wih4vPrSyF2pgA3pRMLOFNRymO
ao3rE/tYggiEySy8KwBXM+UMIsmz/Ne+AIDlp+rt2sqC/xeKSaa48LKHNiim
FFyA7b8HWaUs3v6HEjPcBfHo/MCTptrPkoh0fXXBrv/P27hY5c2b7GhgJEgV
/xwbHWGst2FQFpW0m9ObVhMiZ29fEi9pkCzgXL9WJNjQkgbxmnYghiYW2B3/
aJjgkParQQTQkl0iNoW4gfJ2v7Tt5UTkjV+mtU30cK4ewyJ8yJSNKRx1yUTc
tA8ZUGwP/dDoUPPvPWKLPoEsP8+b/52RvLTcz5bbsW8NAKWZF8P6RHI0+JDk
1gIzeetfjMH/934Wo8KEqz4L2N7wQF000z1P7zXB3yTmUS+wE3PG/MbuWhWv
HLxihPKmq6L07CGLqA5ANwiBqas1BUiH1VYOKjOMaDz/XAaidJq7m00Avkfl
+7XRLp4tp107PIoW3ly03yTcQdAarzYgyRDwD+JTKg5BcwaUDySc+GkOK7oR
c4SKgvsUPihqrwIgms+aBSHdJjvzQ/fbE8OG1sujwy7tDsH3kZdbOihHsDXb
D/zZpgEnlFbAHcQGty/Bka1tTgmBvhZxXYJL5SdIjcMY6+Vn1C76CL560v7l
vYOzBRS7uocCDZ5JEeiI/PXlsAM4sGfZrjJWGZLdsuZjPjciYQ+D3+u4qmOo
mIkwaHxBT/SBnjmherefrYftb/i32pYrEjlgNk8js7hpMRFYx0SJ1JO8UpXA
PVt3hHgaOaNHI7tFi3aSZb8vW3I6/g9YyoiVFkG25kD7ItiQfh7qZNC0rEg2
mu6xaG7Vc56fWQ6jzNi5BPzLHYx2DOcdUxtPFPNQQvwi7qUS0jobvLNpBmyN
byL98MxjenefN6t7XSYTyHKrQhCOMkvTWyf4/ZU0Ej8cR5kImw0Fzr+fwWP/
iVbKcS+gMxMW+XqAyMhjZvE70JAVHPvsBPFu/rmqgmSMYE58KfISow4W/m+j
CF3ZL0InNBWfxGMAZg6gAHWyLNb5siRG9J4oHXNrU/sG2s6xU29qvH17KEjj
X9q61BTI71AXBPhDpbA3sjy2tEz8lJv4JMZQ0oQDHSCS97NHjbdjNO7TQv6E
80c0fhR7+PWbhdZfAVkfem0W11b7FbMnUS7qZtYuPPs54uUUer8UVs/unsCr
XsTM+Yr15SnnuEc3Vvu5V4YbSrtveFUQlg4Vq2y0Ah1/bZrW6Hto9+xpW9ft
ATEhC86LZf241LWCM6LpXLorGCvzPre9F6LMWfwXkw+AXMFJTELQ2miqlE5f
ypCGKEK990tjg0Hxsjp31502lxE9yzkaD0KDKofQ8bSbJAY/cQP5xWIP3qAf
3yu6T5AVRxv3RzPR53O0WLWwbQMTQaCrJYkAVWdD2r4i8mJBSRpy42Bw9pmM
Uob7EaBkVD9g+/JPMeOsQ/PTwB3X5B1E13l7n82OnZq8Pa9MFt65MslIx/tp
f/AesiodHnOulGhDuBfLIlUeVU8NLVPHz/DC3z769L5QIn/2SNCyiZJ88dXS
+s8CP9KG4X1sfPhmpPaBIHeW8VshAm7FZSIkzV7VFwGbq8YGGOiRToezphMv
pC8Fb4w/UBwDBDP64H34JmPvxq1hNqQPiQXcWdBpYwIZsIiRUTyRFrunJ2k6
rH19sEN8VKXpezpY0KD/IoAwaOP0HbsF55uPBQbyhQaMl4zEenN6PUkC3LOW
oUhe2rS23Aa6y02v9LaGdtUDP4yTjRzdYk69LmMqK6oksyHIk5l6/xTqgeuz
03EA7GFan2Zo7Dnk+F8Elt9d+PMMlwvklMfXk/0f0LfjzJxyb7Ewp3SxW1f5
WZUhLgVHWqtJrc1wJgB+EKwG1+4DdjepwTDKPJLkNMFVnXD4YC9yNB7YQ+16
2tqeh0iV0rdewpy68ALVrW6MgBptS7odkJfsHlRM7dWvDK9UBE25iWBtznVP
xFp2jiVJ2y7XoGlSYwtVzF80FWGyToIMkKJNfIqa3D4NC+9KT6gswLA2ga+T
yEOs75OBKgsAP7wDsq4vFTeOiyQ57o8PUyUvLP8wlbyTaLkqs4l53AocsWIT
8oUTfTWk05I41efQSpWNXKMSBwxpGzlVkmV31w2oh/uTadyaK28DMTI5+dPI
MZlmJwTQT5gSGWNfF57zP+5cx77q4MgjYhXnRKXILWiyyvyuPOPPWzzOrKiq
qOUPQSFKLRhU8avHEtVqKeb3iYBjwcq5fn+8JRCtTtGo/65HeCFj7IK3OqKa
XRMhTRv09bf0qFmltgSUaFxOMkgR9BPQxGlTUjfjMnc20c9HP7k3qGvkr/6r
vaDYo0gmUY8sdX9GLaGAmsEkxYsDpsCGxNdJTGD6PCdp/xgq9xpIJVOVVWiv
i0I1CxNWMy7ApGTquCsTnXMOmg2f6Q7gJNtIj2zAuU/SHEUL8LG3JibxU5Gf
U9AXLHd75TS3QUCQw/VOwjtd7JhRX8Tg2eJWWShe44etMAyOp59T4gjusJud
FVjEwyaOO6ULvnMnqsSVKRDsZxj6VMVByod8WaEYLVtkKprzx0VQx58HA1IN
nAiyMGOzAdO2Ui7+yTvSHbW0P+KMGJZhMENpIz86YkfEBHKcEaWmxNpOhu4h
VmLLFJqA1PXx4nhmitrcLz8kAMoA9wtttRvE2T3A24IjuiXszj1BhiF2zSsM
nsukowx34WxrQ+2hiNAQerLst1RfhAHTrT68pDKemZk16uXFKZXm5T1e+t1r
G4vN9+Qi8xDSRroCJA58h0jU92DdHx5FxglF/vaBDe/GPNQ4eyGD1hjR7pHC
4qdP9JHQ89znjVHy6W6e2QFxE2ciSDd6uTd5kCWtyNvLB4g58awxXC0IR1oW
64MgKCfk5pCZlJfMppJOCu0VZGSUwBRRLGpOaeC/j9hVka/WnYdC+3zG08qX
aVO+NkBxuPy5QePoeTFUzd5nu6+avcreyZINu9b71xDojQVD91PR64WsUXYh
PC1+nqJfFQZrLZljsbsI2fswsDf43jQnHF7zvowkzARKbDrzmgOXQJgkIq6t
yagvz13rP5V4Sw8ogrPQKiMV0sBnBier1OU9M4kead73oEcxvSSBgrWW/wGC
DTdgewa96FOoHZu3uepIm4jFPSr/Fcpc2qDBokIa9hzW4u3nj6q5F2jYlHfN
AHoNzmSk42uH7ZbR2HxX7jnKMq0Srp0aP0wszXe3F7ZHm9DJ8OCx7YkMMK1H
GW5lSYTGN9dgQ34r+h1C3XXedw7ehkAvddATMjXTWpEryBgfToDq6Rrzbv9k
5zj/EoDSQ/Siv+UvqVx0EO+LcmZ32bePJ+WqiCzpieKkggcnT7lt9EOLB50S
9E4j5t1Kku0ZPgFL0VojvmvTZsidUc8QG51dVDrgzkVUB51co32pUvVkl1+q
QBpL3I33jslzCmKu12IYeY2AZAFGTFW3J1YmONGah23tpxFLNX5Oubm9KNp9
hdYUkSZcUnUmHstQNDbhSk4Kj0TXn+Mk0ldudMAWNIfClnSfBDJ79o4q/rHp
KtyyKMFv+jJCVBxUUFZ7B1UlOQYPJj500Pc8Igv5GLYseQ/jAmmP8DCYFgnw
aZxC81rICNCADuMWKuNuoOFj17cD3vpuQ6sy0pCpl4D5zZz79n3Nbnfuhqf+
Nq/1jrMo9IrodUdU8fyPtxzCC02MPayqqaRFEzKWE1ZZWeO1dlDSMQTbi2i8
KRSVp7IBTLmMbowPr77KRfBGXZD1Pod6IVoK0JbR6bUPYl9nW+hZzmFKxcoq
rmcPd1nNinaT9roD/SSIXZW46tL5psaEiBiafcdsC/WbvBaNFpszZS4+27Ii
g8vYBCtjXF0moXJYGkhS2FxWoojsko4OZOPjQVOA85sPjEniGEK8nF/3YLJw
Y64z7r8ytODy1UI+l8h5BKOc9Y4oBd2Tu6Iso3TE016ygKT9zMVKMPZDGbhe
PgRZrnoJYeWJTFDEZLOG2hm3W4c/jMzpf7o6XSCQarKPw7Anuv3P4zMjrN4v
UsRFh/wU/XF2w3wsE1JoZsc/S6Ugsl1YBD1hbBt1N4bDnlGbZ2r8hJ1ay1co
WzwmcTqhAydCy+pCd0fMIimBRP0qK0lcIpmHYDrJpOKCA6dMkbgluFQ41hif
2JNkhIAWkOGOBfIf+cJcZWhjCInKmxyZeosyExraMmwFIYRSqx7ubLJsxtm6
wUNzotyH9bRbFgrJfoQwxZVYef4glX7ax2immsiU5/Vxsx6/xQ75nBnWJA7m
HcC1WXqD7NLcy9Wh7SNRfBb/JiPAgCYpGqjSDZY+byKndtXS6E7AvmFk6ngO
2ETPXcwCbVv7rLl7vMf13J1AkcEVsiZHYrC+9AmFLwOyu4Q1jk/6aH2f66Sg
lSwUQxY69eE929CjKaks0a+GpT8cGkD5TRs1kMxhMVCcrZPzOXnK4F9tI+Zg
ArOpi5jbiiMxFsyz1v7JFYw/spkTsB3hGlbWZIRQ1q6ygzRfWBM6/NoOjugI
aKySbANrlmVu8QWROCrwZ5AUkO+z4eQ8zCPk+M1EY89ijxiuOV4ki28xYa67
5qvF0p1M5mTKTQqWQX3Tlw+5AteYcKV9j48D/eamAHRcyOwBk81Jmop6KgP5
APwXY7sVJ2tVsZkZzZlxdmMjGUvchTTkDNnDoy4TKJCIQ1nPlhvIs3R4F5RJ
i6OGmxAJDFLswcJ78R3IK/hvA02NEmAmFcYsl0Qg7w87lVri1C6+VibuigT3
eXdDxad/Tq8TrZCVe+wWwe7hll49WwcdbmUG5m3t7hecteWTEnchFKeUjYiP
830DK2RzcVFlI8D+gN/lcvMX5HvAgeuus68KCpJPsl3HuKVtZuQ5JNdL6pQq
K9O4sjWPUpca1uOaxGIwF11ZoVeELJgQQCzavoYIvzLYulJ6WZYQk2cbLi4v
0ZpD1/PKCAVbwMkPwnAQvARHsM1/naKcB2tZO+KjqqkDGHh1Ygp43Gsx6MwB
ZJXEhTlKW14mYrfHBxiDbMyNwmGRbzCM1BrGGg4pHxPNdvuk0rVgYUG49HAI
eQNmgu9Y0mQp9kJ9Nn08fnAJ8iYDVfiKmRmSU3Giok+TZm7mL/cGWjMUkWuL
IuoeXCGbg5yy7ebNHyO+KTdD/gIOvwVZjC11iw5RSY869sZLeQVi0qzE5l5o
dudA5XW/9rQbDL3qufLrRIN7mEfIN3GcgIPUQNSchP/7wtGQ9D9VRc1BbTC7
7I5liPlq9v/0RhjcDeNm0RPsrXknVkrQAVMTPMapBwzXsr9sW0AydhO3b1/T
VjfTaBFnFGVq18zJifpoLE53Cg7/R1wrh7rWiC8WZ4xg+xX6AzaS/7/eXLdl
AwP6GR999LHUZQY4WSQeWIG9vBNiWgAlRK04zIhEkRyCC6Xm4hX+wWqkex39
WyHZ6Pzm1HGznIliai+tDs+uwhJgKVQFshfSutevWxNiAs3lJQGfcp8wJ4rs
d6fOwtDfIwZ2TXlBMcje5cdceEqfRzBLqcQlzxKR/dpmXMGMaTBzrVh8KAkC
3mA+b1u7upTDb8DJ6OtH+pxzk+gIR5S1YakMXARIzYwx6S055udYuO2Iyp6q
uou1YQt+f7ZaIQx+qDBcwXF1tdsSyH9ZGoSrQxIHWfGOPeFt7I77qIhIGD/p
WudGnX98NV/8xSGVVE6BqnWCt0bd6zdb93xBs95m11PGWAH2JBs2y612NgZp
U+Xw9u3m1hyCRKxY+Q91R8vIKETYAEPB8KTmUu6V039d05sj1pxPPwDeYPwv
vXWfIAalfrHWSxaJqh0BgafsL07QpEG3VQpl2rSxH5H1qdfvtWXt0RCh2sUs
g/3W4IOaEnaaimmzS9WojR9lOgkrLwBAFIko5p+4vfH/xgy5q/MLYVfSkwgv
5zNUJg+yswqV7NctEYJa0g7w5oWPDy0fIiVGc2woDWQ0oxFhDS3GmY+jLKJC
6MiBadbIXxtoZpAf8Aj0n8y+Ko2mPAwW0p3D35QFQe3FFexOiTH4hugLkdkY
wuDrOGgXc5NAVAVEPDrayv55rYv8g7uAZdkbqfyKxu2jCXETlpo2bRohR63z
3cfm27yzB/vhduUBtf+wkF7y/a4XwVx+uHc5P8ASUhHNWW6/6KlITdU/TNw9
f3bIu5+8RJ8QVGu0Xghn6PoKnbab0PePzWjmKpfDYQeXGAWLDxfSoF4a4Flx
2iDJln1GD6Ia7m09lo/+JzZrjDLCbg9buLLOb+jsDJdrd3edTZhe23DR5DWJ
KJKMP5LZTgfGuyfiAQh3U22m/dLgYD6JHfncqMog+2DnMvpVT6wpVk9z6Krl
AesWyrzpLMC2MTql5s6V8BCFHFprU6QmsupiRFY+i+V8C+VsNgFDl/GS/lDK
fP6JQcQTs8lWTHbUW0ysAz/zB//IQ3qOP5OsMHT0zEoinpn7bOYk0sXlBEvo
YgCuXbwGmUqWlzgt5qah+HoQolNp4Qc8gnlOG6eV61aL0pvD9YXF1pCSnRyB
iEcGtGSE/Xd33ifVF+VjtoZfM5kFttbNBBitYjhu6CmocMq87kOwthG6yC/B
msGyXgOXBomBGZ0mP1pD2r61FTKz+i871KsiHNLOfoln4mHKT88/kWBfvzEX
e3McFk/ft7SrGRxgqxXimmoo+VcwipJlVSa1Xfx+fntNIc4hXff6qecb1Zu+
KNoFtVP68dwMsE8LsaNOWAc1yx1+FJwtLa4atca00ufez4mAArK0b0AZv54O
TEke1BCe/yvuWE6Zhu4lPHJJn++kVqLpZKG41Jheam2nQ68wPvnPMrvg8s4S
4QNx1OVyW+Bxj0+ajEzj0956BZFUi/+u+43Z02XSLKAlPl2rvnUShSQ005uL
Je51i8TEtj5TiqtnMmKX5TQB7l2hHkLOgkkNbJ/OEGkr/ii1f4oKcp7gvt73
BvVoFubphV30CpIYnWgwrPQyQtFlYaM8fxyYpEjQkOGmj+4kMX2jQeqpV0bP
AZtYNMeUwHHEB0GtZRi1by2vCO7AZDs5zowrTHDSSttSh1s5wYC+xfCigrd/
HQdky6+iV6gN8xZD9900/7ZNvN4nSus847KWGao4gPHcX+ifGoRfFaxAiGhB
Y/STyN2u/Zs1/ty1Q6IIar5eKhmPZyjzw0gtjPsk6cShKqwMbMI+kUqTo7Ea
HXP12zw9TOKa4YC7n5kPt8uUx5HfCKptZlYOKMcHwSVav45KRn3E4DbcnyBS
At3TTp8qu0NSrmrb6Aaxyf4yMaq/+JtGRWT5a+VkaWuljb1RMmtxUiqfJJD9
f4Ras2iQJ2k8esmtIYkjtf3DdA+i0FnFESWB0w/o4hOeVFcc2TFXFKoTWLZF
E5KFiWfIr3FtHcnSlta0y/TRolBDZZHutBmzZc2fmpAZp4/JetJoETnef4+q
EdyNXQAwjNKkXam9Ii9UQxkwxU2krMm3jmJpkhYrmoYSiBsZK2nJhb/Df4RP
K+UKFAXHNO0KxhfZCKDTnD3nLT0iMKP3g3RMmECBhDm+acyspN2gUx9Xg8gr
51CxnJVz3iejDcS/YsvkHx4a3AGr1/HWC10PBZFo5CzPGeUJg/lNWNmCEp2p
i29r9kxoVWVzZbdDGwzd9+pIzTpUwRVMedLghcmbUxCY8nq40inRZt95bUfe
KL/M/fKkH1Co4EsP+5eItHuRQeXlHQ1TsSW5DMjWzq68uGrvhlwys87p0NYm
6gBz22IgCU9YSTkupC/PtL3AeKsU8l1Qt4FK5keRsFHo51kF1lIcRtNeYo7D
Rg8csEEkPBzPNaRbR+SqDVkXMVG4r0Yngq7//WZCWZtMVoYiQanerwJgjo9u
w2selPe/gFY0TziwfQdqNIKRv6Ekey9sSV+gL3jv2PahNzTx5ITPFabEB8Jy
uW9EjmV9niqIIlxAODTvHYTIqOzuGOVxhj1ueI12RLDpb5Z/4I2BkwJ4fIFH
Xl4r2+lY8jvGh97L67d9ZXsOIWr/XSePaQbq0Ou5D11tDkzcw7zND2vOju9W
L6XPl1y53Ehz7m6rR4z2VBL9Wwli0scEulmvMFyYeE0fnVIWtIq+PnmboCDV
+Hr2rsORw5N8jydpVdjXy8oYCYBpno6l9Z/D6+LCmSWff6ffEHM7Ds9lU7vi
lc5Rn32/LUc+8RViRU0AophvU3Q+5jCIh9sLMx3SpVZ2z1FBNXr+WCMcI7Au
WiggEgYR5L8T9J2Fl3u0y1j5PRcngcsVqI3CqHDzYJgl1I6RPM8uNP74yOkx
uKAYSOi3t9Otdxq1I55xwTJQ72jEY9xW3z2g4qlxP4fNkaK+XtLFcxsN/31t
zcEAhAK760rBtQuqqjZYgMgdqkz+p+4jrZtCA/XF8S5Q2319GXg4lFo3HFy/
UKXZcPDqfYLQz4vgWSmZFKWntH2bs9817pSkaeJU9nHY10azq49HfAm2uzyI
Y4IQjHbjtn5aCiLN5tSoont0EGTeA7U6Hp9xrchUWm8zO9qiWH3ZM209F3gz
vBSZ+nYj1e8gTicJQ8210yboXZfVVmRg9tUA7ezzmS7eVpDxxIaMw9LFVm2n
RsB5qa8SirruyEaY0EqjylbM5hPpN/v1FSIML12hrR3mGdZLfUINAW7PQEF1
2LFvBAAKVMXmpYNAXDx36VM0MdhJv/8lvpDnh58tvwH9lZYGPHt8o/+n0/SZ
UxVyGVR2AEpbszP3q1upV92cN+1L3enCKzRNF2izgTKttP0jVmwAF7NNiMBU
CzjyF18MD3bojSSYLMAJYPGac9e1tEYsM1ewutTPZFsZ58I1czdCFz/w0eYO
olZZuJxQMhEjaw8y8vpesUoXFTwuC7cqywxlxvq4/9AJkcCX6H03zLvdySeC
SEL1uYFek081vpKS3NAsiO5jK4XPdK/abPa3yRqMHdusy+MXg93o0poXNhzi
cqre6RL+N1Gjo3s8zPsgkNdBZ024iuMEclBUcp7AqYTuBV59xLN+5pwVdQQV
pP1qxUcRtqRpSePSBwgAklcc7TPT5XoqFTwOD8RbsxGgWnfO0oHDC/SVzjmp
D87UT2o/jJjABq3qhUGtluL0lu8ECbuNzmVxeoHv7e48LkuK/JxZpJnQbg0v
qIstDt3ZiqJsil8VkfXcs1S/8Yyf+aMG1YJmdw976o3ELEYiiW+Qt1tNdbxt
5dZp3E9EIdfHQNozaTMss8sPR8CnPVsBgeH3axA8ICH0iHc5+vYFNuFvzkyP
C/QtGpgjsTNUHdJeHcCVLWMke7785f7FRttVzW85vaHcxoH0omtS3Z3hBQ4M
Ybrm7lCr8hJIycFOTokQE0u/FRdfTfnVeFk+vHvggAkzywvauUe8fl04Tm4t
82YkdQj3Jsdo+w7ViQVzLGxm6Y8b7WyZZrpV6tA03Nbu45RCYtwsSM+4yrH5
ip5VWzEilK3HmHxNV+i/pOMcx5vnn4XWHrBAMRXcBrVE2gp4TioCIKNEclJz
7UciKpLYYvCzMeZok+LGj3dwAW9snvwpOLiUsH54ivMe9zcOueyHH6jOYrPE
Zo0dVrC2s4Ol4amTtn4W9oio+Uwb1Z2Ivn4L/3rRLZbi6kfs7hsN+vXmYqjy
uNjgMhGjHLCVR/ejxbALIWnQOY43Mmqzw5kpt2oWBFt2s4OvEGkPlHIvbKCI
lfDZJFrjxj10+5O1TksyQPhBEhl2EL2ACypqcwrL2AJVx2+HaeG557+2EDX3
PHGH+aYi3eZGGI3hR511yySUMsM0Z8RVOMYZP5IImcshSkI25EJ4tycm9bB+
ZZScAjWEhqSlhDZ7GVFL5fSOIZaPqZ6TA2lGeYeTJ//m6KMGKJM88hrmAws1
JLYWBxzmEfihJyQ/Afka7CefxJEcjoDn/+Ng/tHQfcWXaGXPTs7FY6LkEbO9
xkFNrZhUsaG9WoBB4zgbGCLH7zQer2AL5wUXdvBMUDj5Qtkt55WAGX2KBHzM
RN6/wX5MIpXXNEB2sF20K0hB9+HfoaS5+7zoPEXvMVD6VYl2sKpc5kViViXz
wJY5Uso+opLIbEKhgujzx6JFPkf3vgcxctLquzVt1OXs/fOSqsUSgYr1lMn0
hyMmVmQ0D6CEDnA2JRzmb/bI1DuUh13N0jXpDuFzepHjkosx3TlSnzARVZ33
HxHCs9JhpJvlW2/yOvCAu8XPSu+YNsIcEEdHbt0LsqzJsC08gNvyLOiZvq7/
ponNYIxq2ZA3CgyzTN8BuVtt1f/QUmc/k4jXlOdTjNGoLdCPrfQuPBYNtOsc
BOh3wiWLarRw1RsvYLANyJ6EbtshurF+apyh8/3GJITRjI7+t9sXn+yK8Emc
gKguPjcepJtvrpxNchfHJBE/2boZsSp7rmfsk4afl9huuvC7DbOC0jkHqZ9E
tlKosas3uvedE8+d0fi3vLIcROpIG/M8/nbpylaRHYWSQXRXvlyOSWaV8pt1
PVLAt6YjAxqFzgjhGoOA1Y4BM/yT05pciSjtWaMxZ8PY4xEu3PW8Gk3AmVWY
MRq8Ht7Qc+A9RJmdQy5y6qxjhU3nvRMMGe5GIOAKOomnLeTo76CdleA9dPfJ
3j+UumnMCql2+hAuWXIRn6/zZPx11qehAX424hupodrgJT1vSWo8WfkOCSKz
t35PfP4Xv0HhMcYTJ4w0y3kzHudXdbll+PxL51U/fnShqrDMB4SiI/IjILGs
PxL7trRrNNgMaX8PbDLbJsVA9Tn2aXbCirXYkxds2qMu2ydyqZubLnQM8+c4
e0777p5CSnoZjyWNZ4XjsTNTJRM9dd4PRcPek4TO5VKjSwXEbr3TtKPC+WHS
yNmOgp+I2os1A94jQ+6M11SM6FTMqUnHsPZXTpnhNzOtkbXWy89p0hjKUkqf
zNB370CTW+/nOZ4fFVoFlGXjCCEnCikFjz2G9CQvCtDLZ0aKWC5HGgIriQII
LHYqlpHdUeOQ6RPsj8uKFkRrJWjUWvcVLcUJJi2ULlcyYxJ1u+wxD0KVP5fe
WvmESirBG1Uj/NlN3716dCzAInDzlufJCW19xOsBQvB0D+FYZHM98GEbFAWf
+ZHCQpJGN9WWrDUjvN8Wlo1RMfYG6HG9luh9Z+rmbV+4VO4+9YuxKQeFJA9M
3kORspU41le6FvZdFoLA1Q2+Z1KFsSyAWL3TOB7Iuy+VguHGfCvoQAQ2A8Rv
oo37ISkZMnimHa1Lp6hR9p36G2mwQAz4icRW7P9OiYcK31PYzeJIn3YHz+4M
Hkj8qP1Ojf7hV7T10+DMks4RrPOhFOAxE5Z14CAsZF38SkqIGNSZKOszMl5L
Z0NZdVWrtZTLuWVaiz6PDjtT0P40P/0t1wER73EcWmOKtieuk6FkHos/SSic
0SYrhaJToOn0XDSxnEDkoQO1NThmXGdMSuJ96Hep21UkqLpOSDB0YEhAlZCZ
e6l1wSevxSk6dStOQPkk+W1u0LcrOdBX0K2U5a3rRZGiXpjF8vdNIqK5gWHS
jeucDBByZlsXBPqZ5Hjs99l0RuE8Qy3C/njulf6tLESUjUGwlh4yAaO3uhG1
/uTW6zaa+EflDkKWGn5r0jMm4biHDwjTp962OXCThtBWFnT9sj4p87I3pciR
446qlnGZmMMZ/DIJJJNCONAbw9fPyAsw1l9J7h1lunvFIoy3wgX8O5rc1Vdx
rS5S2YrZMqIMlgZIkrFDtUTArqns3Fy7cQyBWgGMgxPIs5/eq0NNLG6sYDCc
aLozmw4GDNmbw1NdSlFEf2z9oRoB3sfmBda6l0iZnL/1uhkLxauvZpTwSuA7
ApCL+UMk0Rg9nb4fAb29S9kpqsNCSNEwrsMjdHQjxqKIMgqxhkksVgjWeKxT
/jfY7teo+Z9n0MQnO2kjSdmz3yaCVI+d6+3EVLNtKUmHor6BuTHM2Hy2/OfT
TGJhp2d6e0n+ASoq6/xgwoaDAKAUOLKj2YtK/JPdx1bsDd++8+V8fW++WKzH
pMELpDI5iu3AiP/sWwsV3W1jmDGpOi3ziJlVab0kNimcpJjTnoq+BMjY5ly+
m9eOEBKjDfo8Oz4WExLVjvHTSSqeSs7uAT1olTUXJq0E8Ypr0F40KkHInKz8
IqwpjNl7NmWnGHfdIylRq3uCI4vQycgdvTEIYaneGcPPuABpvxqNodLhUv0Z
8iNFaB0eQWvoBg6o/SOjh1xcVbDRNO/El+qX9Zol3Bl5hBu1FCZ3CBLYVo2N
ATzjsh0iskcgez36mS7csecuEnieBEgJVakh8Xm4w9zyuLaYVc+2EflWisKm
29a22eQlp4f+LTI712jEev+xSKcXjL7cOtAPQ/vQkXR3D/RdTTX4gLRcQCI9
cmTuHr0DRa+Oq2CC7TeMl715H1if/ljc2k+QOI8qLelNEyZ4xFzVVYQpsoLq
AZhrSp5Ot8pplI2InjEQlITzK70bkYkeAvuL4ca0EKXrBMlMbVajA/ywc8eZ
Si2q1nhFE7xiE5GPA9wfCqkGkEFPq2Vnlh7NwnsebduTdKAGSAIXkYRBB1rn
W0Y+BLT9/hmKHcc/LU3cI1wjWkSGDm+dEDMWdmK9XtSPzsdmEBSWVf25a2Ej
qvYFr9qxxYIeAMHhoUbeCtk12zUFNn24b3pC4kTLtFf5tHDSu3U2LUZfc7U7
9r2UBT/YUhOR2LbkQ1blr59jcUaUqrgJr2wAVzmCAup/jdBfCxiEV2CX9LHA
aI00yH9SgUT4pBvgJVnplogahDO2j8RE/3wyzN2GBGKXs0NsGxLtwBedb2zf
EChgSzhSSjQMBCxFbp3PNC5drvAnwudE1w6g6/4B7eoaXKgf0bbbP6Wx//oU
qciSj8ov3HOel65n/Iz7196Diybo6W8Q/MRF2BUAkawY5XbIlOjgoRh0oXyE
27ZExN+vWhTMU4BvXu5jqT//oGxdK811rN1jkyXmC1XxIJC6ITdmITRhdWf6
VvtX07wCILzLP/PtxIRJ+LJwzg8TwZzFWk6tipXXSCBmRtNB081ZtixyTxyj
b4EPbAegPIxMQ0DlC1r7aK1CHSww2GAcwRpwyImZOai0cS+hGUYUBb/bjL4t
t7V8O80OVoYiKz6aWBZkkQPRlCKT2r+G8sL58ceKzgNjWXAM5dfzLsJc2h3s
g7IeFIAdKBjQM3MYPKthPZXRj5W4eoAGxjfQiNWyUUT1iYv5UCKFJUdsx1Zl
xwQdk+HW29vuFZneVqimSU9wX6jXzfZjPbIrs0HmiKrEI3HPzTdOg+b1WqJz
ec9y1s5h3OKyfAD2x6Pl0J/gkvlzAT6D7Mgq6IQTKFZWUq0TleNptPOp/q1D
R/gPuA4i1O92mibQaxQrzP4Y+VzCWI+DlpIafI9GTO55YCjQFVrDak0k2856
AO6dtMuVeU9arcWCXaVhdkhP2PsMdlaLZsiiT78b6zNZ+wUQVOBiE7zI9pRG
eGRrhq9CY+sEWH5SHXBrbWVgYeZM21pOgRANyrXA7KUZRJSo9dc8JEUy9Y1Q
bR2mBOFIEfkhtzLTxVXieNyYqDVBpD9UnTBtNuZf7sN3Klezt0v2DyfZB+Xr
SYVPPJYGBvxAOMGfz/ClwnubNmOwPtwvH5TXQV2vTPzUgnuoNViNmwyyw0lh
LXDYSIQicB3MztLDD1fIVlysJ/8o9O6G9uJL2S5Odq3IVJbwiEkrXJvty9xO
IpeSqqhggAHWKaQy1KKVYBTq0DGjqRQ7In9DIe42Rj73Gk6wAYfwZxVFxLvt
20dak9zT7Kdgje0o3jw9+/N+gVjHPPJKsbPyxaDQlCUhI+uyEMtDuZiX+NUG
DUel/Wl61LsNVy4Ef+61flf5WdCfX6pDwda+C/f04asaf+id/tRE5aknjw/P
PDtEFuaDeR2A293R8fShIGJ4s56Um6k6KZ/lWoF8A6vxLd8bLmYFwWl9H4eZ
Vc/fcqHKB/bDLhWA6uBcAR9C6LUDYi1BV6lW12muFHv+sapN/wn7OmvQZZtc
9XkgGiyUkBShDkHGjToWZ53Ee+DDaEdZef0AphZO9M8lHt0qoHNq0G2qZn24
eyXiVoA9gAArBixsCMlmWSYzmi3/lxY1M8i1/HFOos+ir9V3mBSH1IScamJM
y3Kx0z7qVzFdg9+WmOo+hmqJ/VenKGmSV2PG9NK/WfnA9ojHIusGWlRQ8C0e
ygdn/jMC9jHE3ky12mQKWKNHiQFNFqtNjPxUztfixSHIrkeP4tls/xNrrZLU
JQO4kwlgtMxOLCuJ9mn5YCQx4a9AC15/YVgZWSXNOMOtyyVu8TbkbjLu1DC5
6+1012iJEkKj7JzttbeC/BkSvaTudvLKJ/BxZgm8b0/sQrN89j3VfRMrq/hJ
3DRTxC2gNXwH52ZZ/KuQRfmYxD84Tg+D16N4BzfJT1cgH6bstfTCGx9TAdSV
Auf7Gjl/uSfrSVLHqX6F9zg01C5fqfXNucrQ8CKgFAjnWsE4ZLGnJ4u2Wvaz
Os3C9042Cg392qBRns92sApl/sHycDXFoofyMhtHXq5k56JoHccdO8Vh27e1
dPyMqpSsmHmsr0Gylry9zuk6Zqz8WQOWKMKZF8VdNMinbvdgjzScVzW/c29Q
xi1BQybVIbcDkkjf0iwELlgKpFdLXaRMurQpIGVhtOTsY39Nxt2WYFDFAbrX
anOVb1O7L4O1xibhClP2SMY0oMcBwZqo8r1Ksz1wxnd5du0jOSRouKUoUjR1
XGpo30tRjrBQh7Ow+KRZvS8AzNICqx+NP8wRx5QFahAhLlDnvndZSyQcX2kR
c9kU03Pgo8VBtpuBGqfuzIRAEri4Dp62SQ1/IXlCmB5I0+9jVyx9jtZN1fxe
zhnskpyrG4hGi3HTDnVmjmRwcCyKji4moDYNVuZ1rP0TU14sXBnWUs2RlCOX
NTgZCqLg9o1QDo26gmijzNHyD72jeBsCGCgrYz22paq/JAoHXmb4pfO5061Q
GRqoA7gAgOaEiGJ0S/KNRvIK/ROsz7WOvpFL+Hnzh7oxVJiw1HemRIqk7cSc
SEmy5p9cA0wKlehQ8C5rnanIPdKJ7S5ruMzUqDjJ/2XQSWijnc0gmkeTjzwY
QhzlDKrriMElRU/VenQxZZ6pT56zl/TvBjW6Z9P8CyXL+I6F2bpqx1rPr4E7
FdS4MPASwdmsgM9uiAPaIMFEEvG3hvY7rD5TUBo1IHOpxkOlnJ9wDfPMc2GO
M96Qh2RLXonvLRKJn0DjsbGNo/JY0EeulUA7szKBeDRllaULRaO7Tp3jGBX2
7UdKGCL/v43WkApvpuTwnIu0hT/tuuuL+6PTSiEW5Vbi6xvwINlSrOSCoiyd
bwcTr0aPpOeik8lXWxvQ5fOJD51CTz8mLW3Fhpe3dpOraID41uuE/Uhj/kq7
X/9nXLDtkqNkiGi02an0p4bH8bys+41hxnaO4MglwQiZpbNlFPav53rhMqEH
4Tw6AS3IdqPJiqteN6XJeMoDn0EO6OcNmbRa2yurrDYr/NEbjeOctc2VJfOc
eA+YVZSzDCcRFXM9jUdoe7pkh95Qw5VCJV/pjfnW6l7ibb4aXrbtgTUEZ8BK
Z0NYVSldy8584Twbp52GdmMHJmAvhqFZVlYfNyABRQDubP7YW00QaVl4d7Kx
RuD4VcyIklpCBZyBo7be7UzXr+GKH3P+xc0rPipmzbgfWgxSjg9Lqn6cbAaE
AAVG+7xNaOCfnpLaXEYDhG3kwl77cvN2Qo/PF5Jcrg9aklj+cq6NYtsS2vmF
kRvkNmb7R+jnih30o7p0R2ujnyytBFChyREpY9WIbwK4QcoZjpIhB5T5vipQ
+d0DFuMgR9Dx1MsfbQUsoxxfUO1JPU66fAXgOtyAo6euCalKdiXW8lsY9V9M
ERsa1ESVzTABsCPOCsl9Q0WZeDUGwkeDHbcNc5JA0cFY2LJjArWMlo0NIM2H
H6LC1rx8jb3u7U10Mm8f1cCiYLEd0DLK/PEEhxq6GduvrNugkCTlLE9ZTan4
i8OntLimPVm9eidyvG/7nHUlvQ8IbtBShgfZrYzSBG20n0Kim7IwlQ7kkGDe
cD4YWeB1AghFMG+2q7HUvm5O1KR0KWsllOlS2DFnHYNmXth4Iiyr1SBUVPnt
bmnyJW8iIQ3Wr28ThmF1611L/y6mnGpImmvlLLtPi9SNleHw7WDKmkh3lvUQ
tDdyKCZXzt4AlXHEt1oQ0PREaXdvRim7U/YZ1KfK1H87qHsUCmKap0zBZ+5T
kwVNBAlKL0eB16/gXhL1P9HgJNXjyj3gwvwOAJ0ZUxrFyP8C9shAU56GzZoX
IRjDd7rCQdQ1oTpdFqsxqyTdCjMyM7oMGxtXfokkD4EWSdIeKZEZbufh5048
aLSDQztJdfd8cVgS4RQTtPH4aYJk1to6/1sfdIVT3ns/+IudFAPE4ar1gZN8
z8SSLuunklwDHfAK9De4Ba4nvwoULRwRNlv3RfDrPo5d3+9PY5YNmcz41i+u
y4Zs2KIl8y22xnOeXu0DvPBJ9vnzkGwD+FsFMJyq2AawftYPU/0MSQgIkacc
Jd2nUtTpbKiuNiU6JH2M/NCz4cE1VjWNmKgWptQFZskCXk5Zg8Sq529gI4pP
899ILZWengomObAy7I0I2dtTroRlnCbR9yrfZukSgRC0NEb4TnIalttgypb1
18almqnyyi9UjIsziDTPOzGgEqHHYltmra2Kd82LPqS5MDxSXKlW0g8hRMmh
qy5ssOlzkQQ5KLYFoyy1tyk2u2/OScq7X/wGKgLZYibKoGhaXiP3s13m+KE9
ET3797sKoNJorwEfFu/3Lv1ckkmsW7utwKJLbUw4wWCGVzqeDRHBZP4KD03s
WALIPLmAqiEDV+I7AenSG5ChAig5QDjouUbLKuPBWaGHB3hM6mVr44jflmbD
2MdKwFUA9kzPweNjzDQ/psxzFYoojdM0noNwz6JTDgvj2wObaw9n3edsMJTS
B1r8FnyR+IkgT2u7qGD9NLVnk3cK7mmPGPIkmpchZhR+yWtwIcgRC3zexAeQ
SUT73tUfnRS2AT8SUiPVb94uTwxH+RgA/7tCQWTeSQm5IEL3s+qXlDEVt4Hk
W7wxc6RWULyPiWk7ZTaRNvBN8d+IZURIVPWvG5mePuxAS/Fp7VhX3TOGXbdt
H225JISc4M84ZTPozIBXHrUHHV9gPxhIonolzlQ7yfUp2ExNwGBaMoCn9Bqo
ciBxx77X3mUKHUW+fldsu0DeDpOlk/q0X4riTzUwzheEjpv97U19nDA+qk9t
uiwj2uluGpuEBNFSriegJtySzN60FkVzrwh1gWncdyFXJHilybz/DlJ6jhWA
5q2mL/DzQ7M2NqC03KM4lgRliGr07VuePhCy9YdfCBybQnkf0ARVa6uDQ3yx
WstaUOZfO9cQpzwYVMWwjkOUs7OKGZGHhc9vusmryrHE2GHip2mcSmSIMtwl
zyZJ9j7ykLS94qvFopMWnFbLfs7HFavGIpp4ptgOrR3msZaMQ6LTP3TZbWx1
a2L3wWbDzkvPCofbW+54WpZyr6A57GRd17NAvAL71mGcCW+S86srLuh3hoTs
fPJOnkG+Fq/b6hYVNPZF6XrCfIouU+8i80Q5jYwbfkQnxlYsnki5DoXiAISz
MjCG0yJPyMmVKZQPitFCH6gcDAIdafKtrbOBkwhnSRQXwCl0wI2DDmJdHnFy
UoRtjwW9vobVB9oizlw19kI0ECaVrK/RAAKBpPdJGcW7vNDdPi/Rm+sSp2M8
FK+Ikcdcrd6Aya/fIdP5ceCEoZrc52Z8m0OaH/MxoT+JXmzUgjYToBPlqZCh
V00Bh7wWVgThZ1NJ9FX3+zrJqIlTq4GrZ0xhiRro4Q2lKgvmkz+BDg7mAiov
qFpTeOl/GdKZ2vcVI2DJ3s7pi75hyjZrKAyE/UFEiEPBeAY2VBwplJH7tiIH
4NUuRRcaeXGPQT2OTYMpVOcmJwIUCGAMKb1R8h8+ZQgWHsI1T/Xdv+HB7fG0
9nZ+CjRT+OEQN6DCr+ZMdN3BcByRA1zqPKbcoPbG1Z6j5UBmoZwugs1ZUQJJ
Xe5VnCHh4rD/EvT0Sw3BL5UPmbEEXV2kYJ6WD04XU4RXNNvxXb+EeyeCcadn
GH4PPzNxUmZ3HrFHRkGFcqWlaU28mTWgTIhebUKk10Kp8vx6LmsTC+B8p0Wj
rWOgF8b0PtuUJmnhdanNwsHg6S3zQZZIArhHP0VgFBn6gMeHzScP5AYR5G2e
vibvkpXTJFtF2GqvexKavIGAsoEEx9edzNx5hvooDJJg30dqL9YCD1BqRuK8
9JCnVrN9oxZPAMjJgoQqbw1JtMzCMhXWQyzyrJoylx1SIsrQitbNXFpU79u9
NLZUdsGA3RRbMaw/uSj43+rqdeVTX8vifPeSHC+UGkRNlYSrRIoDdUSIm0qX
TH3ORtOisNFncyDWdd5gOHiIPjQFDQtihgtmF/Zv5oHMYNfrkahP6UswLC/D
3BbqaYd4MvBm9pSUiJsJOm8AtIC3GwFAWICczR0SSnW5hQqfk/qOWYB3N74i
B/Cnuf0OG4opGoAyrgG39rYHai/FTmdMuQf7RfkyEM4CtFFBJPS0EwByIN7w
4pvBSe8=

`pragma protect end_protected
