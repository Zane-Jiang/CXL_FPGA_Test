// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
FJR3Cu3naEz8M+ZlGNtBbPhJP54hxC7qAihDmIaY9bwonMXYAV7GSCE8NzfuA6TD
rD9q+sd1C9+BCNTfuIGnkm4bQHOJWuzRnyU5kLkXRUZqPrRas2nGspyvtSdgh/Qy
Dh8rKxlvIx1fppWJ8KDQvk5DAGCoJd4PePX4Ar5G0ZU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 9616 )
`pragma protect data_block
DQtrHKKG0oAl4ayYo2Jeesl+Se3taLWakCBlguq0FZdw1Sasw3B1dbWrAMuGZALL
7xiLaRGbvIj1NiTus0WIWbjb5B11fczyEELkIVfXICFJJzjKqPHtUyWuTSBDHK8t
mt+BzSyaeEP/ug3I2Sv2Q2CacXPx4Ox4MvY0AAAjm8Nb9n15W6j/CniO90nKn13i
7AA2rCZcuAjuO8ToMrrULQxVearWn8SkV6XKMVUSDcxxCX4IcYAqD/HPHc0F0637
2kdKxlFGnoWwRn0DsADD4YA4S8QijsSO+Se1yKK+NmbyVOWpOv2UVy5/4cMQGC5D
yMPrZCWNdRLJP3ZK7SQe4rRnXUvReFNMoNYcg3CdVtyJk1bvKItAfVIgZO7eWCX3
qzlG59BjkfXvUPiB0YeZa8UZ0K/7diS9EI+lnPh1hyJpmsOc4XaUFkiC/wCuquUS
k0vrqySXaY0dYg8VbkcI9W73fd2Fx5+DsyNLtNKb5gep5oCvONNLS7P0mtn52WhJ
v1MRdoOQOanqgHSoTL7fbZwr3/xr5+Ey5JrPySqgbCh0QlD79jv/BskQfs6uuQgL
SQJaLOPr9WCYNzFusiQIB/jw50I8MsOGSAZ26CwOIXRAxNudAcxjw0R+sxEf4j7u
QT9CjcPFJ8pMraVq1F3WQrvdlSVR548KGgtK5xX3F0CHQANaSxJhKSNTSURUAzN3
fe6vDn9TSxXj+qTi5QOyiJ1D3arCSBjq2bKLbI51n2mZMFJs4Mmd7sLXgPN9QrKh
tqqixu5bcqvTY4OouFe+DkVXchv+g3rz+Pi5itqIUCkYMKq/GsAGXqPqJ7XkhM5h
k4gABLKwjETvfK4S9R7p8G7sczNsZ2naggT+axfeo4w2OAmgoZJfYHuDajUCwo5s
oSaUfz2UNKl8zGm3dJysj1RzYCByJgldoTCQdvzmwDRkCAybJ7twHVJioCIO/rRM
nIl/Is9koKrzdk6/Nv/i1dy3C5x0Ko3adOFIVikG9Xi/QBf5dgRH+yLkQ81wcvap
bZ5WM7qGfYvY2hI7jyDtdEWTA6IiRxpu9wGa8/mIipEB7I2gF/ot63HtXfs0sNah
DsJK8FVHLySFruFTihLjdjMr/Ei8qviI05OAKVC8dTASozIkuha9vfYi8xBvZFvb
szJ1hfzwpZ6AFsBSUqGCVFdp/7aDtV8Q1/4jGxMf/73D8SoIXAXee0gl7Bt53i2L
bXiaI6N858ARa+1K7Fa2t4fTtfCqL76D3F/0l4t6rtTFPUi6bdTJfZuFn8XQCc+Z
Ukb1I4cO+cu3efQfH2kCr61RmDhOI2qzp0ENNQ1FtUlVU/nGZdOKPWsRNAWxwQyH
E5UU71tUn3duClgu0JrL4pRj7bvxeshOPFpTzktA+uKqXQTwKrwmIS7iHGUo1beN
zObt+/Oot0BmxcDp+/n+r/6kHDU90DksTbIROh8Zo+MaXX3Wu/CFgGRKov7oDVwR
aQltg8WUswATdYmGkplL77DJWGhZA6YV64QTuvHgIsanCFu3GggJ2biGT1i/uWVq
QuvOIJYiLVKLZ1L1oW2gqXnGWo5BdUBD+/zaEkPgV1JFRxhdsBW21tFgSNVgnAy5
AYv4CxT6gKrUtDrnE2Qg2TeWyHu5IGaVuc0H/ZPCKleo6Vc4vT1thx7ZLF6R9pIZ
bFco2//lPd13VuHiqlu346CCrrSjiPqrtN1coZmduZzCKDZCSXDmRqvilz473p2w
SQ5X7PafIhCkq2BCDX4QsPQNkbO2ypjb9K7EKA9UlNYOWPm+/rn/uRLmwUaCm2gL
Pp2HAOz5hkpmNcZsALKLP4HlgQN2AEUqqK2tSnKiBdltSQXtkdmVvL5M6UY7v9XG
L9ohLsahoN49sX+EQNWnxd26TqzJOuETcBaCAhSLn794SRnzutV019zbWRioZkX5
75wye58c8eRz5qPgMEW02f1B/CrVMn0MeGsa7GDAPRqu6bdWs4hMuOp5vcyZkjxU
zof6J2/gePjZet+ZLUCLV7i4djWfl31XfQ7zBZDiKmPFSrMlIAPIWxB2v7z8UlBU
efxt2Lr5I3e/80FZuOu4bsqpRWEN1qhMxH70qzLjHtn9xlEYXI0+gnO1NzN/qxaD
FlUAfYv/d6kIlFQ7DY6oeNalzKjyTANsoOySfZF9/iJzoChiYWlKKG8Zh+cttbOO
k4b201iahWdvjY+C6Xg3DqzlTjNaiJ2HAdyTHbYdlDwuN0pdAsLodeMscM4zT7sI
T+vqKwrgVbP7JrlXU+AYfmVcdAuhL7Zqq18u2orhi/m3z4bmvIWQVjSsPCUwBXaT
1Cm/3vqLeT/Hj2ENRyIkgJ1jL0aijzTUO0ES/L/bBU9k+P2vZpssliRaYOfP4Ubn
DOvmLaEy9kQxe9vB4Qg+UXmIhH65hLChtdv2HOvDJt9VgStFCvQdEX2yYKVvGGxK
KytUWnYo2+QtfQ1Z2QLu7DpuIOMIyT5Zawma+Pe8epCrsGIKEksA4YLFsXaEGBSi
Jwt1DJAgBRNbvfZWaRo5KIN3y1Z+gzFMhyWU0OnbzaCq/KNZyZJ6z9PLhFx9y60z
Fl0ZHQCx5RNQLqC9sr+nRQhhnqBAZ5gBcjJsWLjw3YXs9zeYVLr3YKm8u/J7Qtg2
junxLSBgtc3AzFrCNAkz/arb/0UuaeGDnlfZnCmgynlKd70gDCzbyS1thTn/bLa6
OOIslBLJZ01a5bVmgCr2qr+hfj3oGVufpFLa0Q7kWJlmeOitZnjcB1hgla/QbH6S
3E/pjzEM4CxOMeVUQCi5Z9VaoeR+Ptynr2tH5hvkWbTNNzny7drWU9pcRF4LQME2
eZp9CR7N+1EY3FMY57VDx7S0Faq95mnbCCIqDPW+HtiS5mVzfvhHd75+r6tugeTs
wEu+6Z1qlUKGUOtwjznAtt8Pt7LrRjZR9EFn31MEBTntYE9kJpeBaAMZfDkzVXCf
dPrF2X3uGRQl8AJddDdjZsBu/6f0NpfrvPGOBs6hLMkIF2Blafs+gRdZHtM3fTqm
YEL6KpLpeGTSpoAHKDcoFCZ3tMve8uz6q+XiVlXMAS54zmwPp2v/btVSeZlygh8w
Jakp5lfJKO6uN/EXWuXVkvS+AAfIGzuHjpgNs1bOcYBKWGUVRUqbhnarnwjhwK+d
4kG4fohn+UnAiTdOX5U+nlnvYsPgAlXS7mBCiz6ZQbgsJMN44R24EONdCmbx5fn0
iF5THwXzmPWoHfexcrcU8wksXJc7uEq3m+Dz/iR+v9fMq4oz787qwQokV8x1GmeY
PUU57FPGGdxKlCxwTuJmIfgj0P7vYDFd/c9Pkwi6xhCqaC5EzzdvVwHN3v7UG+V4
3ic7IK+RPYO6fmfEux9dO2QPqY1DxslEU35T4QBreKyCnyvlG9LGX02HJq5b3phi
nLcHSjXQ6F4K9IhLr//QcQcOJQmvF++TcspM3T1RfXjcapNj6YPR/D/417FAcl6w
5OVMhd/nozsEv5SxKClHJku3S+6u0QM74XpZEtMgnG0fx9f2oyuggBUXie/cOxpz
CiEnpwefEKxnxfdqxaoBl+838WsufX8K8iSUjYVnp818g5Qte2Rq2E6zWTkuh8BV
2zcIOFtom1jNc0PW9NHkz3xs5sPE5NoNMgYailHccFIQNvOdKcZB7Vsgo5zm7qXF
9n3ZwhhuS2XYDCROjPJc+zkAkXxq1NuzsaFZ3EGYYRObSq6dzqX0OxLZMaDZbIkq
ev5x496Gx2w2rtMsO5hYAZkI3B6/xUDsw0nEXO4d+lzS2PMe8AEir6B6U92NR+Cs
dhYDQ71Z1FJs6v9mHu9/gD7D4RolIJvn+nTnLIoJWNpyxGpuGJ8tB9BouAfucvhB
aHUyunFKbPru7UKimOf1mPjl2NpWYVmrvud+5EJ5QfKkWkoW+Pqomlh1u0qGmEEb
pB9ABvIsD0DVo5KmXu02MkILyvZ38XIdRdpgJWyoDCOXxzXscp0DaQ+cySBm8hfJ
Oj1mPApO8Vpm10OGwwsdxLgqYKVthxMav3l15G7aI546apnywp75bcTlWKaaEDmo
dIC9G1HKcjmj8DgDnKGI3e1le3CwJvqxztia+rc0jUhFKhX7Q4f9HUtuZt41gtHb
FJwdpUIB3iC+5jXBqEdZaNznm7wJIfqrXl7N4Icm6gCKWwhKqhNmrA7fMAX9IKhh
WwFEk4GShVp+7IUOzFDBKJnAnT2xKDiIYD//TDGmScVKiCJX22gzyl1EsgjRVfMf
90rWi90uhi2hatPFqk1DAgYYKeP61+BwXZn6kpWe4dMY1dl/+PXN28LTmiAeSfqo
1a3CJn+dP2vBHdYTjoPyWL8rM4uBcGAdcj7PPmjd/y/dVlCOK6VUAXk4AkAC89NA
EZRavIh+dvY5Fon5Mkqr2s52HRS4JaFEoJ19UGSHDGygbI1JFufVRDslK2GXvLut
+nq2Zcc+QHcc34HhNTzbUxPkjv9EW165zRTu/ELaBdq1eCmruVPBk40Nlz6hCjW1
01p2qbrAmsznVHWvXKvQShlVz212ZMR7CJESWylfkik4gMxQwUJmWsJRuKIfiu8d
pslw2b8+AEiOPfTjpal4cUmYWOl29Zg3MIKJd8GY52IVy93Kf13/BBnPqnfL+thk
znN3Sck9amlMWg+Fo0q/In9p0SYBvUMoDkL5RtbaZv2nccsGpVErBClpFpnwnz6i
5C/ZYfz+t5W7Hnrm9yx6zjMgwzhygA7pZ9ZJegg+9DYHO48uZOAJeKkVAIStpUTn
ZGlz31qC3u0uYawxPlwOK4m7RaLxIIu5QHmIqV/Q+S1BzHRRFszZTk4aJqjGAdMA
j7Uf4CDhB+Dg12BzCjW6p67YYXPJaXeWPdV0qgvRThrYf7StSes1XmxBoHuX5+DX
Veq+dlMlS4+aYQ/p1c8A605InmpdzydG1TMPAquxEjH1XZBTwXsX1twV7Nue4N9Z
I+8B0yFdDgfyIasMVeKkakT/vi3RBxv/1psM1nkwzwE+i6gyK/brq8d/EyH0iHMZ
T6og7TEuQuamCv5fHAPtrXMDIrjkXgkYYAXsebuvfm+sx/QM7PK6SFJ50z7+edtR
iQwJ/cXViiVMsCI0QzwaaDbJ26iE/yV9VwIRg/YPJXseT/LWao85K86ZgCIl0LI+
8FDiWSco76jNMay9rHaR7tE96qgN6ZQSKeW2wdmdH8K/9mBJRBfQSeg45aXa2snf
HiIqSvwJuKUfK/0q4y9iKOJDA+3SMRdKsK0f1MsAG5JCzLONHliayArU99RwzYeX
A4sMdO7aUpTZyYy2bcTMAKPe8re/NU8K9lnsMDiEALvlGKWkVreuINggF6dHrH/a
vFt/y85+1ttWP59sDtFnET5wJ/k8ljDC2HGD8XdQcsTYNSSlB90t9PBtSpDE2cgD
4//79nvmBjYpgUltF0MghW74TKXuv4aCgsDlbV343QbH6/nh4a81eMiYptok16Fa
RFC3TTzmla8FJl029n4XgO2Wj8zy/oAZHxU4bw2uU5fAFJ8qb0Wd8JVRGaO6zPow
jYXoEGYmnUyiW1oFz7jvJFb4uPU6A0YFMV0SJRGXSh7sNCmkKaBra9S7PqKPG4xM
AbiNsKvklWX3mxB6Ov4CZa0YaNwgJP9a2ykTbDJ34kNDh6HhLn2tUMMCc6hVHQIr
H5xCFRFXSJNaeYeEvMUfHVNG/5URLoSnqun2FOiqg8Cv2MBMP6gD7GWykbVYGKXu
qMnBvTq8SICsaRyZPGhPuMhONbK1Do6aXPsvyOugEGEHwKnzZ1wGVd4YaO0bqm6y
hKqstAVrDw9k3ikoGXV4U2QTMLpEodIQig8xBFegGpFjRg/4sIvNB+XLZNffSdlC
dJSEuUA0xip9vaafGrjt2HzulinaEghBuQKM0/WQE35HxZDUmApsEtjQJGjcJpJt
8h5hdKxZOWbA5ckvMXy34DtyJwvFxYX044VtEoy3UOqI/2mOVg8JZ5RipcLLTUwf
iKuwVGjxLQdcQl3G9BOLCtxzh5V3pjQD8fUw+3IH0xorLRmlj3OiRJE+caaRFPDD
megAJNCh9IUDIBl2lsbWEnLMS8WflfCMmd8BoRQPwdkBMfMhSGhvuAP1CCt3FDaF
U2pmvvJLCvnbyOOAe5RUvsxEpheCTPT2vfBEUn4ZBPt++hwGzryJ4mLX9nUbjMLf
1gerqXKzPI0q1BdMr59arkHU9bzlnn1qxDpejkkZgha1FyRO28M053Au83zZzT5u
he1HV5+E65JZKIwNc4zZJ1NH21anLrIYITZQe0Cr7TMefKOPhmvRV629TsmLnS3g
uI1GQc+eoojCV9cg/A1OvFtgxD/HgG6riY4NxuwsqI4NG+hNlRf1QTY4LakZrFIp
HOrYbrmaBpWqKfoDB7bsrgQZuaJed1LyYnteXVXkEh+wTmMeVJ59gUwEJT8KHpJ2
MGILcqi5hxexO5DgeP/cnwmdir7Qvd29jadeGhXtO6LxeLSoO0zcUoGH0sUG071V
1YuKqVL1r1HgJyTnQjsGedJaCd+AIbSb0m/G/3oiSFpjq8WgHOgACgBKkeiOxzj5
6XqriYuSEw7VhY1T4CUS71WDooyOLJ6ojhC2kHrZ5MDS89yCCX5AqCw6hBoSk1+E
Vyye9LJ0gboenDy1cfSlM31aIfOXuBzr+WV6aJXW3TM+OCcjWZtO8mpX9XsPVMb/
Adk24N7sSbO2/o5yoVqcDeJKQ1jgiIr5CmM4mGSJjyX/v5THMiy365GVYA1e6LL+
wCD3JIT1vTFFFv/cVN7VmwEB1Guc3Ao5k4D/H0KOGsbaIqWi0L3WhJ8w05NGlOFa
pI5YdxqQh2oZxcUQHuprqzRAMkzIIAJ5VdGv4YCSksT40hhtlHp+aV/vi90Nodx3
yF17NpP8eNrpduzJTxjXwNtkdMiuoHlPNSV0Acd0g41gE0vXaE3f8RRf0Zz7l1V1
Dt5i1jFAZL0EZzWMTPjS798bWdhOToFKlOAL43Vc6CTPgZtaxvPsJWVIHIBBUvU3
Cy9wPjAr5pEULlZJoR7FrGB20Gshan7O7UHa38tS4bOyUOHBHjyEtD6/UHKRt3VX
QZRuZE851Oln08l915zyTzyAnx2gqDlpqKsNIgIkf6YpbAazfbiQt+QyTrUGsaSk
tRekLmpI7NI3AJ19EbcOJbuGh6ydlr4FPAd3nAc7CjDmmRS/9cgj5kBXLTRr/yqY
K4oDHTCaPy16CSPViZscWLGP4K/ZySi8wVsZ/5C4qLphflpn/zc5e4Geb8wwEVEs
l0YCYttqiK7OsHaqIpqUOpZyorJpbpyOjh82SbxwiQZqfAdcyV6NQT+UkTWQu8Yw
4S9PrAWSE+uEWPgrn8hMa5pZlWZ3uAZg64qCgDi5l34jCGZN47h00Ld/OKgRMLwZ
38V4xau5QcZefRh4M8HBVWGrvycGprUWTNau1vkihZFCvJS2vVsgTZUB+xLuIlvm
q7n6JgjVv51sVZOKAynXLOiAEaeO9pyqVeXugUt5lptNUjzCvBTCwIhQFI8GeWNu
YWqI388KH620tx5dbBdcSAZib9tC//dWzheYIEk2keDz3ejsOlatfbWQIvMottH2
UbQQbsbIkiWLsf83WAZOApoSFloWjemRCBEe0vtHRV82tvGaiVONsGTU2E00UU76
hDhPiXRgV6nVtlgBLjsEoAy6cfIDGFQRe69zed6mTnagRgkjaMFJ5t0ibqRS3l6p
OU+9F6fK8IP7EWNPSVsvMHGyvbhDFQZGpRjZL2Asip99Hf3FDsm8AfFHGOBaih+/
vl7e4JWRu4qmlACFsJoB5MZA5NJe0XPZ9IG9auWlCezC6P838qEnZtXRabDzEM7Q
w2NN2DoHLPZjYvPAN23H7khqe1S5MA5QFPSLF9mvfZEiHLfLAxM06WjEXZrwveAh
yizIbb3xgr67k6lLADTU4prHAY8jjxI2PF73eKOn4mCxygKlJEESDB6JDivXJNGY
f3L0ZzfCiyZ0N7ptu1323Qp5Jo07o+RMHWRYKsbejQPg8Lehnzk1Q2wQmLhGHrDY
tX80s3YAuzo5aJY5NMzKt6m1siPopQvoqSPCySYmcmC8al8HdofDA2G9MqRoqFuQ
a6zJyaqUXdrLwr7dWq+72DxY9pyOl3gx0v+VjJZP7mz2PcwwTXKrxjgVpFbPeDM0
neJQUVgaVf1rWGg4b3oO6fQY/2o75ZMImFs9nkAbw29KvBTQ6sWh959oo1Pybnd4
BvqhRFa2FZLAWYbZix4cwjIc8yScVgJ4LcWLMNXSX1EbwyoZ4bgSo/cZWS0Pycr8
+7mqrr7sY3qjPJxVgQfHBxl1OoUSIilTAaOk13QxiGqsBLAj/PQKT7hq1Uckozy/
89eWrD17BVY5+nvEXJwMtMvEihW+3Bse7ZekCJElgB8SvTNhf7++K7blRRIejOy0
MXVfkArkTy8V65uROIAEVY2PdvKj7OFKcAnj7lhWsyF2njCTpVMkQODJsLNCHRqk
VoRmfArNPJ9myWjZf+CkJqDfuh6WpdMbRrxs/0s7gOfCoB2kKwfhTYhoQom+zpUg
lm3ctJLHotGU+ziYvB/uCCd7JCGSWSE5ojejYMKOotZe1J+VeoTEFCxO3sBWjGxU
eREJ+fHOwgHB20Jl1pIpSFQ0sxu1fk2yd9KQ0fZWjhdw92MoZYk4vqbNiTn/BRpU
HFc9vsWHndcfGjY/Z0MN5UK729VSoPWSs6V8b3shA9ivUZcJhvwyVzpbkit+zPEC
leY4t9LJ4cw9KPp8z6Kwns0ZpGQoXDPyHp7naCu7rZWXtmsO6dhPX88N2YnByCKC
eVCdj89ux9TKeFycTeQDpOKxEzhSr/BNxVSUSVidg2WS0GEkcazbqzYuakyyZX9I
qkI/psydGvaOI6o+jf7pXABV2QMp+cxRT1X7qXqmXvkaD76t7O9VzrAnlDruU9UB
Vk5MbMG9Ech3Ou+5LW+IR7L8HsCBQqMRf1TheRVfs32MXLrujvK2GsKDmit0qPrV
98PDxsjpcVLl2m1EEEkJzZsug7As1XxxcpbWtLjoNfY8AIaWgZeuV2cWw6y75hMX
hpr8S/APLNCfqYOQw2QkCR0QJPwMbTfN6MZnCKVsSdFX7+7z3OFKTbxtOYNqwddi
uG9Imor5aWzVMXyStN1cufE15dDXyH00RPvkQILJtDdKDuRFmkdBmygjWB+ky6B4
G4fYSPZZ6GlC4KGysaD/2nYUE1u6LcKSew6TcilCdzh7bEm5dFO3Y54FFlMwtXHb
S8psd9BANJUrxaJ+MlZ4fAJ3CDsk9Dit3XHPdXZM49LU9VR2aLaM7GGrfplYsSFy
/v7t+PZVdQ0uJDulH5ltQq7O7BRWfVj9tOuNDKDVFVyzbDunDB8bXqqLTUNX1kEN
VoflrjQVwVNhh2Y7g7W/YVd2GMkCq6fT+vFua+9y8cgBrMefz+wZBIaTzP48kVd4
LeEu7O8EZBto5hm3P9kOEPoqsOd7rRx6u1cgJVH+cWO0n20BBQLkWWFqYW4Pbcrn
hQb/OW5RARLo+c4vYVFnPsLZ/NulJuezptaAcU5cjaH8fXv8uU0yZs5h1QOmUl1O
rLEsHMPHY24CPtdsK5ynST2Egh0AEDI27MiuVzqq8e7jl9Ypt/sKWlyDWBMwKwMB
6jSNNBc9meGypnaFio2ZkasL5D+0RbdwCW1v74Sk9v5w9+3LlJ5fKai4ACBi+btv
8C2uzClZAhyQb5z3BtBZsfpIY7sOSmjeceQKSnCqZKcHznp3SX5FV0DZ0NcTMnqW
kn1WmlIFKVXEpxj/tMhhLPKzh9WnXVYu9vELTRbCeJ5fxvkmAaJ45WvDUoHnRr2P
LLoX3bPaoAcbiEVJqE8E1Hi65PbkQrAuqfTlvQ6WWX1rfbBkkukM3YLDRDLiy+EL
lXoqFEVN8+i4v5+WTJzb3i8I4oyO//x0x7gHYBiJkJDbjC1b1Z8bVsyC2Us+UpSV
1E3aBREm3EUWsjX5dd7DNKikb4MWojw5jWt3JuQb/6zlkkojQ611omaFNVhCJ4n4
DPh2rfHd6T4tUj+cS6B3aRCeCCOEXheY2REukr+88R3Sn0wiEIXa6Bt1pBel1FoB
MK+xNW413h7s2Uv5yrFGujqWykahv2bIdjoeRgFkAEXmFWWnaa81KXu7bNHtwJSQ
PbIEKTcj09d62q4w4p2emS558imatb5bkEWrE0fMK1cRmE6iISxjcgyzTLj79kh/
LgPijyuO3tDQi/U8SFgZS1gsNiSICphsBUgKYrsk32/7Y5SpOdYOD1sJiE3SzMPe
fX9qLKVPep8zkL+LijOG2Gw1akZQ9D510sUGrTosOm6oERHtgA/p2qDgH38neqTF
STeVXaS57og0ND5ULQHBMl7OtMT9WBg2BD/XBYX0mENFuAqL9cu8P3NNw3ykbFOu
zsT1Pg/PrNgi9gx/819CGi+mwVxoRS0XGLFhu9dWPYgEsT7Am+nW3S+pksW74XG9
Dn7liorDZEvDLAAQjcZHCmuVDM+69tv0DdX0SDSIY4EJv9cwkJzjH+CgEuf/+VOu
XvmEos0OlbYCgXqxtHKwonzi4+yGwLivEi+wz+0MMBGfZPg9GVzArEybXJsfV8Mo
li4P9BGzqYUwrOpQ/tFGCJ04JCasjwcGT+/5r8UK4P1OjQa/BnyUx99cm8IRBfal
2G68DYlymz2JQ1kBEjvQlWhv7rx0398yjsu8Uu3pV+LuzLqp6yWoCv2ESV1EmvaA
yk9eGLvgqEJWQHgG8SKa2aEtmkH5RD6G+zVU2j+2/Yzf+7wCD1t6zlrq2sjLp7g9
Un3+7w7u7p6cxTv0mE5OMiGGXW6JvgRroaBBLg691l+jS8MSHo1rDrezW5UVhYZz
nGCdMslKdFbL1jDqoTEsnE/HBfKN73I3IR1/Rx4GwzvdosM9cifdy13IbrJefwFk
uygsNXSnytuCqnGeicHkvaXKWfPUncTvVQ1RwwaafNmnUUibZII2rpgxiVeN2R9e
fpL7c5ZOa5IGv0dyW+CQWGYVp39SPIqEqYBlkcSz42q81r7NrojWYr9Kb6BkYoKB
aVWjlUcp1pckKaOKEb5aPkGR9/IPnMbpKJPDlVlK1uko0YfZ5MgM2XH2paZcZTx9
ZH2Iraqclgd+upLXq2l05YeGryjQOt2YM3nT2+TcrK9NHnirRbG9ZiMg8s81AiE9
93SdNUxWngOSYBiJgK0EnTi539xEB3LLQUWcp+wLKN9G6XsOEJ6M2iGhoWzEfDZO
7VZ2RdQgRJa51EXqlusIUgu8n54sME0YdUg9XoAGFQvC95MXioCrs3Xde6frdWKf
aL5tn5mJL0RZBDJ5rlLQ3YuS1S/d+VoW8sRXU99bK8nOW3O3cqPW6jpChpJptT/R
/SB66RoE9JVEJLZZEgmeXeetB133/KI6qWhwPcWdrw7zuqiUqE4sV7E2g/7dI14M
STHBaVW73VeOynRipyQpSN1z1JBL5lkyaExMAWjC0urh5ZO8tdkC+cywUU56HUKE
+dl+hIHdqHOK0pZj2luCG4QESb/Q62nQGmdceeSzAdKs0p6bxNYtTmGkkSCfptU8
TJokAWXEpjvtS3xnlR6TahWPueDEXaxV3Wg6DqWfth3v/GIG9u0Uv7WrEGLmSHOm
NuHfQa3lrs8BTOFL2nFuU52CyVgNTQcXP57XYcGvISS0w/T2e9SnrEyGl3eY7oal
Vgk0xliV3LHbkig15rhQ3F/8Of3fw92K3eeWo9jyT2+dsu5qUJLJlyMwWM+hyHR7
hrz7MdG5ocm7Lt35s1yK62kgkUxeeozbANxwkiZuu6gWmqOWv8znh5HmiChMW2T0
mcV7PjJmgc1KSxffElL1iDwTsIPCRdWC1+PMH/TUqqVQ9jNYhW6v+3NXJoS2eCaj
ZMMRa99URw7/iauvBpdy104jNIaQ67y1QmfqVhpZc0BoYAdoKj5WhbErElRjsqTB
66e8U4+c209z9q2Q9ociBU07d3G9sfYvrMLkxCca4afWzIFBXuabR+PNwEsUAXZT
ouWbNAPYoh2gjPr8S6YRin92yH6rW6NUVjutkFNlw9SFJcJFZ366ak6tzb0Yuttp
o9L6i5QzXDCElP1iNip7jNmo4tfrhymikGcJO5xuJgJqkMrKtPE4RkbNCCh8SK2y
61g9qErG9DC6PtEmzVA5UnehpKgiIzWYfXJoGj+Bsbu+2VOYKtMVfvrmNGfKnIpZ
NMB8XPsIvAUu4bnjpRzPibIul2wCc86rDRbtJV2IPYN4Gp5sgNj8dRziDY9T+aCu
gGJxkzDxJJcJCL0uHpCCeCf0GKcB/36bceW8G0HxdJ/pp4NTBz8i9ONbiYL8xPi+
UK7JnWc/hCsuqKP4Mk+CxBj2cnmFjvWJq/7dpapDOpbOoAuaIAWZSuqw9XvvCyHK
91WRC0LawxJlXHKRWT5NyAKVhd4soQgj3r0ItVzWV72EIwKDUHthZsfyTskVpPMG
mdjYLLhAguPcKX1DHabqcZZZcrWflJlbqyDmoVpORPYr/w+nguDX5cqk6ppBqTiP
ul3FfJyNaoRJQz/Vy4sJUtWtbTtw/PBVdqOuxuaZyHGLZhsIE7mVoXPwhv8eC4dX
enkgVG6DOvFg3s3luQzxA3F0o1CXVnJSv1y9M4CtV2EUtClT0gDJJGL06URcfN+t
p80RT9+ipqlZPVDFS5h4UHbb/xAuyRczWLn4NFM5p4NjsJChDMXU0iLFAGUu/f5v
xQXv7HcNjO+sR2ogiojEJ2EKgNYNrrgclgFHE+/lspzblZw5PESVEbuZbyz2BTvL
7CtoK7OSHSP/L/A4JmgHEI3nMYlkoY4e+fkz23FnSRyGFKWttsl+uW9JnqsCjcT0
KJ2vrbQ3W9X6vBNfOTzMBA==

`pragma protect end_protected
